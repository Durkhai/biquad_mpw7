* NGSPICE file created from bqmain.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

.subckt bqmain bq_clk_i nreset vccd1 vssd1 wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11]
+ wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18]
+ wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24]
+ wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30]
+ wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8]
+ wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12]
+ wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19]
+ wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25]
+ wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31]
+ wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9]
+ wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15]
+ wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21]
+ wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28]
+ wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5]
+ wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rst_i wb_stb_i wb_we_i x[0] x[10]
+ x[11] x[1] x[2] x[3] x[4] x[5] x[6] x[7] x[8] x[9] y[0] y[10] y[11] y[1] y[2] y[3]
+ y[4] y[5] y[6] y[7] y[8] y[9]
XFILLER_140_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13855__A1 _13761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18869_ _18869_/A _18869_/B _18869_/C _18869_/D vssd1 vssd1 vccd1 vccd1 _18909_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_95_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20900_ _20961_/A _20961_/B _22937_/Q vssd1 vssd1 vccd1 vccd1 _20901_/B sky130_fd_sc_hd__and3_1
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21880_ _21880_/A _22173_/B _22057_/B vssd1 vssd1 vccd1 vccd1 _21880_/Y sky130_fd_sc_hd__nand3_1
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20831_ _20830_/Y _20840_/B vssd1 vssd1 vccd1 vccd1 _20906_/B sky130_fd_sc_hd__and2b_1
XFILLER_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15830__A _15978_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21551__B _21551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20762_ _20827_/A _20827_/B _20827_/C vssd1 vssd1 vccd1 vccd1 _20762_/Y sky130_fd_sc_hd__nand3_1
XFILLER_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22501_ _22501_/A vssd1 vssd1 vccd1 vccd1 _22745_/D sky130_fd_sc_hd__clkbuf_1
X_20693_ _13022_/B _17007_/A _20697_/B vssd1 vssd1 vccd1 vccd1 _20695_/C sky130_fd_sc_hd__o21ai_1
XFILLER_168_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14446__A _22965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22432_ _22432_/A vssd1 vssd1 vccd1 vccd1 _22715_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13350__A _13350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22663__A _22663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14165__B _14165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22363_ _22355_/A _22356_/A _22356_/B vssd1 vssd1 vccd1 vccd1 _22364_/B sky130_fd_sc_hd__o21ai_1
XFILLER_176_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17521__A2 _17523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21314_ _21466_/A _21466_/B _21467_/A vssd1 vssd1 vccd1 vccd1 _21316_/A sky130_fd_sc_hd__o21ai_1
XFILLER_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15532__A1 _15530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22294_ _22294_/A _22294_/B vssd1 vssd1 vccd1 vccd1 _22294_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15532__B2 _12571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17809__B1 _20972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21245_ _21245_/A _21245_/B vssd1 vssd1 vccd1 vccd1 _21247_/A sky130_fd_sc_hd__xor2_2
XFILLER_151_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14181__A _14181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21176_ _21176_/A vssd1 vssd1 vccd1 vccd1 _21179_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20127_ _20502_/C vssd1 vssd1 vccd1 vccd1 _20249_/B sky130_fd_sc_hd__buf_2
XFILLER_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20058_ _20010_/A _20058_/B _20058_/C vssd1 vssd1 vccd1 vccd1 _20058_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_86_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21445__C _21445_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22899__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _11900_/A _11900_/B vssd1 vssd1 vccd1 vccd1 _11900_/Y sky130_fd_sc_hd__nand2_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _12868_/A _12873_/A _12875_/X _12879_/Y vssd1 vssd1 vccd1 vccd1 _12880_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_172_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20592__B2 _12928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11837_/B _11833_/A _11831_/C vssd1 vssd1 vccd1 vccd1 _11831_/Y sky130_fd_sc_hd__nand3_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18537__A1 _12157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18537__B2 _11563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14863_/C _22876_/Q vssd1 vssd1 vccd1 vccd1 _14551_/A sky130_fd_sc_hd__xnor2_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11762_/A _11762_/B _11932_/C vssd1 vssd1 vccd1 vccd1 _11762_/X sky130_fd_sc_hd__and3_1
XFILLER_42_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20358__A _20358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ _13501_/A _13550_/C _13550_/A vssd1 vssd1 vccd1 vccd1 _13559_/A sky130_fd_sc_hd__nand3_1
XFILLER_92_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _22763_/Q vssd1 vssd1 vccd1 vccd1 _14775_/C sky130_fd_sc_hd__clkinv_2
XFILLER_42_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14023__A1 _22873_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11561_/X _11563_/X _11566_/X vssd1 vssd1 vccd1 vccd1 _11693_/X sky130_fd_sc_hd__a21o_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _16473_/A _17129_/B _16947_/A vssd1 vssd1 vccd1 vccd1 _16476_/A sky130_fd_sc_hd__nand3_1
X_13432_ _13635_/A _21177_/A _13192_/B _13572_/A _21848_/B vssd1 vssd1 vccd1 vccd1
+ _13433_/D sky130_fd_sc_hd__a32o_1
XANTENNA__22097__A1 _21841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15771__A1 _15350_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15771__B2 _15389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16151_ _12065_/A _13024_/A _16153_/A _17006_/D vssd1 vssd1 vccd1 vccd1 _16151_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20647__A2 _20452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13363_ _13421_/A _21367_/C vssd1 vssd1 vccd1 vccd1 _21177_/D sky130_fd_sc_hd__and2_1
XFILLER_42_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16571__A _22702_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19585__C _19602_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15102_ _15101_/A _14987_/C _15101_/B vssd1 vssd1 vccd1 vccd1 _15103_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12307__C _20461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ _12447_/A _16256_/D _12802_/C vssd1 vssd1 vccd1 vccd1 _12314_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__17386__B _17386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16082_ _16082_/A _16082_/B vssd1 vssd1 vccd1 vccd1 _16082_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13294_ _22729_/Q _22728_/Q vssd1 vssd1 vccd1 vccd1 _21188_/A sky130_fd_sc_hd__or2_1
XFILLER_181_152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19910_ _19851_/B _19909_/X _19907_/Y vssd1 vssd1 vccd1 vccd1 _19991_/A sky130_fd_sc_hd__a21o_1
XFILLER_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15033_ _15033_/A _15033_/B vssd1 vssd1 vccd1 vccd1 _15034_/B sky130_fd_sc_hd__nor2_1
X_12245_ _12245_/A _12245_/B _12245_/C vssd1 vssd1 vccd1 vccd1 _18272_/A sky130_fd_sc_hd__nand3_2
XANTENNA__19265__A2 _11351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater127_A _22877_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__C1 _19061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17276__A1 _16944_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19841_ _19842_/B _19842_/C _19176_/X _17927_/A vssd1 vssd1 vccd1 vccd1 _19909_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_122_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12176_ _12173_/Y _12174_/X _18162_/A _18165_/A vssd1 vssd1 vccd1 vccd1 _12177_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_96_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22512__S _22512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16984_ _16908_/X _16909_/X _16982_/Y _16983_/X vssd1 vssd1 vccd1 vccd1 _17027_/A
+ sky130_fd_sc_hd__o211ai_2
X_19772_ _19900_/A _19772_/B _19772_/C _19772_/D vssd1 vssd1 vccd1 vccd1 _19848_/A
+ sky130_fd_sc_hd__nand4_4
XANTENNA__19017__A2 _19176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17833__C _17833_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18225__B1 _12221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18723_ _18723_/A _18723_/B _18723_/C vssd1 vssd1 vccd1 vccd1 _18724_/A sky130_fd_sc_hd__nand3_1
X_15935_ _15935_/A vssd1 vssd1 vccd1 vccd1 _15935_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__18648__D _18648_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_884 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18654_ _18654_/A _18654_/B _18654_/C vssd1 vssd1 vccd1 vccd1 _18670_/A sky130_fd_sc_hd__nand3_1
XFILLER_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _17385_/B vssd1 vssd1 vccd1 vccd1 _20806_/C sky130_fd_sc_hd__buf_4
XANTENNA__20583__A1 _12968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17605_ _17605_/A _17605_/B vssd1 vssd1 vccd1 vccd1 _17611_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14817_ _14727_/B _14726_/C _14816_/Y vssd1 vssd1 vccd1 vccd1 _14821_/A sky130_fd_sc_hd__a21oi_1
X_18585_ _18427_/X _18428_/Y _18773_/A _18274_/Y vssd1 vssd1 vccd1 vccd1 _18586_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ _15797_/A vssd1 vssd1 vccd1 vccd1 _15797_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_149_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17536_ _17401_/Y _17532_/Y _17533_/X _17535_/Y vssd1 vssd1 vccd1 vccd1 _17536_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18664__C _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14748_ _14750_/A _14750_/B _14836_/A _14749_/B vssd1 vssd1 vccd1 vccd1 _14839_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17467_ _17467_/A vssd1 vssd1 vccd1 vccd1 _17467_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_189_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14679_ _14868_/C vssd1 vssd1 vccd1 vccd1 _14934_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14014__A1 _13904_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19206_ _19211_/A _19418_/B _19211_/C vssd1 vssd1 vccd1 vccd1 _19206_/Y sky130_fd_sc_hd__a21oi_1
X_16418_ _16418_/A _16418_/B vssd1 vssd1 vccd1 vccd1 _16419_/C sky130_fd_sc_hd__nand2_1
XFILLER_73_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17398_ _17252_/Y _17535_/A _17643_/A _17394_/Y _19768_/C vssd1 vssd1 vccd1 vccd1
+ _17399_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19137_ _19137_/A _19301_/D _19137_/C vssd1 vssd1 vccd1 vccd1 _19141_/B sky130_fd_sc_hd__nand3_1
XANTENNA__20638__A2 _12607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11402__B _11503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16349_ _20357_/A vssd1 vssd1 vccd1 vccd1 _20582_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19068_ _19074_/A _19074_/B _19066_/Y _19067_/X vssd1 vssd1 vccd1 vccd1 _19149_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15514__B2 _15707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18019_ _17953_/B _17953_/A _17957_/A vssd1 vssd1 vccd1 vccd1 _18019_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_133_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19792__A _19792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12879__A2 _20870_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12514__A _22823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21030_ _21030_/A _21030_/B _21030_/C vssd1 vssd1 vccd1 vccd1 _21031_/B sky130_fd_sc_hd__or3_1
XFILLER_99_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16490__A2 _12774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21932_ _21917_/A _21917_/B _21836_/A vssd1 vssd1 vccd1 vccd1 _21932_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_27_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20574__B2 _20449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21863_ _21861_/X _21726_/Y _21633_/B _21862_/X vssd1 vssd1 vccd1 vccd1 _21865_/C
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20326__A1 _12577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20814_ _20813_/X _20810_/B _20810_/A _20812_/A _20812_/B vssd1 vssd1 vccd1 vccd1
+ _20816_/A sky130_fd_sc_hd__a32oi_2
X_21794_ _21664_/X _21671_/Y _21793_/Y vssd1 vssd1 vccd1 vccd1 _21794_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_196_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20178__A _20178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20745_ _20745_/A _21017_/C _20745_/C vssd1 vssd1 vccd1 vccd1 _20745_/X sky130_fd_sc_hd__and3_1
XFILLER_168_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20676_ _20676_/A _20676_/B vssd1 vssd1 vccd1 vccd1 _20676_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22393__A _22439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22415_ _22426_/A vssd1 vssd1 vccd1 vccd1 _22424_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16822__C _16822_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15505__A1 _12930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22346_ _22346_/A _22346_/B vssd1 vssd1 vccd1 vccd1 _22943_/D sky130_fd_sc_hd__xor2_1
XANTENNA__15505__B2 _12111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22277_ _22277_/A _22277_/B vssd1 vssd1 vccd1 vccd1 _22277_/X sky130_fd_sc_hd__and2_1
XFILLER_117_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15438__C _16488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17258__A1 _12294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ _12054_/A _12054_/B vssd1 vssd1 vccd1 vccd1 _12088_/B sky130_fd_sc_hd__nand2_2
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17258__B2 _15541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21228_ _21226_/Y _21227_/X _21238_/C _21238_/B vssd1 vssd1 vccd1 vccd1 _21230_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_151_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21159_ _22948_/Q _21165_/A vssd1 vssd1 vccd1 vccd1 _21164_/A sky130_fd_sc_hd__nor2_1
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13981_ _14122_/A _14073_/A _13986_/A _13884_/X _13883_/Y vssd1 vssd1 vccd1 vccd1
+ _13992_/A sky130_fd_sc_hd__o32a_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15720_ _15911_/A vssd1 vssd1 vccd1 vccd1 _15960_/A sky130_fd_sc_hd__buf_4
XFILLER_37_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_832 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12932_ _12933_/A _12933_/B _12927_/X _12931_/X vssd1 vssd1 vccd1 vccd1 _12957_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16233__A2 _16227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _15329_/X _15319_/B _15321_/Y vssd1 vssd1 vccd1 vccd1 _15651_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12863_ _12863_/A _12863_/B vssd1 vssd1 vccd1 vccd1 _12864_/B sky130_fd_sc_hd__nor2_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13047__A2 _12894_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14602_/A _14602_/B _14602_/C vssd1 vssd1 vccd1 vccd1 _14602_/Y sky130_fd_sc_hd__nand3_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _11542_/A _16276_/A _18092_/Y _17427_/A _12116_/A vssd1 vssd1 vccd1 vccd1
+ _18370_/X sky130_fd_sc_hd__o32a_1
X_11814_ _11814_/A _11814_/B vssd1 vssd1 vccd1 vccd1 _11930_/C sky130_fd_sc_hd__nand2_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15582_ _15579_/X _15581_/X _15571_/Y _15566_/X vssd1 vssd1 vccd1 vccd1 _15583_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__15992__A1 _15649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15901__C _15901_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _20123_/A _12704_/A _12844_/A _12793_/X _12788_/C vssd1 vssd1 vccd1 vccd1
+ _12794_/X sky130_fd_sc_hd__o311a_1
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17321_ _17311_/X _17127_/A _17323_/C vssd1 vssd1 vccd1 vccd1 _17324_/B sky130_fd_sc_hd__o21bai_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14561_/D _14561_/B _22875_/Q _14273_/C vssd1 vssd1 vccd1 vccd1 _14541_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_11745_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11745_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11503__A _11503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17252_ _16225_/X _16227_/X _20129_/A _17401_/D vssd1 vssd1 vccd1 vccd1 _17252_/Y
+ sky130_fd_sc_hd__o211ai_4
X_14464_ _14461_/Y _14462_/Y _14463_/X vssd1 vssd1 vccd1 vccd1 _14472_/A sky130_fd_sc_hd__o21bai_1
XFILLER_169_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11676_ _11668_/A _16482_/A _15435_/C vssd1 vssd1 vccd1 vccd1 _11706_/A sky130_fd_sc_hd__a21o_1
XFILLER_169_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16203_ _16421_/C _16418_/A _16418_/B vssd1 vssd1 vccd1 vccd1 _16203_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__22914__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17397__A _19687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13415_ _21268_/A _21259_/B _21259_/C _21270_/C _21270_/A vssd1 vssd1 vccd1 vccd1
+ _13416_/B sky130_fd_sc_hd__o32a_1
XFILLER_179_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17183_ _16982_/A _17105_/Y _17188_/B vssd1 vssd1 vccd1 vccd1 _17184_/C sky130_fd_sc_hd__o21ai_1
XFILLER_127_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14395_ _22771_/Q _14322_/X _14379_/X _22739_/Q _14394_/X vssd1 vssd1 vccd1 vccd1
+ _14395_/X sky130_fd_sc_hd__a221o_1
XFILLER_167_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16134_ _16134_/A _16134_/B vssd1 vssd1 vccd1 vccd1 _16137_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13346_ _13344_/X _13345_/X _13326_/Y vssd1 vssd1 vccd1 vccd1 _13346_/X sky130_fd_sc_hd__a21o_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13770__A3 _14181_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16065_ _18130_/C vssd1 vssd1 vccd1 vccd1 _19470_/D sky130_fd_sc_hd__buf_4
XFILLER_185_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13277_ _13210_/B _13210_/C _13210_/A vssd1 vssd1 vccd1 vccd1 _13282_/B sky130_fd_sc_hd__a21boi_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17249__A1 _12696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15016_ _15015_/B _15015_/C _15015_/A vssd1 vssd1 vccd1 vccd1 _15017_/B sky130_fd_sc_hd__a21oi_1
X_12228_ _12039_/B _12039_/C _12039_/A _12029_/Y _12081_/Y vssd1 vssd1 vccd1 vccd1
+ _12231_/A sky130_fd_sc_hd__a32oi_2
XFILLER_64_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18997__A1 _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18997__B2 _15887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12730__A1 _12602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19824_ _19293_/X _19294_/X _19761_/Y _19881_/B _19818_/B vssd1 vssd1 vccd1 vccd1
+ _19892_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_151_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18659__C _19507_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12159_ _12157_/X _12158_/X _15377_/A vssd1 vssd1 vccd1 vccd1 _12162_/A sky130_fd_sc_hd__a21oi_2
XFILLER_110_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_648 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12988__B _12988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16472__A2 _18797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__B _19455_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19755_ _20025_/A _19749_/X _19752_/Y _22920_/Q vssd1 vssd1 vccd1 vccd1 _19827_/B
+ sky130_fd_sc_hd__o211ai_1
X_16967_ _16967_/A _16967_/B _16967_/C vssd1 vssd1 vccd1 vccd1 _16978_/A sky130_fd_sc_hd__nand3_1
XFILLER_65_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18706_ _18706_/A _18706_/B _18999_/A vssd1 vssd1 vccd1 vccd1 _18707_/B sky130_fd_sc_hd__and3_1
XFILLER_83_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15918_ _15918_/A vssd1 vssd1 vccd1 vccd1 _15918_/X sky130_fd_sc_hd__buf_2
XANTENNA__20556__A1 _20548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16898_ _17502_/A _16660_/Y _17215_/B _17215_/C _17064_/C vssd1 vssd1 vccd1 vccd1
+ _16899_/C sky130_fd_sc_hd__o2111ai_2
X_19686_ _19350_/X _17647_/A _17391_/A _18718_/X vssd1 vssd1 vccd1 vccd1 _19689_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_65_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18637_ _18778_/B _17400_/X _18626_/Y _18629_/Y _18953_/A vssd1 vssd1 vccd1 vccd1
+ _18637_/X sky130_fd_sc_hd__o311a_1
X_15849_ _15849_/A vssd1 vssd1 vccd1 vccd1 _15970_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15380__A _15415_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18568_ _18568_/A _18568_/B _18568_/C vssd1 vssd1 vccd1 vccd1 _18569_/C sky130_fd_sc_hd__nand3_1
XANTENNA__15983__A1 _11904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14708__B _14857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1112 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17519_ _17054_/Y _17078_/Y _17518_/Y vssd1 vssd1 vccd1 vccd1 _17519_/Y sky130_fd_sc_hd__a21oi_1
X_18499_ _18499_/A _18499_/B _18499_/C vssd1 vssd1 vccd1 vccd1 _18526_/D sky130_fd_sc_hd__nand3_2
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18691__A _18691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20530_ _20532_/A _20532_/B _20568_/A _20534_/A vssd1 vssd1 vccd1 vccd1 _20531_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_138_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21808__A1 _21805_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20461_ _20461_/A _20461_/B _20461_/C vssd1 vssd1 vccd1 vccd1 _20462_/A sky130_fd_sc_hd__nand3_4
XFILLER_192_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19477__A2 _19839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22200_ _21908_/X _21911_/X _22024_/Y _22160_/Y vssd1 vssd1 vccd1 vccd1 _22200_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_146_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20392_ _12500_/X _12501_/X _22827_/Q vssd1 vssd1 vccd1 vccd1 _20393_/C sky130_fd_sc_hd__o21ai_2
XFILLER_173_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22131_ _22131_/A _22131_/B vssd1 vssd1 vccd1 vccd1 _22132_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22660__B _22660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22062_ _22062_/A _22262_/A _22190_/D vssd1 vssd1 vccd1 vccd1 _22113_/A sky130_fd_sc_hd__and3_1
XFILLER_88_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21013_ _21083_/C _20972_/A _21081_/C _21012_/X vssd1 vssd1 vccd1 vccd1 _21013_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11524__A2 _18116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20795__A1 _20792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21339__A3 _21498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22964_ _22964_/CLK _22964_/D vssd1 vssd1 vccd1 vccd1 _22964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17412__A1 _12234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17412__B2 _15355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21915_ _21908_/X _21911_/X _22024_/A vssd1 vssd1 vccd1 vccd1 _21915_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_16_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22895_ _22952_/CLK _22895_/D vssd1 vssd1 vccd1 vccd1 _22895_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_167_1034 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17963__A2 _17227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15974__A1 _15504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21846_ _21846_/A _21846_/B _21846_/C _21846_/D vssd1 vssd1 vccd1 vccd1 _21847_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_169_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15721__C _15960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22937__CLK _22937_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21777_ _21841_/C _21777_/B vssd1 vssd1 vccd1 vccd1 _21790_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11530_ _11578_/A _11581_/A _11529_/Y vssd1 vssd1 vccd1 vccd1 _11533_/A sky130_fd_sc_hd__o21ai_1
XFILLER_169_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15726__A1 _15723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20728_ _20728_/A _20728_/B _20728_/C _20818_/A vssd1 vssd1 vccd1 vccd1 _20818_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_196_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17929__B _21011_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11461_ _12090_/C vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19468__A2 _19839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20659_ _20656_/B _20656_/C _20656_/A vssd1 vssd1 vccd1 vccd1 _20659_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_104_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _21473_/A vssd1 vssd1 vccd1 vccd1 _21185_/A sky130_fd_sc_hd__buf_2
XFILLER_125_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11392_ _11502_/A _11503_/A _18984_/A _18984_/B vssd1 vssd1 vccd1 vccd1 _11392_/Y
+ sky130_fd_sc_hd__o211ai_2
X_14180_ _14180_/A _14180_/B _14180_/C vssd1 vssd1 vccd1 vccd1 _14180_/Y sky130_fd_sc_hd__nand3_1
XFILLER_180_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20483__B1 _20593_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _22725_/Q vssd1 vssd1 vccd1 vccd1 _13131_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16151__A1 _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22329_ _21473_/Y _21579_/A _22306_/B _22055_/Y _22306_/C vssd1 vssd1 vccd1 vccd1
+ _22329_/Y sky130_fd_sc_hd__a2111oi_4
XFILLER_180_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16151__B2 _17006_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input55_A wb_dat_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ _22735_/Q vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_180_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12712__A1 _12689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12013_ _12013_/A _12013_/B _12013_/C vssd1 vssd1 vccd1 vccd1 _12013_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__11993__A _22792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17870_ _17785_/X _17954_/B _17860_/B _17860_/A vssd1 vssd1 vccd1 vccd1 _17907_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_120_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16821_ _16014_/A _15939_/A _16810_/C _16810_/D vssd1 vssd1 vccd1 vccd1 _16822_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_120_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_bq_clk_i clkbuf_4_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _22916_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_87_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19540_ _19540_/A _19540_/B _19540_/C vssd1 vssd1 vccd1 vccd1 _19540_/Y sky130_fd_sc_hd__nand3_2
X_16752_ _16598_/A _16598_/B _16599_/C _16599_/B vssd1 vssd1 vccd1 vccd1 _16753_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_98_1120 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13964_ _14583_/C _14583_/D _13849_/C vssd1 vssd1 vccd1 vccd1 _13973_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12476__B1 _12493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15703_ _15703_/A _15703_/B vssd1 vssd1 vccd1 vccd1 _15704_/B sky130_fd_sc_hd__nand2_1
X_12915_ _12602_/Y _12613_/Y _12916_/A _12916_/B _12601_/Y vssd1 vssd1 vccd1 vccd1
+ _12915_/Y sky130_fd_sc_hd__o221ai_1
XANTENNA__19943__A3 _19461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16683_ _16664_/A _16683_/B _16683_/C _17065_/A vssd1 vssd1 vccd1 vccd1 _16685_/B
+ sky130_fd_sc_hd__nand4b_1
X_19471_ _19476_/A _19476_/B _19476_/C vssd1 vssd1 vccd1 vccd1 _19479_/C sky130_fd_sc_hd__nand3_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13895_ _13820_/A _14583_/C _13963_/C _14383_/A vssd1 vssd1 vccd1 vccd1 _13899_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_185_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18422_ _18216_/B _18216_/A _18417_/C _18417_/A vssd1 vssd1 vccd1 vccd1 _18423_/C
+ sky130_fd_sc_hd__o211ai_1
X_15634_ _18512_/A _15718_/A _15638_/A vssd1 vssd1 vccd1 vccd1 _15634_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13713__A _14165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12846_ _17144_/A vssd1 vssd1 vccd1 vccd1 _20129_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _18354_/A _18354_/B _18726_/A _18520_/B vssd1 vssd1 vccd1 vccd1 _18353_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20249__C _20249_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15565_ _15567_/A _15565_/B _15565_/C _15565_/D vssd1 vssd1 vccd1 vccd1 _15566_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12765_/X _20177_/A _12886_/B _12776_/X vssd1 vssd1 vccd1 vccd1 _12777_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17304_/A _17304_/B vssd1 vssd1 vccd1 vccd1 _17475_/A sky130_fd_sc_hd__nand2_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14505_/X _14516_/B _14516_/C vssd1 vssd1 vccd1 vccd1 _14522_/C sky130_fd_sc_hd__nand3b_2
X_18284_ _12204_/X _17388_/A _18296_/A vssd1 vssd1 vccd1 vccd1 _18291_/A sky130_fd_sc_hd__o21ai_1
X_11728_ _11941_/A vssd1 vssd1 vccd1 vccd1 _16256_/B sky130_fd_sc_hd__buf_4
XANTENNA__15717__A1 _17128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13151__C _21609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_743 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17839__B _17839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15496_ _11721_/C _14439_/A _16226_/C _15495_/X vssd1 vssd1 vccd1 vccd1 _15523_/A
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__16914__B1 _15690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17235_ _18200_/A _19351_/C _20870_/A _20870_/B vssd1 vssd1 vccd1 vccd1 _17235_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_147_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14447_ _16226_/B _14439_/A _22967_/Q _16242_/B _18259_/B vssd1 vssd1 vccd1 vccd1
+ _14448_/A sky130_fd_sc_hd__o41a_2
X_11659_ _11712_/A _11659_/B _15482_/B _11659_/D vssd1 vssd1 vccd1 vccd1 _11660_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_122_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17166_ _16932_/Y _17133_/Y _17288_/A _17385_/B _19772_/D vssd1 vssd1 vccd1 vccd1
+ _17169_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14378_ _16324_/C vssd1 vssd1 vccd1 vccd1 _20069_/A sky130_fd_sc_hd__buf_4
XFILLER_183_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16117_ _16115_/X _16082_/Y _16169_/B vssd1 vssd1 vccd1 vccd1 _16118_/C sky130_fd_sc_hd__o21ai_2
XFILLER_31_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20474__B1 _20579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13329_ _13337_/A vssd1 vssd1 vccd1 vccd1 _13329_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17097_ _17341_/A _17310_/A _17341_/C _17341_/D vssd1 vssd1 vccd1 vccd1 _17103_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12064__A _12064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16048_ _17539_/D vssd1 vssd1 vccd1 vccd1 _20745_/C sky130_fd_sc_hd__buf_4
XFILLER_131_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17574__B _17574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22911__D _22911_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19807_ _19807_/A _19807_/B vssd1 vssd1 vccd1 vccd1 _19809_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__16445__A2 _15630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14456__A1 _11667_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17999_ _17999_/A vssd1 vssd1 vccd1 vccd1 _17999_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11408__A _22956_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19738_ _19742_/B _19808_/A _19742_/A vssd1 vssd1 vccd1 vccd1 _19746_/A sky130_fd_sc_hd__a21o_1
XFILLER_37_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18198__A2 _19353_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19669_ _19669_/A _19669_/B vssd1 vssd1 vccd1 vccd1 _19669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_610 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21700_ _21700_/A vssd1 vssd1 vccd1 vccd1 _21700_/X sky130_fd_sc_hd__buf_2
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22680_ _22943_/CLK _22680_/D vssd1 vssd1 vccd1 vccd1 _22680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19013__C _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21631_ _21631_/A _21638_/A vssd1 vssd1 vccd1 vccd1 _21635_/C sky130_fd_sc_hd__nand2_1
XFILLER_52_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15708__A1 _15397_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21562_ _21423_/Y _21561_/Y _21426_/Y vssd1 vssd1 vccd1 vccd1 _21562_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_178_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20513_ _20323_/Y _20328_/D _20512_/Y vssd1 vssd1 vccd1 vccd1 _20513_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_166_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15184__A2 _15056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21493_ _21725_/A _21725_/B _21741_/B vssd1 vssd1 vccd1 vccd1 _21493_/Y sky130_fd_sc_hd__nand3_1
XFILLER_193_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20444_ _20444_/A _20444_/B vssd1 vssd1 vccd1 vccd1 _20754_/B sky130_fd_sc_hd__nor2_2
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19855__C1 _19795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12942__A1 _15774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18393__A2_N _18407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20375_ _20375_/A _20375_/B _20375_/C vssd1 vssd1 vccd1 vccd1 _20376_/A sky130_fd_sc_hd__nand3_1
XFILLER_107_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22114_ _22113_/B _22113_/C _21939_/A _22119_/A vssd1 vssd1 vccd1 vccd1 _22115_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__21287__A _21423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15892__B1 _11504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22045_ _22045_/A _22045_/B vssd1 vssd1 vccd1 vccd1 _22045_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12702__A _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19622__A2 _18107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13517__B _21480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15435__D _15435_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11318__A _18690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22947_ _22948_/CLK _22947_/D vssd1 vssd1 vccd1 vccd1 _22947_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_515 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12700_ _15774_/C _20579_/C vssd1 vssd1 vccd1 vccd1 _12700_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13680_ _13558_/C _13557_/X _13612_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 _13680_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_71_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22878_ _22944_/CLK input72/X vssd1 vssd1 vccd1 vccd1 _22878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_356 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ _16488_/A vssd1 vssd1 vccd1 vccd1 _15901_/C sky130_fd_sc_hd__buf_2
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21829_ _21568_/A _21827_/Y _21706_/A _21828_/Y vssd1 vssd1 vccd1 vccd1 _21832_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15350_ _16302_/A _20605_/B _18876_/C vssd1 vssd1 vccd1 vccd1 _15350_/Y sky130_fd_sc_hd__nand3_4
XFILLER_141_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12562_ _12546_/A _12769_/A _12645_/C vssd1 vssd1 vccd1 vccd1 _12562_/X sky130_fd_sc_hd__a21o_1
XFILLER_196_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14301_ input9/X input8/X input11/X input10/X vssd1 vssd1 vccd1 vccd1 _14302_/C sky130_fd_sc_hd__or4_1
XFILLER_169_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11513_ _11511_/X _18203_/B _11493_/Y _11501_/Y vssd1 vssd1 vccd1 vccd1 _11551_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_156_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15281_ _15287_/D _15271_/B _22881_/Q vssd1 vssd1 vccd1 vccd1 _15282_/B sky130_fd_sc_hd__a21oi_1
XFILLER_141_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12493_ _12493_/A _12520_/B vssd1 vssd1 vccd1 vccd1 _12493_/Y sky130_fd_sc_hd__nand2_4
X_17020_ _17020_/A _17027_/C vssd1 vssd1 vccd1 vccd1 _17020_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14232_ _15050_/B _14231_/A _14231_/B _14231_/C vssd1 vssd1 vccd1 vccd1 _14233_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18649__B1 _17421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11444_ _19061_/A _18288_/A _16711_/C _15912_/C vssd1 vssd1 vccd1 vccd1 _11444_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__22445__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17097__D _17341_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19310__A1 _16711_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11736__A2 _11503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18113__A2 _18278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19310__B2 _19470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11500__B _18131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ _14163_/A _14163_/B _14163_/C vssd1 vssd1 vccd1 vccd1 _14248_/B sky130_fd_sc_hd__nand3_2
X_11375_ _11421_/A vssd1 vssd1 vccd1 vccd1 _11980_/B sky130_fd_sc_hd__buf_2
XFILLER_113_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_0_0_bq_clk_i_A clkbuf_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13114_ _13344_/A _13345_/A vssd1 vssd1 vccd1 vccd1 _13513_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14135__B1 _13748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18971_ _18788_/A _18969_/X _18970_/Y vssd1 vssd1 vccd1 vccd1 _18972_/B sky130_fd_sc_hd__o21ai_1
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15907__B _16781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14094_ _14094_/A _14094_/B _14094_/C vssd1 vssd1 vccd1 vccd1 _14178_/C sky130_fd_sc_hd__nand3_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21628__C _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17922_ _17922_/A vssd1 vssd1 vccd1 vccd1 _21082_/C sky130_fd_sc_hd__buf_2
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13045_/A _13045_/B _20304_/A vssd1 vssd1 vccd1 vccd1 _13045_/Y sky130_fd_sc_hd__nand3_4
XFILLER_26_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16427__A2 _16402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17853_ _17853_/A _17853_/B vssd1 vssd1 vccd1 vccd1 _17910_/C sky130_fd_sc_hd__nor2_1
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18821__B1 _18666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12331__B _16256_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16804_ _16972_/A _16971_/A _16971_/B vssd1 vssd1 vccd1 vccd1 _16908_/C sky130_fd_sc_hd__nand3_1
XANTENNA__15923__A _16011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17784_ _17855_/A _17855_/B _17778_/A vssd1 vssd1 vccd1 vccd1 _17784_/Y sky130_fd_sc_hd__o21ai_1
X_14996_ _14934_/Y _14996_/B _14996_/C _14996_/D vssd1 vssd1 vccd1 vccd1 _15001_/C
+ sky130_fd_sc_hd__nand4b_2
XANTENNA__12050__C _19490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19523_ _19536_/A _19536_/B _19523_/C _19523_/D vssd1 vssd1 vccd1 vccd1 _19528_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16735_ _11821_/X _15935_/A _16466_/X _16261_/Y _16842_/B vssd1 vssd1 vccd1 vccd1
+ _16735_/X sky130_fd_sc_hd__o311a_2
X_13947_ _13947_/A _13947_/B _13947_/C vssd1 vssd1 vccd1 vccd1 _13957_/C sky130_fd_sc_hd__nand3_1
XANTENNA__21184__A1 _13050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19454_ _19651_/A _19896_/A _19454_/C _19602_/C vssd1 vssd1 vccd1 vccd1 _19454_/X
+ sky130_fd_sc_hd__and4_2
X_16666_ _16669_/A _16670_/A vssd1 vssd1 vccd1 vccd1 _16667_/A sky130_fd_sc_hd__or2_1
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13878_ _13984_/A vssd1 vssd1 vccd1 vccd1 _14889_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__20931__A1 _20806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18405_ _18177_/X _18178_/Y _18163_/Y vssd1 vssd1 vccd1 vccd1 _18405_/X sky130_fd_sc_hd__o21a_1
X_15617_ _15617_/A vssd1 vssd1 vccd1 vccd1 _15617_/X sky130_fd_sc_hd__buf_4
XFILLER_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13162__B _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ _12396_/A _12823_/A _12324_/X vssd1 vssd1 vccd1 vccd1 _15370_/A sky130_fd_sc_hd__o21ai_4
X_19385_ _19240_/C _19240_/D _19343_/A vssd1 vssd1 vccd1 vccd1 _19385_/Y sky130_fd_sc_hd__a21boi_1
X_16597_ _16599_/C _16599_/B _16598_/A _16598_/B vssd1 vssd1 vccd1 vccd1 _16602_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_50_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19768__C _19768_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15548_ _15548_/A _15548_/B vssd1 vssd1 vccd1 vccd1 _16964_/A sky130_fd_sc_hd__nand2_2
X_18336_ _18137_/Y _18139_/X _18141_/Y _18150_/B vssd1 vssd1 vccd1 vccd1 _18345_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__18888__B1 _18128_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16473__B _16473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18267_ _18088_/Y _18252_/Y _18262_/Y _18266_/A vssd1 vssd1 vccd1 vccd1 _18268_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15479_ _15479_/A _15479_/B _15479_/C vssd1 vssd1 vccd1 vccd1 _15502_/D sky130_fd_sc_hd__nand3_2
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16192__C _17401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17218_ _17371_/A _17371_/B _17370_/A _17373_/A _17370_/B vssd1 vssd1 vccd1 vccd1
+ _17219_/B sky130_fd_sc_hd__o2111a_1
X_18198_ _12050_/B _19353_/B _19353_/C _18195_/Y _18197_/Y vssd1 vssd1 vccd1 vccd1
+ _18571_/B sky130_fd_sc_hd__a32o_2
XFILLER_128_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18104__A2 _16711_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17149_ _17149_/A _17149_/B vssd1 vssd1 vccd1 vccd1 _17149_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16115__A1 _16053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20160_ _20167_/A _20167_/B vssd1 vssd1 vccd1 vccd1 _20162_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14721__B _14721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14677__B2 _14057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20091_ _12803_/X _20214_/A _20090_/Y vssd1 vssd1 vccd1 vccd1 _20093_/A sky130_fd_sc_hd__o21ai_1
XFILLER_130_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12522__A _12522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_919 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22801_ _22801_/CLK _22801_/D vssd1 vssd1 vccd1 vccd1 _22801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22369__C input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22372__A0 _12876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20993_ _21062_/A vssd1 vssd1 vccd1 vccd1 _21006_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13652__A2 _21195_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15390__A2_N _15665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22732_ _22733_/CLK _22732_/D vssd1 vssd1 vccd1 vccd1 _22732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22663_ _22663_/A vssd1 vssd1 vccd1 vccd1 _22951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21614_ _21614_/A vssd1 vssd1 vccd1 vccd1 _21730_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20186__A _20314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22594_ _22594_/A vssd1 vssd1 vccd1 vccd1 _22786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21545_ _21545_/A _21545_/B _21545_/C vssd1 vssd1 vccd1 vccd1 _21546_/B sky130_fd_sc_hd__nand3_1
XANTENNA__15562__C1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19694__B _19694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21476_ _21476_/A _21749_/A _21476_/C vssd1 vssd1 vccd1 vccd1 _21596_/A sky130_fd_sc_hd__nand3_2
XFILLER_119_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20914__A _21019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12915__A1 _12602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20427_ _20427_/A _20427_/B vssd1 vssd1 vccd1 vccd1 _20427_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15727__B _15727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20358_ _20358_/A _20358_/B vssd1 vssd1 vccd1 vccd1 _20368_/A sky130_fd_sc_hd__nand2_1
XFILLER_161_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17645__D _17645_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19056__B1 _17632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20521__A1_N _20337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20289_ _20198_/Y _20158_/B _20167_/B _20200_/X vssd1 vssd1 vccd1 vccd1 _20290_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22028_ _21986_/B _21986_/C _21841_/A _21220_/X vssd1 vssd1 vccd1 vccd1 _22075_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15880__A3 _16402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14850_ _14832_/X _14829_/X _14828_/Y vssd1 vssd1 vccd1 vccd1 _14923_/B sky130_fd_sc_hd__a21bo_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17648__A1_N _17645_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13801_ _13897_/A _13833_/B _13833_/C _13869_/C vssd1 vssd1 vccd1 vccd1 _13974_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_75_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input18_A wb_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14781_ _14781_/A _14857_/A _14948_/C _14895_/A vssd1 vssd1 vccd1 vccd1 _14895_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_95_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11993_ _22792_/Q vssd1 vssd1 vccd1 vccd1 _18313_/A sky130_fd_sc_hd__inv_2
XFILLER_91_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16520_ _16520_/A vssd1 vssd1 vccd1 vccd1 _16534_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13732_ _13798_/A _13733_/B vssd1 vssd1 vccd1 vccd1 _13869_/B sky130_fd_sc_hd__nand2_2
XFILLER_45_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16451_ _16451_/A _16451_/B vssd1 vssd1 vccd1 vccd1 _16734_/B sky130_fd_sc_hd__nand2_1
X_13663_ _13663_/A _13663_/B vssd1 vssd1 vccd1 vccd1 _13665_/B sky130_fd_sc_hd__or2_1
XFILLER_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15402_ _12094_/D _15394_/A _12598_/A _18512_/A vssd1 vssd1 vccd1 vccd1 _15403_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _12584_/Y _12601_/Y _12602_/Y _12613_/Y vssd1 vssd1 vccd1 vccd1 _12618_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_19170_ _17421_/X _17422_/X _12108_/A _12108_/B vssd1 vssd1 vccd1 vccd1 _19170_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _15673_/A _15673_/C _16372_/X vssd1 vssd1 vccd1 vccd1 _16636_/B sky130_fd_sc_hd__a21o_1
X_13594_ _21250_/A _21750_/C _21250_/C vssd1 vssd1 vccd1 vccd1 _13663_/A sky130_fd_sc_hd__and3_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18334__A2 _11786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18121_ _11377_/A _18116_/D _18677_/B _18128_/A vssd1 vssd1 vccd1 vccd1 _18483_/B
+ sky130_fd_sc_hd__o211ai_4
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11957__A2 _11503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15333_ _12576_/X _12577_/X _17532_/A _11627_/A vssd1 vssd1 vccd1 vccd1 _15333_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_40_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20677__B1 _20913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16724__D _20593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12545_ _12543_/B _12543_/C _12543_/D _12469_/A vssd1 vssd1 vccd1 vccd1 _12546_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20141__A2 _12696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18052_ _18069_/C _18051_/C _18051_/A vssd1 vssd1 vccd1 vccd1 _18077_/A sky130_fd_sc_hd__a21o_1
XFILLER_145_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11511__A _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15264_ _15176_/A _15260_/B _15262_/B _15262_/A vssd1 vssd1 vccd1 vccd1 _22816_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_126_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12476_ _12335_/A _12403_/A _12493_/A vssd1 vssd1 vccd1 vccd1 _12501_/A sky130_fd_sc_hd__o21a_2
XFILLER_144_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17003_ _16098_/X _17091_/A _16997_/A vssd1 vssd1 vccd1 vccd1 _17005_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11868__D _12050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14215_ _14203_/X _14185_/X _14214_/Y _14206_/Y vssd1 vssd1 vccd1 vccd1 _14215_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15918__A _15918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _11619_/B vssd1 vssd1 vccd1 vccd1 _18674_/A sky130_fd_sc_hd__buf_2
X_15195_ _15161_/A _15161_/B _15197_/B _15223_/A _15163_/X vssd1 vssd1 vccd1 vccd1
+ _15210_/B sky130_fd_sc_hd__o221a_1
XANTENNA__18637__A3 _18626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16648__A2 _21086_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _14146_/A _14146_/B _14146_/C vssd1 vssd1 vccd1 vccd1 _14147_/A sky130_fd_sc_hd__nand3_2
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ _15484_/A _11605_/A _11334_/X vssd1 vssd1 vccd1 vccd1 _11594_/A sky130_fd_sc_hd__o21a_1
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11590__B1 _18797_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18954_ _18952_/A _18952_/B _18953_/X _18627_/Y vssd1 vssd1 vccd1 vccd1 _18955_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_14077_ _14068_/X _14072_/Y _14075_/Y _14076_/Y vssd1 vssd1 vccd1 vccd1 _14147_/B
+ sky130_fd_sc_hd__o211ai_4
X_11289_ _22968_/Q vssd1 vssd1 vccd1 vccd1 _11411_/A sky130_fd_sc_hd__clkbuf_2
X_17905_ _17954_/A _17869_/A _17949_/A vssd1 vssd1 vccd1 vccd1 _17908_/B sky130_fd_sc_hd__o21a_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13028_ _13028_/A _13028_/B _13028_/C vssd1 vssd1 vccd1 vccd1 _13028_/Y sky130_fd_sc_hd__nand3_1
X_18885_ _18333_/X _18875_/Y _18880_/B _18881_/X vssd1 vssd1 vccd1 vccd1 _18887_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17836_ _17900_/B _17900_/A vssd1 vssd1 vccd1 vccd1 _17842_/A sky130_fd_sc_hd__xor2_2
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17767_ _17768_/B _17768_/C _17768_/A vssd1 vssd1 vccd1 vccd1 _17769_/A sky130_fd_sc_hd__o21ai_1
X_14979_ _14919_/C _14978_/Y _14919_/B vssd1 vssd1 vccd1 vccd1 _14980_/C sky130_fd_sc_hd__o21ai_1
X_19506_ _12170_/X _12171_/X _17532_/C _17532_/D _19651_/B vssd1 vssd1 vccd1 vccd1
+ _19506_/Y sky130_fd_sc_hd__o2111ai_2
X_16718_ _16714_/X _17087_/A _16712_/X _16710_/Y vssd1 vssd1 vccd1 vccd1 _16719_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17698_ _17579_/Y _17585_/Y _17583_/Y vssd1 vssd1 vccd1 vccd1 _17699_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__16033__B1 _16034_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19437_ _19296_/A _19434_/Y _19436_/Y vssd1 vssd1 vccd1 vccd1 _19437_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16649_ _16635_/A _16895_/B _16650_/C vssd1 vssd1 vccd1 vccd1 _16653_/A sky130_fd_sc_hd__a21o_1
XANTENNA__15387__A2 _17424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13398__A1 _13339_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19368_ _19368_/A _19368_/B vssd1 vssd1 vccd1 vccd1 _19368_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20437__C _20554_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18319_ _18319_/A _18319_/B _18319_/C vssd1 vssd1 vccd1 vccd1 _18512_/C sky130_fd_sc_hd__and3_1
XANTENNA__12070__A1 _12064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19299_ _19299_/A _19299_/B _19299_/C vssd1 vssd1 vccd1 vccd1 _19299_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__12517__A _22825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21330_ _21330_/A _21330_/B vssd1 vssd1 vccd1 vccd1 _21850_/A sky130_fd_sc_hd__nand2_2
XFILLER_176_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20734__A _20734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_1019 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21261_ _21266_/A _21261_/B _21266_/B vssd1 vssd1 vccd1 vccd1 _21261_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__18204__A _18204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16650__C _16650_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17297__C1 _17304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20212_ _15617_/A _15370_/B _20341_/C _20213_/A vssd1 vssd1 vccd1 vccd1 _20339_/A
+ sky130_fd_sc_hd__o211ai_4
X_21192_ _21192_/A vssd1 vssd1 vccd1 vccd1 _21970_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20143_ _20143_/A _20143_/B vssd1 vssd1 vccd1 vccd1 _20143_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14114__A3 _14491_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19589__A1 _12207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20074_ _12761_/X _20429_/B _12792_/Y _20073_/Y vssd1 vssd1 vccd1 vccd1 _20077_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22593__A0 _11306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16809__D _19317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12833__B1 _12519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20976_ _20917_/A _20975_/B _17806_/D _20910_/Y _20919_/B vssd1 vssd1 vccd1 vccd1
+ _20977_/C sky130_fd_sc_hd__a32o_1
XFILLER_41_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22715_ _22747_/CLK _22715_/D vssd1 vssd1 vccd1 vccd1 _22715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16394__A _20793_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22678__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13389__A1 _13339_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16825__C _17539_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22646_ _22810_/Q input53/X _22652_/S vssd1 vssd1 vccd1 vccd1 _22647_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16327__A1 _15645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22577_ _22577_/A vssd1 vssd1 vccd1 vccd1 _22779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12330_ _22818_/Q vssd1 vssd1 vccd1 vccd1 _20346_/C sky130_fd_sc_hd__buf_2
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21528_ _21393_/C _21393_/B _21387_/Y _21386_/X vssd1 vssd1 vccd1 vccd1 _21529_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_194_684 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12261_ _22688_/Q _22689_/Q vssd1 vssd1 vccd1 vccd1 _12276_/A sky130_fd_sc_hd__nor2_1
XFILLER_108_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21459_ _21216_/B _21352_/X _21349_/X vssd1 vssd1 vccd1 vccd1 _21460_/D sky130_fd_sc_hd__o21ai_1
XFILLER_147_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18114__A _18279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14000_ _13902_/A _13902_/B _14618_/A vssd1 vssd1 vccd1 vccd1 _14002_/A sky130_fd_sc_hd__a21o_1
XFILLER_141_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12364__A2 _12403_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ _12191_/X _12007_/Y _12014_/X _12088_/A _12088_/B vssd1 vssd1 vccd1 vccd1
+ _18214_/B sky130_fd_sc_hd__a32oi_4
XFILLER_1_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput86 _14374_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[13] sky130_fd_sc_hd__buf_2
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput97 _14407_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_49_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15951_ _15951_/A _16210_/A vssd1 vssd1 vccd1 vccd1 _15957_/B sky130_fd_sc_hd__nand2_1
XFILLER_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14902_ _14902_/A _14902_/B vssd1 vssd1 vccd1 vccd1 _14904_/A sky130_fd_sc_hd__nand2_1
X_18670_ _18670_/A vssd1 vssd1 vccd1 vccd1 _18826_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15882_ _15970_/A _15826_/C _15826_/A _15828_/X _15836_/X vssd1 vssd1 vccd1 vccd1
+ _15883_/B sky130_fd_sc_hd__a32oi_2
X_17621_ _17375_/Y _17376_/Y _17513_/B vssd1 vssd1 vccd1 vccd1 _17622_/B sky130_fd_sc_hd__o21ai_1
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14833_ _14828_/Y _14829_/X _14832_/X vssd1 vssd1 vccd1 vccd1 _14836_/C sky130_fd_sc_hd__a21o_1
XFILLER_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11506__A _11506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _17552_/A _17552_/B _17552_/C vssd1 vssd1 vccd1 vccd1 _17553_/A sky130_fd_sc_hd__nand3_1
XFILLER_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14764_ _14745_/A _14745_/C _14745_/B vssd1 vssd1 vccd1 vccd1 _14764_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_189_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _11976_/A _11976_/B _12013_/B vssd1 vssd1 vccd1 vccd1 _11976_/Y sky130_fd_sc_hd__nand3_2
XFILLER_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _16475_/X _16480_/X _16493_/Y _16502_/Y vssd1 vssd1 vccd1 vccd1 _16519_/A
+ sky130_fd_sc_hd__o22ai_1
X_13715_ _13856_/A vssd1 vssd1 vccd1 vccd1 _13821_/B sky130_fd_sc_hd__buf_2
XFILLER_60_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17483_ _17490_/A _17490_/B _17490_/C vssd1 vssd1 vccd1 vccd1 _17483_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14695_ _14695_/A _14695_/B _14695_/C vssd1 vssd1 vccd1 vccd1 _14696_/A sky130_fd_sc_hd__nand3_1
XFILLER_44_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19222_ _19208_/Y _19209_/Y _19210_/Y _19221_/Y vssd1 vssd1 vccd1 vccd1 _19400_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16434_ _15879_/X _16206_/X _16432_/Y _16686_/A _16433_/Y vssd1 vssd1 vccd1 vccd1
+ _16664_/B sky130_fd_sc_hd__o2111ai_4
X_13646_ _13672_/B _13672_/C _13672_/A vssd1 vssd1 vccd1 vccd1 _13674_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _16369_/A _16627_/A _16369_/C vssd1 vssd1 vccd1 vccd1 _16365_/X sky130_fd_sc_hd__and3_1
X_19153_ _15888_/A _18493_/A _18514_/Y vssd1 vssd1 vccd1 vccd1 _19156_/C sky130_fd_sc_hd__o21ai_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _13577_/A vssd1 vssd1 vccd1 vccd1 _13662_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__21311__A1 _21185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18104_ _12162_/A _16711_/C _19587_/B _12156_/X _12163_/X vssd1 vssd1 vccd1 vccd1
+ _18109_/A sky130_fd_sc_hd__a32oi_4
X_15316_ _15326_/A _15325_/A _16256_/C _12003_/C vssd1 vssd1 vccd1 vccd1 _15329_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_9_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12528_ _12528_/A _12550_/C vssd1 vssd1 vccd1 vccd1 _12771_/A sky130_fd_sc_hd__nor2_2
XFILLER_158_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19084_ _19004_/Y _19237_/A _19035_/X _19037_/X vssd1 vssd1 vccd1 vccd1 _19088_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_16296_ _11462_/A _15412_/A _16295_/Y vssd1 vssd1 vccd1 vccd1 _16296_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21862__A2 _13305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20554__A _20554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18035_ _18035_/A _18035_/B vssd1 vssd1 vccd1 vccd1 _18036_/B sky130_fd_sc_hd__xnor2_1
X_15247_ _15247_/A _15246_/X vssd1 vssd1 vccd1 vccd1 _15247_/X sky130_fd_sc_hd__or2b_1
X_12459_ _16465_/A _12734_/A _20255_/C vssd1 vssd1 vccd1 vccd1 _12459_/Y sky130_fd_sc_hd__nor3_1
XFILLER_126_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18024__A _19983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1030 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15178_ _15178_/A _15178_/B vssd1 vssd1 vccd1 vccd1 _15179_/A sky130_fd_sc_hd__and2_1
XFILLER_67_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11895__B _11895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16484__B1_N _22967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14129_ _14191_/A vssd1 vssd1 vccd1 vccd1 _14727_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17294__A2 _17286_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19986_ _19985_/A _19985_/D _18023_/X _19941_/D vssd1 vssd1 vccd1 vccd1 _19986_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12072__A _17006_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1088 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18937_ _18937_/A vssd1 vssd1 vccd1 vccd1 _18937_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18868_ _12114_/X _18330_/X _18849_/C _19013_/B vssd1 vssd1 vccd1 vccd1 _18869_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_95_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17819_ _17819_/A vssd1 vssd1 vccd1 vccd1 _17927_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18799_ _18795_/X _17388_/A _18613_/B _18797_/Y _18798_/Y vssd1 vssd1 vccd1 vccd1
+ _18799_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_48_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20830_ _20830_/A _20830_/B _20830_/C vssd1 vssd1 vccd1 vccd1 _20830_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__22820__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_719 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20761_ _20761_/A _20761_/B vssd1 vssd1 vccd1 vccd1 _20827_/D sky130_fd_sc_hd__nand2_1
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22500_ _22745_/Q input52/X _22508_/S vssd1 vssd1 vccd1 vccd1 _22501_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20692_ _20587_/B _20577_/B _20584_/Y vssd1 vssd1 vccd1 vccd1 _20695_/B sky130_fd_sc_hd__o21ai_1
XFILLER_149_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22431_ _22715_/Q input54/X _22435_/S vssd1 vssd1 vccd1 vccd1 _22432_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16309__B2 _15319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16942__A _18192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22362_ _22359_/Y _22360_/X _22368_/A vssd1 vssd1 vccd1 vccd1 _22364_/A sky130_fd_sc_hd__a21oi_1
XFILLER_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21313_ _21313_/A _21478_/A vssd1 vssd1 vccd1 vccd1 _21467_/A sky130_fd_sc_hd__nand2_2
XANTENNA__15558__A _18107_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15532__A2 _15531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22293_ _22291_/Y _22292_/Y _22251_/B _22208_/A vssd1 vssd1 vccd1 vccd1 _22294_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_190_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21244_ _13339_/Y _13353_/Y _13359_/X _13387_/X vssd1 vssd1 vccd1 vccd1 _21248_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21175_ _13343_/A _13364_/Y _13265_/A _21174_/Y _13635_/A vssd1 vssd1 vccd1 vccd1
+ _21176_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_132_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20126_ _15355_/A _15355_/B _12718_/X vssd1 vssd1 vccd1 vccd1 _20126_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20057_ _20057_/A _20057_/B vssd1 vssd1 vccd1 vccd1 _20058_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11857__A1 _19418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19982__A1 _19983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _12083_/B vssd1 vssd1 vccd1 vccd1 _11831_/C sky130_fd_sc_hd__clkbuf_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18537__A2 _12158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19212__B _19587_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11932_/A _11932_/B _11932_/C vssd1 vssd1 vccd1 vccd1 _11761_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ _20959_/A _20959_/B vssd1 vssd1 vccd1 vccd1 _20963_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13470_/Y _13474_/X _13475_/Y _13476_/Y vssd1 vssd1 vccd1 vccd1 _13550_/A
+ sky130_fd_sc_hd__o211ai_2
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14583_/B _14583_/C _14583_/D vssd1 vssd1 vccd1 vccd1 _14775_/A sky130_fd_sc_hd__nor3_2
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11842_/B _11842_/C vssd1 vssd1 vccd1 vccd1 _11692_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13431_ _22846_/Q vssd1 vssd1 vccd1 vccd1 _21848_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22629_ _22629_/A vssd1 vssd1 vccd1 vccd1 _22802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15771__A2 _15646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18770__C _18770_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11388__A3 _11404_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16150_ _16150_/A _16150_/B vssd1 vssd1 vccd1 vccd1 _16168_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13782__A1 _14199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13362_ _21964_/A _13361_/X _13274_/Y _13281_/A vssd1 vssd1 vccd1 vccd1 _21249_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20647__A3 _20454_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19585__D _19585_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15101_ _15101_/A _15101_/B _15205_/B vssd1 vssd1 vccd1 vccd1 _15103_/A sky130_fd_sc_hd__and3_1
X_12313_ _22819_/Q vssd1 vssd1 vccd1 vccd1 _12802_/C sky130_fd_sc_hd__clkbuf_2
X_16081_ _16081_/A _16081_/B vssd1 vssd1 vccd1 vccd1 _16082_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13293_ _21188_/B vssd1 vssd1 vccd1 vccd1 _13297_/A sky130_fd_sc_hd__inv_2
XANTENNA__17386__C _20675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15032_ _15031_/B _15088_/B _15031_/A vssd1 vssd1 vccd1 vccd1 _15033_/B sky130_fd_sc_hd__a21oi_1
XFILLER_181_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12244_ _18239_/B vssd1 vssd1 vccd1 vccd1 _18249_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19265__A3 _19941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18779__A _18779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19840_ _19768_/B _17401_/C _17401_/D _19945_/C _17929_/A vssd1 vssd1 vccd1 vccd1
+ _19842_/C sky130_fd_sc_hd__a32o_1
XANTENNA__18473__A1 _18770_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12175_ _12175_/A vssd1 vssd1 vccd1 vccd1 _18165_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19771_ _19771_/A vssd1 vssd1 vccd1 vccd1 _19945_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_150_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16983_ _17188_/A _16981_/A _16982_/A vssd1 vssd1 vccd1 vccd1 _16983_/X sky130_fd_sc_hd__a21o_1
XFILLER_1_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18722_ _18722_/A _18722_/B _18722_/C _18722_/D vssd1 vssd1 vccd1 vccd1 _18723_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18225__A1 _12220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15934_ _15934_/A vssd1 vssd1 vccd1 vccd1 _15935_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__22843__CLK _22937_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18653_ _18653_/A _18653_/B vssd1 vssd1 vccd1 vccd1 _18654_/C sky130_fd_sc_hd__nand2_1
XFILLER_92_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16787__A1 _16178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15865_ _16192_/D vssd1 vssd1 vccd1 vccd1 _17039_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20583__A2 _16611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17604_ _17058_/A _17603_/Y _17516_/Y vssd1 vssd1 vccd1 vccd1 _17605_/A sky130_fd_sc_hd__a21oi_4
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14816_ _14816_/A _14816_/B vssd1 vssd1 vccd1 vccd1 _14816_/Y sky130_fd_sc_hd__nand2_1
X_18584_ _18437_/Y _18440_/Y _18586_/C vssd1 vssd1 vccd1 vccd1 _18587_/A sky130_fd_sc_hd__o21bai_1
XFILLER_18_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _15775_/B _15775_/C _15795_/X vssd1 vssd1 vccd1 vccd1 _15801_/A sky130_fd_sc_hd__a21o_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17535_ _17535_/A _17535_/B vssd1 vssd1 vccd1 vccd1 _17535_/Y sky130_fd_sc_hd__nand2_1
X_11959_ _11949_/X _11952_/Y _11957_/Y _11958_/Y vssd1 vssd1 vccd1 vccd1 _12220_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14747_ _14747_/A _14747_/B _14747_/C vssd1 vssd1 vccd1 vccd1 _14749_/B sky130_fd_sc_hd__nand3_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17466_ _17466_/A _17466_/B _17467_/A vssd1 vssd1 vccd1 vccd1 _17469_/A sky130_fd_sc_hd__and3_1
XFILLER_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14678_ _14673_/Y _14674_/X _14677_/X vssd1 vssd1 vccd1 vccd1 _14745_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__16944__D1 _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14014__A2 _13924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19205_ _11859_/X _11861_/X _18629_/B vssd1 vssd1 vccd1 vccd1 _19211_/C sky130_fd_sc_hd__o21ai_2
X_16417_ _16418_/A _16418_/B _16417_/C vssd1 vssd1 vccd1 vccd1 _16695_/C sky130_fd_sc_hd__nand3_1
X_13629_ _13650_/A vssd1 vssd1 vccd1 vccd1 _21399_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17397_ _19687_/B vssd1 vssd1 vccd1 vccd1 _19768_/C sky130_fd_sc_hd__buf_2
XANTENNA__20099__A1 _20486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19136_ _19136_/A _19281_/A vssd1 vssd1 vccd1 vccd1 _19137_/C sky130_fd_sc_hd__nand2_1
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16348_ _20582_/C vssd1 vssd1 vccd1 vccd1 _21011_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__22914__D _22914_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15378__A _15378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19067_ _19043_/X _17819_/A _19046_/A _19065_/X vssd1 vssd1 vccd1 vccd1 _19067_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16279_ _15568_/B _15563_/Y _15558_/Y _15559_/Y vssd1 vssd1 vccd1 vccd1 _16595_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_69_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13525__A1 _13350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18018_ _22906_/Q vssd1 vssd1 vccd1 vccd1 _18051_/A sky130_fd_sc_hd__inv_2
XFILLER_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20271__A1 _20261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19969_ _19974_/B _19974_/C vssd1 vssd1 vccd1 vccd1 _19972_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12530__A _12771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18621__D1 _19418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21931_ _21931_/A _21931_/B vssd1 vssd1 vccd1 vccd1 _22145_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16937__A _19694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22658__B _22658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19313__A _19313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21862_ _13305_/A _13305_/B _21376_/X vssd1 vssd1 vccd1 vccd1 _21862_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20813_ _20804_/Y _20884_/B _20808_/Y vssd1 vssd1 vccd1 vccd1 _20813_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14457__A _14863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21793_ _21650_/X _21653_/Y _21661_/Y _21662_/Y vssd1 vssd1 vccd1 vccd1 _21793_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__20326__A2 _12576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20744_ _20806_/B vssd1 vssd1 vccd1 vccd1 _21017_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1110 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20675_ _20675_/A _20675_/B _20675_/C vssd1 vssd1 vccd1 vccd1 _20676_/B sky130_fd_sc_hd__nand3_2
XANTENNA__14556__A3 _14554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22414_ _22414_/A vssd1 vssd1 vccd1 vccd1 _22707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11775__B1 _11774_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19983__A _19983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22345_ _22295_/Y _22343_/Y _22344_/Y _22324_/A vssd1 vssd1 vccd1 vccd1 _22346_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_191_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22276_ _22277_/A _22277_/B vssd1 vssd1 vccd1 vccd1 _22317_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22613__S _22619_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18455__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17258__A2 _12294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21227_ _21848_/B _21227_/B _21638_/C vssd1 vssd1 vccd1 vccd1 _21227_/X sky130_fd_sc_hd__and3_1
XFILLER_160_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22866__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21158_ _21162_/A _21162_/B vssd1 vssd1 vccd1 vccd1 _22927_/D sky130_fd_sc_hd__xor2_4
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22539__A0 _13973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20109_ _12680_/X _16715_/A _20098_/D _20098_/B vssd1 vssd1 vccd1 vccd1 _20109_/Y
+ sky130_fd_sc_hd__a31oi_4
X_13980_ _14009_/C _14009_/D vssd1 vssd1 vccd1 vccd1 _14007_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12440__A _20461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21089_ _21090_/A _21090_/B _21090_/C vssd1 vssd1 vccd1 vccd1 _21091_/A sky130_fd_sc_hd__a21oi_1
XFILLER_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12931_ _12928_/X _12968_/D _12718_/X _16155_/A _12682_/X vssd1 vssd1 vccd1 vccd1
+ _12931_/X sky130_fd_sc_hd__o221a_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17966__B1 _22904_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16769__B2 _16496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_844 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17430__A2 _19336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _15616_/X _16397_/A _15649_/X _16361_/A vssd1 vssd1 vccd1 vccd1 _15650_/X
+ sky130_fd_sc_hd__o211a_1
X_12862_ _12862_/A _12862_/B vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__nand2_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13047__A3 _13041_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _11809_/A _11809_/B _12024_/A _11810_/C vssd1 vssd1 vccd1 vccd1 _11930_/B
+ sky130_fd_sc_hd__o211ai_1
X_14601_ _14712_/A _14712_/B _14600_/Y vssd1 vssd1 vccd1 vccd1 _14601_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15581_ _16016_/A _15546_/X _15472_/X _12922_/X _15580_/X vssd1 vssd1 vccd1 vccd1
+ _15581_/X sky130_fd_sc_hd__o32a_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _15299_/C _15299_/D _22825_/Q vssd1 vssd1 vccd1 vccd1 _12793_/X sky130_fd_sc_hd__and3_1
XANTENNA__15992__A2 _17539_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17320_/A _17466_/A vssd1 vssd1 vccd1 vccd1 _17323_/C sky130_fd_sc_hd__nand2_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14561_/D _14561_/B _22863_/D _14273_/C vssd1 vssd1 vccd1 vccd1 _14541_/B
+ sky130_fd_sc_hd__or4bb_2
X_11744_ _11904_/A _11905_/A _11611_/A _11611_/B vssd1 vssd1 vccd1 vccd1 _11744_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _17251_/A vssd1 vssd1 vccd1 vccd1 _17401_/D sky130_fd_sc_hd__clkbuf_4
X_14463_ _14475_/A _14475_/B _14074_/A vssd1 vssd1 vccd1 vccd1 _14463_/X sky130_fd_sc_hd__a21o_1
X_11675_ _11675_/A _11675_/B _15482_/B vssd1 vssd1 vccd1 vccd1 _11738_/A sky130_fd_sc_hd__and3_1
XFILLER_169_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16582__A _16582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16202_ _16202_/A _16202_/B vssd1 vssd1 vccd1 vccd1 _16418_/B sky130_fd_sc_hd__nand2_2
X_13414_ _13413_/B _13413_/A _13438_/B _13262_/D vssd1 vssd1 vccd1 vccd1 _21270_/A
+ sky130_fd_sc_hd__o211a_1
X_17182_ _17180_/X _17181_/Y _17173_/D _17178_/Y vssd1 vssd1 vccd1 vccd1 _17184_/B
+ sky130_fd_sc_hd__o211ai_1
X_14394_ _22803_/Q _14381_/X _14382_/X _14370_/A _22707_/Q vssd1 vssd1 vccd1 vccd1
+ _14394_/X sky130_fd_sc_hd__a32o_1
XFILLER_155_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16133_ _16133_/A _16133_/B vssd1 vssd1 vccd1 vccd1 _16134_/A sky130_fd_sc_hd__nand2_1
XFILLER_139_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13345_ _13345_/A vssd1 vssd1 vccd1 vccd1 _13345_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18694__A1 _11800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18005__C _22905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _16064_/A _16064_/B vssd1 vssd1 vccd1 vccd1 _16064_/Y sky130_fd_sc_hd__nand2_1
X_13276_ _21853_/A _21259_/B _21259_/C _13272_/Y _13275_/X vssd1 vssd1 vccd1 vccd1
+ _13276_/X sky130_fd_sc_hd__o32a_1
XFILLER_142_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15015_ _15015_/A _15015_/B _15015_/C vssd1 vssd1 vccd1 vccd1 _15017_/A sky130_fd_sc_hd__and3_1
XFILLER_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12227_ _12227_/A _12227_/B _12227_/C vssd1 vssd1 vccd1 vccd1 _12241_/C sky130_fd_sc_hd__nand3_1
XFILLER_170_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19823_ _19823_/A vssd1 vssd1 vccd1 vccd1 _19881_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18997__A2 _18889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12158_ _12158_/A vssd1 vssd1 vccd1 vccd1 _12158_/X sky130_fd_sc_hd__buf_2
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18659__D _18659_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13446__A _13465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19754_ _22920_/Q _19754_/B vssd1 vssd1 vccd1 vccd1 _19891_/D sky130_fd_sc_hd__or2_1
XANTENNA__16472__A3 _20129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16966_ _16967_/A _16967_/B _16967_/C vssd1 vssd1 vccd1 vccd1 _16966_/X sky130_fd_sc_hd__and3_1
XANTENNA__11892__C _16130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12089_ _12089_/A _12089_/B vssd1 vssd1 vccd1 vccd1 _12188_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12350__A _20323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_660 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18705_ _18705_/A _18705_/B vssd1 vssd1 vccd1 vccd1 _18709_/A sky130_fd_sc_hd__nand2_1
X_15917_ _15898_/Y _15913_/Y _15915_/Y _15916_/Y vssd1 vssd1 vccd1 vccd1 _15917_/X
+ sky130_fd_sc_hd__o211a_1
X_19685_ _19684_/A _19684_/B _19684_/C vssd1 vssd1 vccd1 vccd1 _19685_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16897_ _16644_/Y _16896_/Y _16889_/C _16672_/X vssd1 vssd1 vccd1 vccd1 _17215_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__20556__A2 _20551_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18636_ _18636_/A vssd1 vssd1 vccd1 vccd1 _18778_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _15853_/B _15843_/Y _15844_/Y _15847_/Y vssd1 vssd1 vccd1 vccd1 _15883_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__22909__D _22909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18567_ _18443_/Y _18406_/Y _18399_/Y vssd1 vssd1 vccd1 vccd1 _18569_/B sky130_fd_sc_hd__a21o_1
XFILLER_75_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15779_ _15779_/A vssd1 vssd1 vccd1 vccd1 _15780_/B sky130_fd_sc_hd__buf_2
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17518_ _17603_/D _17518_/B _17518_/C vssd1 vssd1 vccd1 vccd1 _17518_/Y sky130_fd_sc_hd__nand3b_1
XANTENNA__13994__A1 _14686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18498_ _18340_/Y _18349_/B _18337_/X _18343_/X vssd1 vssd1 vccd1 vccd1 _18499_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_178_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18691__B _18691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17449_ _17449_/A _17523_/B _17449_/C _17449_/D vssd1 vssd1 vccd1 vccd1 _17523_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21808__A2 _21677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20460_ _20460_/A vssd1 vssd1 vccd1 vccd1 _20587_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19119_ _19303_/A _19116_/A _19116_/B vssd1 vssd1 vccd1 vccd1 _19119_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20391_ _12761_/X _16179_/X _20263_/B _20264_/A _20263_/A vssd1 vssd1 vccd1 vccd1
+ _20393_/B sky130_fd_sc_hd__o221ai_4
XANTENNA__12525__A _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22889__CLK _22952_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22130_ _22135_/B _22170_/B vssd1 vssd1 vccd1 vccd1 _22134_/A sky130_fd_sc_hd__nand2_1
XANTENNA__21838__A _21838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22061_ _22051_/Y _22054_/Y _22060_/X vssd1 vssd1 vccd1 vccd1 _22064_/C sky130_fd_sc_hd__a21o_1
XFILLER_82_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21012_ _21082_/A _21048_/B _21048_/C _12671_/X _17922_/A vssd1 vssd1 vccd1 vccd1
+ _21012_/X sky130_fd_sc_hd__o32a_1
XANTENNA__21441__B1 _21423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16999__A1 _16098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20795__A2 _17313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22963_ _22964_/CLK _22963_/D vssd1 vssd1 vccd1 vccd1 _22963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21744__A1 _21383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19043__A _19043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17412__A2 _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21914_ _22008_/A _22007_/A _22007_/B _21912_/Y _21913_/Y vssd1 vssd1 vccd1 vccd1
+ _22024_/A sky130_fd_sc_hd__a311oi_1
XFILLER_167_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21292__B _22673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22894_ _22951_/CLK _22894_/D vssd1 vssd1 vccd1 vccd1 _22894_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_bq_clk_i clkbuf_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_167_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21845_ _21897_/A _21897_/B vssd1 vssd1 vccd1 vccd1 _21933_/A sky130_fd_sc_hd__xor2_1
XANTENNA__15721__D _19154_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15974__A2 _15427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21776_ _21775_/Y _21730_/C _21730_/D _21737_/A vssd1 vssd1 vccd1 vccd1 _21841_/C
+ sky130_fd_sc_hd__a31oi_4
XFILLER_168_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20917__A _20917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17612__B1_N _22899_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_21 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15187__B1 _15182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20727_ _20620_/C _20621_/B _20726_/X vssd1 vssd1 vccd1 vccd1 _20818_/A sky130_fd_sc_hd__a21oi_4
XFILLER_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17929__C _21011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11460_ _11504_/A _11505_/A _11506_/A vssd1 vssd1 vccd1 vccd1 _12090_/C sky130_fd_sc_hd__o21ai_4
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20658_ _20658_/A _20658_/B _20658_/C vssd1 vssd1 vccd1 vccd1 _20658_/Y sky130_fd_sc_hd__nand3_1
XFILLER_99_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11391_ _18482_/B vssd1 vssd1 vccd1 vccd1 _18984_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_109_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12435__A _22818_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20589_ _13022_/C _20697_/C _20577_/Y _20578_/X vssd1 vssd1 vccd1 vccd1 _20704_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1096 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13130_ _13449_/A vssd1 vssd1 vccd1 vccd1 _21367_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22328_ _22328_/A vssd1 vssd1 vccd1 vccd1 _22942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13061_ _13138_/C vssd1 vssd1 vccd1 vccd1 _21448_/C sky130_fd_sc_hd__clkbuf_2
X_22259_ _22243_/B _22243_/A _22215_/A _22215_/B vssd1 vssd1 vccd1 vccd1 _22259_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18122__A _18483_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12012_ _11976_/A _11797_/B _11789_/X _11791_/X vssd1 vssd1 vccd1 vccd1 _12013_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__12712__A2 _17401_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A wb_dat_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16820_ _16815_/Y _16816_/Y _16819_/X vssd1 vssd1 vccd1 vccd1 _16822_/B sky130_fd_sc_hd__o21ai_4
XFILLER_66_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16751_ _16751_/A vssd1 vssd1 vccd1 vccd1 _16753_/A sky130_fd_sc_hd__inv_2
X_13963_ _13963_/A _13963_/B _13963_/C _13963_/D vssd1 vssd1 vccd1 vccd1 _14583_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_98_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14870__C1 _22766_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15702_ _15978_/C _17525_/C _15411_/A _15419_/Y vssd1 vssd1 vccd1 vccd1 _15704_/A
+ sky130_fd_sc_hd__a22o_1
X_19470_ _19792_/A _19470_/B _19618_/A _19470_/D vssd1 vssd1 vccd1 vccd1 _19476_/B
+ sky130_fd_sc_hd__and4_1
X_12914_ _12958_/B _12958_/C _12958_/A vssd1 vssd1 vccd1 vccd1 _13004_/B sky130_fd_sc_hd__a21oi_2
XFILLER_185_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16682_ _17502_/A _16680_/X _16681_/Y vssd1 vssd1 vccd1 vccd1 _16682_/Y sky130_fd_sc_hd__o21ai_1
X_13894_ _22761_/Q vssd1 vssd1 vccd1 vccd1 _13963_/C sky130_fd_sc_hd__inv_2
XFILLER_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15912__C _15912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18421_ _18275_/B _18275_/A _18232_/X vssd1 vssd1 vccd1 vccd1 _18423_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15633_ _15633_/A _15633_/B _16450_/C vssd1 vssd1 vccd1 vccd1 _15638_/A sky130_fd_sc_hd__nand3_1
X_12845_ _12792_/A _12487_/C _12721_/A _16178_/A vssd1 vssd1 vccd1 vccd1 _12848_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21499__B1 _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _18355_/B vssd1 vssd1 vccd1 vccd1 _18520_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _15559_/Y _15558_/Y _15568_/B _15563_/Y vssd1 vssd1 vccd1 vccd1 _15565_/D
+ sky130_fd_sc_hd__o211ai_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12776_/A vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_543 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17303_ _17307_/B _17307_/C vssd1 vssd1 vccd1 vccd1 _17304_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18903__A2 _18893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11727_ _12046_/A _15481_/A _11727_/C vssd1 vssd1 vccd1 vccd1 _11941_/A sky130_fd_sc_hd__nand3_1
X_14515_ _14515_/A _14515_/B _14515_/C vssd1 vssd1 vccd1 vccd1 _14516_/C sky130_fd_sc_hd__nand3_2
X_18283_ _18200_/Y _18451_/A _18281_/Y _18282_/X vssd1 vssd1 vccd1 vccd1 _18296_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_15495_ _16226_/A vssd1 vssd1 vccd1 vccd1 _15495_/X sky130_fd_sc_hd__buf_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15717__A2 _16720_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13151__D _21494_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17839__C _17839_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17234_ _17234_/A vssd1 vssd1 vccd1 vccd1 _18200_/A sky130_fd_sc_hd__clkbuf_4
X_14446_ _22965_/Q vssd1 vssd1 vccd1 vccd1 _16226_/B sky130_fd_sc_hd__buf_2
X_11658_ _11712_/C vssd1 vssd1 vccd1 vccd1 _15482_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17165_ _19694_/A _17385_/B _17128_/Y _17288_/A vssd1 vssd1 vccd1 vccd1 _17169_/A
+ sky130_fd_sc_hd__a22o_1
X_14377_ _15369_/B vssd1 vssd1 vccd1 vccd1 _16324_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_183_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18667__B2 _18666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11589_ _11589_/A vssd1 vssd1 vccd1 vccd1 _11589_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16116_ _16115_/X _16070_/Y _16064_/Y vssd1 vssd1 vccd1 vccd1 _16169_/B sky130_fd_sc_hd__o21ai_1
X_13328_ _21367_/A _21367_/B _13502_/D _21448_/A _13332_/C vssd1 vssd1 vccd1 vccd1
+ _13337_/A sky130_fd_sc_hd__a32o_1
XFILLER_155_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17096_ _16919_/A _16919_/B _16919_/C _17095_/X vssd1 vssd1 vccd1 vccd1 _17341_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_127_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16047_ _16047_/A _16047_/B _16047_/C _16047_/D vssd1 vssd1 vccd1 vccd1 _16126_/A
+ sky130_fd_sc_hd__nand4_4
X_13259_ _13259_/A vssd1 vssd1 vccd1 vccd1 _13650_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17574__C _17574_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18967__A _22914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19806_ _19872_/A _19806_/B vssd1 vssd1 vccd1 vccd1 _19807_/B sky130_fd_sc_hd__nand2_1
XANTENNA__15102__B1 _15101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17998_ _17957_/A _17962_/Y _17999_/A vssd1 vssd1 vccd1 vccd1 _18048_/A sky130_fd_sc_hd__o21ai_2
XFILLER_38_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18686__B _19687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19737_ _19689_/A _19836_/C _19419_/B _18028_/A _19607_/A vssd1 vssd1 vccd1 vccd1
+ _19742_/A sky130_fd_sc_hd__a41o_1
XFILLER_111_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11408__B _22955_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16949_ _15450_/X _16758_/A _16946_/X _16948_/X vssd1 vssd1 vccd1 vccd1 _16949_/Y
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__21726__A1 _13423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18198__A3 _19353_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13904__A _22869_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19668_ _19680_/A _19880_/A _19670_/B _19670_/A vssd1 vssd1 vccd1 vccd1 _19674_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18619_ _18452_/X _18450_/A _18616_/Y _18618_/Y vssd1 vssd1 vccd1 vccd1 _18619_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13623__B _21498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19599_ _19591_/Y _19594_/Y _19598_/Y vssd1 vssd1 vccd1 vccd1 _19608_/A sky130_fd_sc_hd__o21ai_1
XFILLER_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11424__A _12154_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21630_ _21633_/A _21633_/B _21629_/Y _21449_/B vssd1 vssd1 vccd1 vccd1 _21638_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_178_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20737__A _20737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21561_ _21561_/A _21561_/B vssd1 vssd1 vccd1 vccd1 _21561_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17563__D1 _16124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17111__A _17111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20512_ _20519_/A _20519_/B vssd1 vssd1 vccd1 vccd1 _20512_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21492_ _21488_/Y _21490_/Y _21504_/A vssd1 vssd1 vccd1 vccd1 _21492_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_21_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12927__C1 _20793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20443_ _20549_/C _20549_/D vssd1 vssd1 vccd1 vccd1 _20444_/B sky130_fd_sc_hd__nand2_1
XANTENNA__19855__B1 _19793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20465__A1 _13022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20374_ _20511_/B _20354_/X _20360_/X _20366_/B _20366_/C vssd1 vssd1 vccd1 vccd1
+ _20375_/C sky130_fd_sc_hd__o2111ai_1
X_22113_ _22113_/A _22113_/B _22113_/C vssd1 vssd1 vccd1 vccd1 _22171_/B sky130_fd_sc_hd__nand3_2
XFILLER_192_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15892__A1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15892__B2 _11505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22044_ _22044_/A vssd1 vssd1 vccd1 vccd1 _22044_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19622__A3 _19772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12421__C _16319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16841__B1 _16842_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22904__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16397__A _16397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13814__A _13814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22946_ _22948_/CLK _22946_/D vssd1 vssd1 vccd1 vccd1 _22946_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18594__B1 _22912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14629__B _14629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_622 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22877_ _22944_/CLK input69/X vssd1 vssd1 vccd1 vccd1 _22877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12630_ _12630_/A _12630_/B _12630_/C vssd1 vssd1 vccd1 vccd1 _12640_/B sky130_fd_sc_hd__nand3_1
XFILLER_169_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21828_ _21433_/A _22674_/Q _21571_/Y _21570_/A vssd1 vssd1 vccd1 vccd1 _21828_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_58_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ _12561_/A vssd1 vssd1 vccd1 vccd1 _12769_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21759_ _21761_/A _21761_/B _21760_/A _21760_/B vssd1 vssd1 vccd1 vccd1 _21765_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__14645__A _22863_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ _11512_/A vssd1 vssd1 vccd1 vccd1 _18203_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_12_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14300_ _14300_/A _14300_/B _14300_/C _14300_/D vssd1 vssd1 vccd1 vccd1 _14305_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_156_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15280_ _15287_/D _22881_/Q _15288_/C vssd1 vssd1 vccd1 vccd1 _15282_/A sky130_fd_sc_hd__and3_1
XFILLER_12_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12492_ _20359_/B vssd1 vssd1 vccd1 vccd1 _20255_/B sky130_fd_sc_hd__buf_2
XFILLER_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14231_ _14231_/A _14231_/B _14231_/C _15050_/B vssd1 vssd1 vccd1 vccd1 _14233_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_184_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18649__A1 _12157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11443_ _15415_/C vssd1 vssd1 vccd1 vccd1 _15912_/C sky130_fd_sc_hd__buf_2
XFILLER_109_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18649__B2 _17422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12165__A _12165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19310__A2 _19480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14162_ _14147_/A _14147_/B _14159_/Y _14161_/X vssd1 vssd1 vccd1 vccd1 _14163_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_165_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11374_ _11374_/A vssd1 vssd1 vccd1 vccd1 _11395_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_180_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ _13112_/Y _13243_/A _13057_/C vssd1 vssd1 vccd1 vccd1 _13345_/A sky130_fd_sc_hd__a21o_1
X_18970_ _18970_/A _18970_/B _18970_/C vssd1 vssd1 vccd1 vccd1 _18970_/Y sky130_fd_sc_hd__nand3_1
XFILLER_124_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14093_ _14094_/B _14094_/C _14094_/A vssd1 vssd1 vccd1 vccd1 _14093_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_140_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14380__A _14380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15907__C _18985_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _17907_/A _17907_/B _17920_/Y vssd1 vssd1 vccd1 vccd1 _17953_/A sky130_fd_sc_hd__a21oi_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13044_/A _13044_/B _13044_/C vssd1 vssd1 vccd1 vccd1 _20304_/A sky130_fd_sc_hd__nand3_4
XFILLER_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1112 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11509__A _12090_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17852_ _17705_/Y _17623_/Y _17607_/X _17708_/Y vssd1 vssd1 vccd1 vccd1 _17853_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__18821__A1 _19651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16803_ _16803_/A _16803_/B vssd1 vssd1 vccd1 vccd1 _16971_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12449__A1 _16465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17783_ _17775_/X _17779_/X _17787_/A vssd1 vssd1 vccd1 vccd1 _17799_/A sky130_fd_sc_hd__a21o_1
XANTENNA__15923__B _16011_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14995_ _14934_/A _15154_/D _14996_/D _14996_/B _14996_/C vssd1 vssd1 vccd1 vccd1
+ _15001_/B sky130_fd_sc_hd__a32o_1
XFILLER_82_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19522_ _19532_/A _19525_/A _19514_/X vssd1 vssd1 vccd1 vccd1 _19523_/D sky130_fd_sc_hd__a21o_1
X_16734_ _16734_/A _16734_/B _16734_/C vssd1 vssd1 vccd1 vccd1 _16734_/X sky130_fd_sc_hd__and3_2
XFILLER_35_803 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13946_ _13926_/Y _13927_/X _13931_/X _14157_/A _15058_/C vssd1 vssd1 vccd1 vccd1
+ _13947_/C sky130_fd_sc_hd__o2111ai_1
XANTENNA__16100__A _16100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19453_ _19410_/A _19410_/B _19410_/C _19435_/X vssd1 vssd1 vccd1 vccd1 _19555_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16665_ _16665_/A vssd1 vssd1 vccd1 vccd1 _16665_/X sky130_fd_sc_hd__clkbuf_2
X_13877_ _13877_/A _13877_/B vssd1 vssd1 vccd1 vccd1 _13877_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__20931__A2 _17816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18404_ _18404_/A vssd1 vssd1 vccd1 vccd1 _18404_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18953__C _18953_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15616_ _15616_/A vssd1 vssd1 vccd1 vccd1 _15616_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19384_ _19340_/A _19340_/B _19332_/Y _19337_/Y vssd1 vssd1 vccd1 vccd1 _19530_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__13162__C _13162_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ _22698_/Q vssd1 vssd1 vccd1 vccd1 _15362_/D sky130_fd_sc_hd__clkinv_2
X_16596_ _16596_/A _16596_/B vssd1 vssd1 vccd1 vccd1 _16602_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18335_ _11511_/X _18330_/X _11774_/Y _18980_/C _18529_/A vssd1 vssd1 vccd1 vccd1
+ _18354_/B sky130_fd_sc_hd__o221ai_4
X_15547_ _15545_/X _15546_/X _15439_/X _15524_/X _16265_/A vssd1 vssd1 vccd1 vccd1
+ _15547_/X sky130_fd_sc_hd__o221a_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18888__A1 _18127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ _12988_/A vssd1 vssd1 vccd1 vccd1 _13022_/A sky130_fd_sc_hd__buf_2
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16473__C _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18266_ _18266_/A _18266_/B vssd1 vssd1 vccd1 vccd1 _22890_/D sky130_fd_sc_hd__xor2_1
XFILLER_30_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15478_ _19316_/A _16059_/A _15309_/B _15472_/X _15574_/C vssd1 vssd1 vccd1 vccd1
+ _15479_/C sky130_fd_sc_hd__o221ai_1
XANTENNA__16363__A2 _16431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17217_ _17060_/A _17060_/B _16665_/A vssd1 vssd1 vccd1 vccd1 _17371_/B sky130_fd_sc_hd__a21o_1
XANTENNA__16192__D _16192_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14374__A1 _14369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14429_ _14429_/A vssd1 vssd1 vccd1 vccd1 _14430_/A sky130_fd_sc_hd__buf_4
XANTENNA__16770__A _16770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18197_ _18197_/A _19351_/C _18197_/C _18288_/A vssd1 vssd1 vccd1 vccd1 _18197_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_162_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18104__A3 _19587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17148_ _20129_/A _17405_/A _17406_/A vssd1 vssd1 vccd1 vccd1 _17149_/B sky130_fd_sc_hd__and3_1
XFILLER_190_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17079_ _17054_/Y _17078_/Y _17058_/B vssd1 vssd1 vccd1 vccd1 _17079_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_143_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11428__A_N _11430_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20090_ _20219_/A _20219_/B vssd1 vssd1 vccd1 vccd1 _20090_/Y sky130_fd_sc_hd__nand2_2
XFILLER_124_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12522__B _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18812__A1 _11502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22800_ _22800_/CLK _22800_/D vssd1 vssd1 vccd1 vccd1 _22800_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20992_ _20992_/A _20992_/B _20992_/C vssd1 vssd1 vccd1 vccd1 _21062_/A sky130_fd_sc_hd__nand3_2
XFILLER_77_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22372__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22731_ _22731_/CLK _22731_/D vssd1 vssd1 vccd1 vccd1 _22731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_655 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22662_ _22662_/A _22662_/B vssd1 vssd1 vccd1 vccd1 _22663_/A sky130_fd_sc_hd__and2_1
XFILLER_129_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21613_ _21613_/A vssd1 vssd1 vccd1 vccd1 _21742_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18879__A1 _15904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12612__A1 _12450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_874 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22593_ _11306_/X input57/X _22597_/S vssd1 vssd1 vccd1 vccd1 _22594_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12612__B2 _15450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20186__B _20442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21544_ _21537_/Y _21538_/Y _21531_/C _21531_/B vssd1 vssd1 vccd1 vccd1 _21545_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_138_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15562__B1 _16779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21475_ _21876_/A _21749_/A _21588_/B vssd1 vssd1 vccd1 vccd1 _21482_/B sky130_fd_sc_hd__nand3_2
XFILLER_181_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19694__C _19771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20914__B _21019_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20426_ _20395_/A _20395_/B _20388_/Y _20405_/Y vssd1 vssd1 vccd1 vccd1 _20426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22832__D _22844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15296__A _22887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16511__C1 _15810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20357_ _20357_/A _20357_/B _20357_/C vssd1 vssd1 vccd1 vccd1 _20358_/B sky130_fd_sc_hd__nand3_1
XFILLER_162_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12713__A _20255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20288_ _20280_/Y _20281_/X _20269_/X _20274_/Y vssd1 vssd1 vccd1 vccd1 _20290_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22027_ _22003_/X _21999_/Y _22002_/Y _21997_/Y vssd1 vssd1 vccd1 vccd1 _22080_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_49_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_195_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13800_ _13820_/A _13773_/A _13799_/X vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__a21o_1
XFILLER_57_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11992_ _18140_/C vssd1 vssd1 vccd1 vccd1 _12135_/A sky130_fd_sc_hd__clkbuf_2
X_14780_ _14953_/A _15107_/A _15107_/B _14781_/A _14895_/A vssd1 vssd1 vccd1 vccd1
+ _14805_/A sky130_fd_sc_hd__a32o_1
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13731_ _13810_/A _13738_/A _13963_/D _13810_/B vssd1 vssd1 vccd1 vccd1 _13798_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22929_ _22929_/CLK _22929_/D vssd1 vssd1 vccd1 vccd1 _22929_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16450_ _19318_/A _16450_/B _16450_/C vssd1 vssd1 vccd1 vccd1 _16451_/B sky130_fd_sc_hd__and3_2
XANTENNA__21480__B _21480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13662_ _13662_/A _13662_/B _13662_/C vssd1 vssd1 vccd1 vccd1 _13663_/B sky130_fd_sc_hd__and3_1
XANTENNA__16593__A2 _16598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _20502_/A _20502_/B _16712_/C vssd1 vssd1 vccd1 vccd1 _15731_/B sky130_fd_sc_hd__and3_1
X_12613_ _12605_/Y _12608_/X _12611_/Y _12612_/Y vssd1 vssd1 vccd1 vccd1 _12613_/Y
+ sky130_fd_sc_hd__o211ai_4
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16381_ _16704_/A _16704_/B _16366_/Y _16374_/Y vssd1 vssd1 vccd1 vccd1 _16391_/B
+ sky130_fd_sc_hd__o211ai_2
X_13593_ _13373_/A _13373_/B _13126_/X vssd1 vssd1 vccd1 vccd1 _13593_/X sky130_fd_sc_hd__a21o_1
XANTENNA__20126__B1 _12718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13800__B1 _13799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _18500_/C vssd1 vssd1 vccd1 vccd1 _18677_/B sky130_fd_sc_hd__buf_2
X_15332_ _15426_/B _15344_/A _15329_/X _15331_/Y vssd1 vssd1 vccd1 vccd1 _15339_/B
+ sky130_fd_sc_hd__o2bb2ai_2
X_12544_ _12561_/A vssd1 vssd1 vccd1 vccd1 _12544_/Y sky130_fd_sc_hd__inv_2
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17542__A1 _20870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18051_ _18051_/A _18069_/C _18051_/C vssd1 vssd1 vccd1 vccd1 _18051_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__14356__A1 _18127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15263_ _15263_/A _15263_/B vssd1 vssd1 vccd1 vccd1 _22686_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__14356__B2 _13973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12475_ _22691_/Q vssd1 vssd1 vccd1 vccd1 _12493_/A sky130_fd_sc_hd__buf_4
XFILLER_126_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17002_ _16714_/X _17087_/A _16719_/A vssd1 vssd1 vccd1 vccd1 _17005_/A sky130_fd_sc_hd__o21ai_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11426_ _18292_/A _11636_/A _11425_/Y vssd1 vssd1 vccd1 vccd1 _11565_/A sky130_fd_sc_hd__o21ai_4
X_14214_ _14259_/A _14259_/B _14261_/C vssd1 vssd1 vccd1 vccd1 _14214_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_137_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15194_ _15186_/X _15187_/X _15194_/C _15216_/A vssd1 vssd1 vccd1 vccd1 _15223_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14145_ _14085_/A _14085_/B _14126_/Y _14071_/Y vssd1 vssd1 vccd1 vccd1 _14146_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16648__A3 _16879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11357_ _11404_/C vssd1 vssd1 vccd1 vccd1 _11605_/A sky130_fd_sc_hd__inv_2
XFILLER_99_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13719__A _13725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12119__B1 _11634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18953_ _18953_/A _19418_/C _18953_/C vssd1 vssd1 vccd1 vccd1 _18953_/X sky130_fd_sc_hd__and3_1
X_14076_ _14085_/A _13808_/A _14721_/B _14270_/A _13829_/Y vssd1 vssd1 vccd1 vccd1
+ _14076_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_152_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11288_ _22953_/Q vssd1 vssd1 vccd1 vccd1 _11404_/C sky130_fd_sc_hd__buf_2
XANTENNA__11884__D _11895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17904_ _17904_/A _17843_/A vssd1 vssd1 vccd1 vccd1 _17949_/A sky130_fd_sc_hd__or2b_1
X_13027_ _13022_/B _20284_/A _12711_/X _13026_/X vssd1 vssd1 vccd1 vccd1 _13028_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15934__A _15934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18884_ _15932_/A _19313_/A _18880_/A vssd1 vssd1 vccd1 vccd1 _18887_/A sky130_fd_sc_hd__o21ai_1
XFILLER_117_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17835_ _17835_/A _17871_/C vssd1 vssd1 vccd1 vccd1 _17900_/A sky130_fd_sc_hd__xnor2_1
XFILLER_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17766_ _17669_/X _17679_/B _17679_/C vssd1 vssd1 vccd1 vccd1 _17768_/A sky130_fd_sc_hd__a21boi_2
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14978_ _14916_/A _14916_/B _14916_/C _14916_/D vssd1 vssd1 vccd1 vccd1 _14978_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19755__C1 _22920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19505_ _18330_/X _17400_/A _17393_/X _11598_/X vssd1 vssd1 vccd1 vccd1 _19651_/B
+ sky130_fd_sc_hd__o22ai_4
X_16717_ _18716_/A _20781_/A _20781_/B vssd1 vssd1 vccd1 vccd1 _17087_/A sky130_fd_sc_hd__nand3_2
XANTENNA__21671__A _21677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13929_ _14069_/C vssd1 vssd1 vccd1 vccd1 _14765_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17697_ _17697_/A _17697_/B _17697_/C vssd1 vssd1 vccd1 vccd1 _17699_/B sky130_fd_sc_hd__nand3_1
XFILLER_62_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19436_ _19411_/X _19555_/A _19435_/X vssd1 vssd1 vccd1 vccd1 _19436_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16648_ _16613_/D _21086_/D _16879_/B _16351_/X vssd1 vssd1 vccd1 vccd1 _16650_/C
+ sky130_fd_sc_hd__a31oi_4
XFILLER_23_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22917__D _22917_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19367_ _19357_/B _19359_/A _19352_/A _19215_/X vssd1 vssd1 vccd1 vccd1 _19368_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_176_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16579_ _16579_/A vssd1 vssd1 vccd1 vccd1 _16579_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11702__A _11702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18318_ _18691_/B vssd1 vssd1 vccd1 vccd1 _19322_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__11802__C1 _15624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19298_ _19298_/A _19298_/B vssd1 vssd1 vccd1 vccd1 _19299_/A sky130_fd_sc_hd__nand2_1
XFILLER_148_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14347__A1 _11771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18249_ _18249_/A _18249_/B vssd1 vssd1 vccd1 vccd1 _18250_/B sky130_fd_sc_hd__nor2_1
XANTENNA__14347__B2 _13896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21260_ _21260_/A _21260_/B vssd1 vssd1 vccd1 vccd1 _21266_/A sky130_fd_sc_hd__xnor2_1
XFILLER_128_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20211_ _20206_/Y _20210_/Y _20208_/X vssd1 vssd1 vccd1 vccd1 _20211_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_132_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21191_ _21185_/X _21187_/X _21609_/A vssd1 vssd1 vccd1 vccd1 _21192_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__12533__A _12540_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20142_ _20142_/A _20142_/B _20142_/C vssd1 vssd1 vccd1 vccd1 _20143_/B sky130_fd_sc_hd__nand3_2
XANTENNA__13348__B _21494_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13858__B1 _13725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19589__A2 _19464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19316__A _19316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20073_ _12540_/X _12783_/X _12796_/Y vssd1 vssd1 vccd1 vccd1 _20073_/Y sky130_fd_sc_hd__o21ai_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22593__A1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20975_ _20975_/A _20975_/B _21083_/C _20975_/D vssd1 vssd1 vccd1 vccd1 _20977_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_53_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19689__C _19689_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22714_ _22746_/CLK _22714_/D vssd1 vssd1 vccd1 vccd1 _22714_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11315__C _11404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22645_ _22645_/A vssd1 vssd1 vccd1 vccd1 _22809_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16825__D _17407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18890__A _18890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1043 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11612__A _18648_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12597__B1 _12697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22576_ _22779_/Q input54/X _22580_/S vssd1 vssd1 vccd1 vccd1 _22577_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21527_ _21514_/X _21515_/Y _21507_/Y _21512_/Y vssd1 vssd1 vccd1 vccd1 _21529_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12260_ _12260_/A vssd1 vssd1 vccd1 vccd1 _22889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21608__B1 _21494_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21458_ _21666_/A vssd1 vssd1 vccd1 vccd1 _21805_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18114__B _18278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21084__A1 _21017_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20409_ _20400_/Y _20272_/Y _20401_/Y vssd1 vssd1 vccd1 vccd1 _20409_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12191_ _11814_/B _11964_/X _12024_/A vssd1 vssd1 vccd1 vccd1 _12191_/X sky130_fd_sc_hd__o21a_1
XFILLER_147_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21389_ _21378_/A _21378_/B _21386_/X _21387_/Y _21393_/B vssd1 vssd1 vccd1 vccd1
+ _21535_/C sky130_fd_sc_hd__o221ai_4
XFILLER_134_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12162__B _15774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput87 _14376_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[14] sky130_fd_sc_hd__buf_2
X_15950_ _15759_/Y _15873_/X _15875_/Y _15876_/X vssd1 vssd1 vccd1 vccd1 _16210_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_62_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput98 _14409_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22584__A1 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input30_A wb_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14901_ _14901_/A _14930_/A _14901_/C vssd1 vssd1 vccd1 vccd1 _14930_/B sky130_fd_sc_hd__nand3_1
X_15881_ _15881_/A vssd1 vssd1 vccd1 vccd1 _15881_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17620_ _17353_/X _17230_/Y _17375_/A _17495_/X vssd1 vssd1 vccd1 vccd1 _17622_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_76_566 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14832_ _14834_/C _14834_/A _14675_/Y _15186_/D _14673_/Y vssd1 vssd1 vccd1 vccd1
+ _14832_/X sky130_fd_sc_hd__a41o_1
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22587__A _22643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _17550_/Y _17410_/X _17399_/Y vssd1 vssd1 vccd1 vccd1 _17552_/C sky130_fd_sc_hd__a21boi_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14763_ _14747_/A _14747_/B _14747_/C _14751_/B vssd1 vssd1 vccd1 vccd1 _14836_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _11793_/B _11974_/Y _11984_/B _12137_/A vssd1 vssd1 vccd1 vccd1 _12013_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16585__A _16585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _15542_/X _16494_/X _16512_/A _16501_/Y vssd1 vssd1 vccd1 vccd1 _16502_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_17_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13714_ _22767_/Q vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__inv_2
XFILLER_72_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17482_ _17341_/B _17324_/B _17324_/C vssd1 vssd1 vccd1 vccd1 _17490_/C sky130_fd_sc_hd__a21boi_1
XFILLER_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14694_ _14568_/Y _14131_/X _14688_/A _14693_/X vssd1 vssd1 vccd1 vccd1 _14695_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19221_ _19206_/Y _19211_/X _19223_/A vssd1 vssd1 vccd1 vccd1 _19221_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16433_ _16433_/A _16433_/B _16433_/C vssd1 vssd1 vccd1 vccd1 _16433_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__19896__A _19896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13645_ _13647_/A _13647_/C _13647_/B vssd1 vssd1 vccd1 vccd1 _13672_/A sky130_fd_sc_hd__o21bai_1
XFILLER_60_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19152_ _19329_/A _19694_/D _19329_/C _19329_/D vssd1 vssd1 vccd1 vccd1 _19156_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_13_872 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _16369_/A _16627_/A _16369_/C vssd1 vssd1 vccd1 vccd1 _16364_/Y sky130_fd_sc_hd__a21oi_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13576_ _13162_/A _13126_/X _13162_/C _13319_/X _13434_/X vssd1 vssd1 vccd1 vccd1
+ _13576_/X sky130_fd_sc_hd__o32a_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _18896_/C vssd1 vssd1 vccd1 vccd1 _19587_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_157_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15315_ _15714_/A _16932_/C _16257_/D _15911_/A _18680_/D vssd1 vssd1 vccd1 vccd1
+ _15315_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19083_ _18908_/A _18908_/B _19034_/Y vssd1 vssd1 vccd1 vccd1 _19088_/A sky130_fd_sc_hd__a21oi_1
X_12527_ _12516_/X _12704_/A _20134_/C _16488_/A _12526_/X vssd1 vssd1 vccd1 vccd1
+ _12543_/B sky130_fd_sc_hd__o2111ai_4
X_16295_ _16293_/X _16294_/X _12094_/D _16302_/A vssd1 vssd1 vccd1 vccd1 _16295_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__18305__A _18305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18034_ _17988_/A _17988_/B _18062_/C vssd1 vssd1 vccd1 vccd1 _18035_/B sky130_fd_sc_hd__a21boi_1
XFILLER_157_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15246_ _15259_/A _15246_/B vssd1 vssd1 vccd1 vccd1 _15246_/X sky130_fd_sc_hd__or2_1
XFILLER_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12458_ _12458_/A vssd1 vssd1 vccd1 vccd1 _17144_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_126_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11409_ _11712_/B vssd1 vssd1 vccd1 vccd1 _11659_/B sky130_fd_sc_hd__buf_2
XFILLER_158_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15177_ _14845_/B _15180_/A _15180_/B vssd1 vssd1 vccd1 vccd1 _15178_/B sky130_fd_sc_hd__o21ai_1
X_12389_ _12458_/A vssd1 vssd1 vccd1 vccd1 _17141_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_193_1042 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14128_ _14237_/A _14128_/B _14128_/C vssd1 vssd1 vccd1 vccd1 _14238_/A sky130_fd_sc_hd__nand3b_2
X_19985_ _19985_/A _20012_/A _19985_/C _19985_/D vssd1 vssd1 vccd1 vccd1 _19985_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18936_ _18927_/Y _18932_/Y _18935_/Y vssd1 vssd1 vccd1 vccd1 _18941_/A sky130_fd_sc_hd__a21o_1
XFILLER_113_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14059_ _22870_/Q vssd1 vssd1 vccd1 vccd1 _14491_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_100_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15383__B _15665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18867_ _18850_/A _18849_/C _18866_/Y vssd1 vssd1 vccd1 vccd1 _18869_/B sky130_fd_sc_hd__a21bo_1
X_17818_ _18814_/A vssd1 vssd1 vccd1 vccd1 _17819_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18798_ _18156_/X _16940_/X _18611_/Y vssd1 vssd1 vccd1 vccd1 _18798_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_36_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17749_ _17733_/A _17873_/A _17880_/A _17876_/A vssd1 vssd1 vccd1 vccd1 _17752_/C
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__12815__B2 _15637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20760_ _20890_/A _20891_/A vssd1 vssd1 vccd1 vccd1 _20761_/B sky130_fd_sc_hd__nand2_1
XFILLER_165_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19419_ _19651_/A _19419_/B _19454_/C _19455_/C vssd1 vssd1 vccd1 vccd1 _19419_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17103__B _17338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20691_ _20110_/B _20689_/Y _20690_/X vssd1 vssd1 vccd1 vccd1 _20796_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12528__A _12528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22430_ _22430_/A vssd1 vssd1 vccd1 vccd1 _22714_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11432__A _18663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17506__A1 _17502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22361_ _22352_/B _22359_/Y _22816_/Q vssd1 vssd1 vccd1 vccd1 _22368_/A sky130_fd_sc_hd__a21oi_2
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21312_ _21312_/A _21312_/B _21312_/C vssd1 vssd1 vccd1 vccd1 _21478_/A sky130_fd_sc_hd__nand3_1
XFILLER_190_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15558__B _18107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22292_ _22094_/A _22209_/Y _22290_/C vssd1 vssd1 vccd1 vccd1 _22292_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_163_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13359__A _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21243_ _21243_/A _21243_/B _21243_/C vssd1 vssd1 vccd1 vccd1 _21266_/B sky130_fd_sc_hd__nand3_2
XFILLER_190_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17809__A2 _21017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14181__C _14181_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21174_ _13162_/A _13229_/A _13162_/C _21173_/Y vssd1 vssd1 vccd1 vccd1 _21174_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15574__A _17436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20125_ _20125_/A vssd1 vssd1 vccd1 vccd1 _20155_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15150__D1 _15006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20056_ _20052_/X _20049_/A _20055_/Y _20049_/B vssd1 vssd1 vccd1 vccd1 _20063_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11857__A2 _16564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16245__A1 _15804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19982__A2 _18778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater170 _22728_/CLK vssd1 vssd1 vccd1 vccd1 _22731_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20329__B1 _20210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13822__A _22866_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14271__A3 _14575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11762_/B vssd1 vssd1 vccd1 vccd1 _11932_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ _20958_/A _20958_/B _22938_/Q vssd1 vssd1 vccd1 vccd1 _20959_/B sky130_fd_sc_hd__nand3_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17745__A1 _17386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19212__C _19687_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _12083_/B _11687_/B _11689_/Y _11690_/Y _11643_/Y vssd1 vssd1 vccd1 vccd1
+ _11842_/C sky130_fd_sc_hd__o221ai_4
XFILLER_187_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20889_ _20894_/C _20894_/B vssd1 vssd1 vccd1 vccd1 _20892_/A sky130_fd_sc_hd__nand2_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13430_ _13430_/A vssd1 vssd1 vccd1 vccd1 _21177_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22628_ _22802_/Q input44/X _22630_/S vssd1 vssd1 vccd1 vccd1 _22629_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13361_ _13361_/A vssd1 vssd1 vccd1 vccd1 _13361_/X sky130_fd_sc_hd__clkbuf_2
X_22559_ _22559_/A vssd1 vssd1 vccd1 vccd1 _22771_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13782__A2 _15008_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20647__A4 _20928_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15100_ _15100_/A _15100_/B vssd1 vssd1 vccd1 vccd1 _15101_/B sky130_fd_sc_hd__and2_2
X_12312_ _12401_/A _12822_/A _12385_/A _12409_/A vssd1 vssd1 vccd1 vccd1 _16256_/D
+ sky130_fd_sc_hd__a31o_2
XFILLER_177_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16080_ _16080_/A _16080_/B _16080_/C vssd1 vssd1 vccd1 vccd1 _16081_/B sky130_fd_sc_hd__and3_1
X_13292_ _22730_/Q vssd1 vssd1 vccd1 vccd1 _21188_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input78_A x[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12243_ _18249_/B vssd1 vssd1 vccd1 vccd1 _12249_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15031_ _15031_/A _15031_/B _15088_/B vssd1 vssd1 vccd1 vccd1 _15033_/A sky130_fd_sc_hd__and3_1
XFILLER_177_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11545__A1 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20804__A1 _20844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ _11500_/Y _11636_/A _12167_/X _12156_/A _12172_/Y vssd1 vssd1 vccd1 vccd1
+ _12174_/X sky130_fd_sc_hd__o311a_2
XFILLER_150_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15484__A _15484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19770_ _19836_/D _19836_/A _19350_/X _17819_/A vssd1 vssd1 vccd1 vccd1 _19782_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16982_ _16982_/A _17188_/A _17188_/B vssd1 vssd1 vccd1 vccd1 _16982_/Y sky130_fd_sc_hd__nand3_1
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16299__B _20678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18721_ _18721_/A _18721_/B vssd1 vssd1 vccd1 vccd1 _18723_/B sky130_fd_sc_hd__nand2_1
X_15933_ _15933_/A vssd1 vssd1 vccd1 vccd1 _15934_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18795__A _18795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18652_ _15981_/X _11786_/X _18508_/A _18508_/B vssd1 vssd1 vccd1 vccd1 _18653_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _15864_/A _15864_/B _15864_/C _15864_/D vssd1 vssd1 vccd1 vccd1 _15952_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16787__A2 _17634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _17603_/A _17603_/B _17603_/C _17603_/D vssd1 vssd1 vccd1 vccd1 _17603_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_97_1038 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14815_ _14815_/A _14815_/B _14815_/C vssd1 vssd1 vccd1 vccd1 _14816_/B sky130_fd_sc_hd__nand3_1
X_18583_ _18774_/C _18774_/D vssd1 vssd1 vccd1 vccd1 _18586_/C sky130_fd_sc_hd__and2_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _12606_/X _12607_/X _15891_/A vssd1 vssd1 vccd1 vccd1 _15795_/X sky130_fd_sc_hd__a21o_1
XFILLER_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _16225_/X _16227_/X _17401_/D _15960_/A vssd1 vssd1 vccd1 vccd1 _17535_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_33_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _14745_/B _14745_/C _14745_/A vssd1 vssd1 vccd1 vccd1 _14747_/C sky130_fd_sc_hd__a21o_1
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11958_ _11938_/Y _11956_/Y _18292_/A _11731_/A vssd1 vssd1 vccd1 vccd1 _11958_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_33_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17465_ _17083_/X _17728_/A _17463_/X _17285_/Y _17464_/Y vssd1 vssd1 vccd1 vccd1
+ _17467_/A sky130_fd_sc_hd__o311ai_4
XANTENNA__16944__C1 _19199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14677_ _14675_/Y _14676_/X _14560_/A _14057_/X vssd1 vssd1 vccd1 vccd1 _14677_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_189_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11889_ _16103_/D vssd1 vssd1 vccd1 vccd1 _16157_/D sky130_fd_sc_hd__clkbuf_4
X_19204_ _18371_/A _17400_/A _17393_/X _12018_/X vssd1 vssd1 vccd1 vccd1 _19418_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_60_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16416_ _16419_/A _16421_/C vssd1 vssd1 vccd1 vccd1 _16417_/C sky130_fd_sc_hd__nand2_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19489__A1 _11639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13628_ _13627_/A _13627_/B _13627_/C vssd1 vssd1 vccd1 vccd1 _13643_/B sky130_fd_sc_hd__a21o_1
X_17396_ _15934_/A _17822_/A _17408_/A vssd1 vssd1 vccd1 vccd1 _17399_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__13222__A1 _13475_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19135_ _19138_/D _19138_/B _19138_/C vssd1 vssd1 vccd1 vccd1 _19136_/A sky130_fd_sc_hd__nand3_1
XFILLER_146_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20099__A2 _16261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18680__D _18680_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16347_ _20357_/C vssd1 vssd1 vccd1 vccd1 _20582_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__18697__C1 _18678_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13559_ _13559_/A _13559_/B _13559_/C vssd1 vssd1 vccd1 vccd1 _13677_/A sky130_fd_sc_hd__nand3_1
XFILLER_145_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18161__A1 _12164_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19066_ _11308_/A _11308_/B _19046_/A _19065_/X _17819_/A vssd1 vssd1 vccd1 vccd1
+ _19066_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_2_0_bq_clk_i clkbuf_2_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16278_ _16595_/A _16596_/A _16273_/X _16277_/X vssd1 vssd1 vccd1 vccd1 _16283_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18017_ _18017_/A vssd1 vssd1 vccd1 vccd1 _22965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17874__A _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15229_ _15210_/A _15210_/B _15197_/X _15227_/X vssd1 vssd1 vccd1 vccd1 _15230_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16475__A1 _16248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22668__CLK _22964_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15394__A _15394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19968_ _19977_/A _19977_/B _22924_/Q vssd1 vssd1 vccd1 vccd1 _19974_/C sky130_fd_sc_hd__nand3_1
XFILLER_114_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18919_ _19091_/B _18920_/B _18871_/Y _18900_/A _18908_/C vssd1 vssd1 vccd1 vccd1
+ _18919_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_80_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19899_ _19899_/A _19899_/B _19937_/A _19899_/D vssd1 vssd1 vccd1 vccd1 _19937_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12530__B _12773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18621__C1 _17632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21930_ _21930_/A vssd1 vssd1 vccd1 vccd1 _22155_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16937__B _16937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21861_ _21990_/A _21963_/A _21990_/C vssd1 vssd1 vccd1 vccd1 _21861_/X sky130_fd_sc_hd__and3_1
XFILLER_103_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20812_ _20812_/A _20812_/B _20812_/C _20812_/D vssd1 vssd1 vccd1 vccd1 _20812_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21792_ _21783_/X _21785_/Y _21789_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _21792_/X
+ sky130_fd_sc_hd__o211a_2
XANTENNA__14457__B _22876_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20743_ _20928_/C vssd1 vssd1 vccd1 vccd1 _21050_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_168_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20674_ _16294_/X _16293_/X _20853_/A _20608_/B vssd1 vssd1 vccd1 vccd1 _20676_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_196_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22413_ _22707_/Q input45/X _22413_/S vssd1 vssd1 vccd1 vccd1 _22414_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15569__A _15569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22344_ _22684_/Q _22289_/B _22324_/B vssd1 vssd1 vccd1 vccd1 _22344_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19983__B _19983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15505__A3 _17427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15910__B1 _15792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22275_ _22240_/A _22240_/B _22240_/C vssd1 vssd1 vccd1 vccd1 _22277_/B sky130_fd_sc_hd__a21boi_1
XFILLER_191_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20247__C1 _16932_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21226_ _22057_/B _21219_/C _21227_/B vssd1 vssd1 vccd1 vccd1 _21226_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18455__A2 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22840__D _22852_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16466__A1 _12118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16466__B2 _12696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21157_ _22947_/Q _21157_/B vssd1 vssd1 vccd1 vccd1 _21162_/B sky130_fd_sc_hd__xor2_4
XFILLER_105_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12721__A _12721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22539__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20108_ _20119_/A _20118_/B _20119_/B vssd1 vssd1 vccd1 vccd1 _20115_/A sky130_fd_sc_hd__nand3_2
XFILLER_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21088_ _21088_/A _21088_/B vssd1 vssd1 vccd1 vccd1 _21090_/C sky130_fd_sc_hd__xnor2_1
XFILLER_101_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20039_ _18778_/D _19987_/B _20013_/X _20037_/B _20012_/X vssd1 vssd1 vccd1 vccd1
+ _20039_/Y sky130_fd_sc_hd__o221ai_1
XANTENNA__19504__A _19504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12930_ _12930_/A vssd1 vssd1 vccd1 vccd1 _16155_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__18612__C1 _19197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_856 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12861_ _20120_/B _12860_/Y _12851_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12862_/A
+ sky130_fd_sc_hd__o211ai_2
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14600_ _14600_/A _14600_/B _14600_/C vssd1 vssd1 vccd1 vccd1 _14600_/Y sky130_fd_sc_hd__nand3_2
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11630_/Y _11807_/Y _11592_/A vssd1 vssd1 vccd1 vccd1 _11930_/A sky130_fd_sc_hd__o21a_1
X_15580_ _15580_/A vssd1 vssd1 vccd1 vccd1 _15580_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12792_/A _12792_/B _12792_/C _12792_/D vssd1 vssd1 vccd1 vccd1 _12792_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14272_/C _14044_/B _14527_/Y _13957_/A _14528_/Y vssd1 vssd1 vccd1 vccd1
+ _14561_/B sky130_fd_sc_hd__a221oi_4
X_11743_ _11436_/A _11721_/C _11438_/B vssd1 vssd1 vccd1 vccd1 _11905_/A sky130_fd_sc_hd__a21boi_4
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17250_ _17145_/B _17247_/X _17257_/B _17249_/Y vssd1 vssd1 vccd1 vccd1 _17255_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14462_ _14770_/A _14771_/A _14785_/B _14808_/A _14693_/B vssd1 vssd1 vccd1 vccd1
+ _14462_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_53_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11674_ _11674_/A _11932_/C _11673_/X vssd1 vssd1 vccd1 vccd1 _12083_/B sky130_fd_sc_hd__nor3b_4
XFILLER_168_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19596__D _19774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16201_ _16201_/A _16201_/B _16201_/C vssd1 vssd1 vccd1 vccd1 _16202_/B sky130_fd_sc_hd__nand3_1
X_13413_ _13413_/A _13413_/B vssd1 vssd1 vccd1 vccd1 _21270_/C sky130_fd_sc_hd__and2_1
X_17181_ _17181_/A _17181_/B vssd1 vssd1 vccd1 vccd1 _17181_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15479__A _15479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14393_ _22706_/Q _14370_/X _14379_/X _22738_/Q _14392_/X vssd1 vssd1 vccd1 vccd1
+ _14393_/X sky130_fd_sc_hd__a221o_1
XFILLER_183_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18143__A1 _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16132_ _16072_/X _16084_/Y _16085_/Y _16086_/Y vssd1 vssd1 vccd1 vccd1 _16132_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__11800__A _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13344_ _13344_/A vssd1 vssd1 vccd1 vccd1 _13344_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_127_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18694__A2 _19160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ _16191_/A _16080_/A _16080_/C _16586_/B vssd1 vssd1 vccd1 vccd1 _16064_/B
+ sky130_fd_sc_hd__nand4_1
X_13275_ _13229_/A _13361_/A _13274_/Y vssd1 vssd1 vccd1 vccd1 _13275_/X sky130_fd_sc_hd__o21a_1
XFILLER_182_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15014_ _15080_/A _15080_/B _15080_/C vssd1 vssd1 vccd1 vccd1 _15015_/C sky130_fd_sc_hd__o21ai_1
X_12226_ _18228_/A _18228_/B _18227_/C vssd1 vssd1 vccd1 vccd1 _12227_/C sky130_fd_sc_hd__nand3_1
XFILLER_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19822_ _19822_/A _22921_/Q _19822_/C vssd1 vssd1 vccd1 vccd1 _19890_/A sky130_fd_sc_hd__nand3_2
XANTENNA__18997__A3 _18890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13727__A _13727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _12157_/A vssd1 vssd1 vccd1 vccd1 _12157_/X sky130_fd_sc_hd__buf_2
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12631__A _16488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16103__A _20390_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21944__A _21944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19753_ _20025_/A _19749_/X _19752_/Y vssd1 vssd1 vccd1 vccd1 _19754_/B sky130_fd_sc_hd__o21a_1
X_16965_ _16946_/X _16948_/X _16956_/Y _20249_/C _19504_/B vssd1 vssd1 vccd1 vccd1
+ _16967_/C sky130_fd_sc_hd__o2111ai_1
X_12088_ _12088_/A _12088_/B vssd1 vssd1 vccd1 vccd1 _12089_/B sky130_fd_sc_hd__nand2_1
XANTENNA__22960__CLK _22964_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__D _18305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15916_ _15915_/A _15915_/B _15793_/Y _15794_/X vssd1 vssd1 vccd1 vccd1 _15916_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_18704_ _18343_/X _18695_/X _11800_/X _18333_/X vssd1 vssd1 vccd1 vccd1 _18705_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_110_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19684_ _19684_/A _19684_/B _19684_/C vssd1 vssd1 vccd1 vccd1 _19684_/X sky130_fd_sc_hd__and3_1
X_16896_ _16444_/A _16894_/Y _16895_/Y _16650_/C vssd1 vssd1 vccd1 vccd1 _16896_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_64_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18635_ _18625_/X _18627_/Y _18629_/Y vssd1 vssd1 vccd1 vccd1 _18635_/X sky130_fd_sc_hd__o21ba_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _15845_/X _15846_/Y _15854_/B vssd1 vssd1 vccd1 vccd1 _15847_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18566_ _18568_/B _18568_/C _18568_/A vssd1 vssd1 vccd1 vccd1 _18569_/A sky130_fd_sc_hd__a21o_1
XFILLER_18_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17709__A1 _17226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _15780_/A _15779_/A vssd1 vssd1 vccd1 vccd1 _15778_/Y sky130_fd_sc_hd__nand2_2
XFILLER_45_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17517_ _17603_/A _17603_/C vssd1 vssd1 vccd1 vccd1 _17518_/B sky130_fd_sc_hd__nor2_1
XFILLER_178_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14729_ _14729_/A _14729_/B vssd1 vssd1 vccd1 vccd1 _14729_/Y sky130_fd_sc_hd__nand2_1
X_18497_ _18340_/B _18482_/Y _18705_/A _16564_/B _19694_/D vssd1 vssd1 vccd1 vccd1
+ _18499_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18691__C _18691_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17448_ _17426_/A _17882_/C _19619_/D _16124_/X _20917_/B vssd1 vssd1 vccd1 vccd1
+ _17449_/D sky130_fd_sc_hd__a32o_1
XFILLER_21_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15389__A _15389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17379_ _17379_/A vssd1 vssd1 vccd1 vccd1 _17388_/A sky130_fd_sc_hd__buf_4
XFILLER_174_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_931 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19331__B1 _19167_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19118_ _18932_/A _18932_/B _18932_/C _18935_/Y vssd1 vssd1 vccd1 vccd1 _19118_/X
+ sky130_fd_sc_hd__a31o_1
X_20390_ _20264_/A _20390_/B _20390_/C _20390_/D vssd1 vssd1 vccd1 vccd1 _20393_/A
+ sky130_fd_sc_hd__nand4b_2
XFILLER_173_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18685__A2 _19687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12525__B _12525_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14156__C1 _14147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19049_ _18797_/Y _19357_/A _18282_/X _19048_/Y vssd1 vssd1 vccd1 vccd1 _19062_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_146_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22060_ _22062_/A _22262_/A _22190_/D _22059_/Y vssd1 vssd1 vccd1 vccd1 _22060_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_126_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16448__A1 _15335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21011_ _21011_/A _21011_/B _21011_/C vssd1 vssd1 vccd1 vccd1 _21081_/C sky130_fd_sc_hd__and3_1
XANTENNA__20461__C _20461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21441__A1 _21440_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22962_ _22964_/CLK _22962_/D vssd1 vssd1 vccd1 vccd1 _22962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11693__B1 _11566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21913_ _21913_/A _21913_/B vssd1 vssd1 vccd1 vccd1 _21913_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22893_ _22951_/CLK _22893_/D vssd1 vssd1 vccd1 vccd1 _22893_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21844_ _13344_/X _13345_/X _22167_/A vssd1 vssd1 vccd1 vccd1 _21897_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21775_ _21766_/B _21730_/A _21742_/A _21607_/X vssd1 vssd1 vccd1 vccd1 _21775_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_168_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19697__C _19774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19570__B1 _22918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20917__B _20917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20726_ _16267_/X _16266_/X _20449_/A _16268_/X vssd1 vssd1 vccd1 vccd1 _20726_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15187__B2 _14942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22835__D _22847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15299__A _16256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20657_ _20543_/Y _20539_/Y _20652_/Y _20551_/Y _20660_/A vssd1 vssd1 vccd1 vccd1
+ _20827_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_177_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12716__A _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22833__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11390_ _15484_/A _11325_/A _11325_/B _11311_/Y vssd1 vssd1 vccd1 vccd1 _18482_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__20355__D _20355_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20588_ _20581_/A _16344_/A _20584_/C _20587_/Y vssd1 vssd1 vccd1 vccd1 _20704_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_137_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16687__A1 _16669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22327_ _22327_/A _22327_/B vssd1 vssd1 vccd1 vccd1 _22328_/A sky130_fd_sc_hd__or2_1
XFILLER_164_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21748__B _21757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12154__C _12154_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ _13096_/A _21307_/C _13095_/A vssd1 vssd1 vccd1 vccd1 _13138_/C sky130_fd_sc_hd__nand3_1
X_22258_ _22258_/A _22258_/B _22258_/C vssd1 vssd1 vccd1 vccd1 _22300_/B sky130_fd_sc_hd__nand3_1
XFILLER_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15746__B _15746_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12011_ _12009_/X _19350_/A _11984_/A vssd1 vssd1 vccd1 vccd1 _12013_/A sky130_fd_sc_hd__o21ai_1
X_21209_ _13324_/B _13300_/Y _13317_/X _13316_/X vssd1 vssd1 vccd1 vccd1 _21210_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22189_ _22231_/C _22231_/B vssd1 vssd1 vccd1 vccd1 _22219_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16750_ _16733_/Y _16740_/Y _16853_/A vssd1 vssd1 vccd1 vccd1 _16754_/A sky130_fd_sc_hd__o21ai_1
XFILLER_98_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13962_ _22762_/Q vssd1 vssd1 vccd1 vccd1 _14581_/B sky130_fd_sc_hd__inv_2
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21196__B1 _22841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15701_ _20678_/B vssd1 vssd1 vccd1 vccd1 _17525_/C sky130_fd_sc_hd__buf_4
XANTENNA__15481__B _22660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ _12913_/A _20972_/D vssd1 vssd1 vccd1 vccd1 _12958_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16681_ _17502_/A _16426_/X _16683_/B _16683_/C vssd1 vssd1 vccd1 vccd1 _16681_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_24_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13893_ _13907_/A vssd1 vssd1 vccd1 vccd1 _14583_/C sky130_fd_sc_hd__buf_2
XFILLER_19_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14378__A _16324_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15912__D _17407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18420_ _18417_/C _18417_/A _18219_/B vssd1 vssd1 vccd1 vccd1 _18423_/A sky130_fd_sc_hd__a21o_1
XFILLER_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15632_ _12378_/B _15631_/X _11627_/A _15633_/B vssd1 vssd1 vccd1 vccd1 _15632_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_686 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _12844_/A vssd1 vssd1 vccd1 vccd1 _16178_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _18351_/A _18351_/B _18351_/C vssd1 vssd1 vccd1 vccd1 _18355_/B sky130_fd_sc_hd__nand3_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15563_ _12844_/A _16274_/A _15557_/Y vssd1 vssd1 vccd1 vccd1 _15563_/Y sky130_fd_sc_hd__o21ai_2
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12772_/X _12774_/X _22826_/Q _12645_/A _12769_/Y vssd1 vssd1 vccd1 vccd1
+ _12776_/A sky130_fd_sc_hd__o2111a_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17334_/A vssd1 vssd1 vccd1 vccd1 _17486_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20827__B _20827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14515_/B _14515_/C _14515_/A vssd1 vssd1 vccd1 vccd1 _14516_/B sky130_fd_sc_hd__a21o_1
XFILLER_70_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18282_ _18282_/A vssd1 vssd1 vccd1 vccd1 _18282_/X sky130_fd_sc_hd__clkbuf_2
X_11726_ _11940_/A vssd1 vssd1 vccd1 vccd1 _16256_/A sky130_fd_sc_hd__buf_4
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15494_ _17379_/A _12719_/A _15498_/A _15567_/A _15567_/B vssd1 vssd1 vccd1 vccd1
+ _15500_/A sky130_fd_sc_hd__o311a_1
XFILLER_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17233_ _17178_/Y _17173_/D _17173_/C vssd1 vssd1 vccd1 vccd1 _17301_/A sky130_fd_sc_hd__a21boi_1
XFILLER_80_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14445_ _16400_/C vssd1 vssd1 vccd1 vccd1 _16879_/B sky130_fd_sc_hd__buf_2
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11657_ _15539_/A _15435_/C vssd1 vssd1 vccd1 vccd1 _11737_/A sky130_fd_sc_hd__nand2_4
XFILLER_31_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11739__A1 _11625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17164_ _17158_/A _17158_/B _17162_/Y _17163_/X vssd1 vssd1 vccd1 vccd1 _17164_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__16127__B1 _12765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14376_ _22702_/Q _14370_/X _14351_/X _22734_/Q _14375_/X vssd1 vssd1 vccd1 vccd1
+ _14376_/X sky130_fd_sc_hd__a221o_1
X_11588_ _18348_/A vssd1 vssd1 vccd1 vccd1 _15988_/A sky130_fd_sc_hd__buf_4
XANTENNA__20622__B1_N _20626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20843__A _20843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16115_ _16053_/X _15997_/X _16110_/B _15972_/X _16055_/Y vssd1 vssd1 vccd1 vccd1
+ _16115_/X sky130_fd_sc_hd__o2111a_1
X_13327_ _13099_/B _13098_/A _13095_/A _13326_/Y vssd1 vssd1 vccd1 vccd1 _13332_/C
+ sky130_fd_sc_hd__a31oi_4
X_17095_ _19615_/C _17739_/A _16810_/C _16816_/Y vssd1 vssd1 vccd1 vccd1 _17095_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_116_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16046_ _16046_/A vssd1 vssd1 vccd1 vccd1 _16047_/B sky130_fd_sc_hd__buf_2
XANTENNA__19616__A1 _11821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13258_ _13662_/B _13662_/C vssd1 vssd1 vccd1 vccd1 _13370_/A sky130_fd_sc_hd__nand2_2
XANTENNA__20007__B1_N _22925_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12209_ _12209_/A vssd1 vssd1 vccd1 vccd1 _17380_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13189_ _13450_/C vssd1 vssd1 vccd1 vccd1 _21173_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19805_ _19731_/A _19731_/B _19735_/C _19804_/X vssd1 vssd1 vccd1 vccd1 _19806_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17997_ _17997_/A _18020_/D vssd1 vssd1 vccd1 vccd1 _17999_/A sky130_fd_sc_hd__xnor2_2
XFILLER_69_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19736_ _19736_/A _19736_/B _19736_/C vssd1 vssd1 vccd1 vccd1 _19808_/A sky130_fd_sc_hd__nand3_2
X_16948_ _17145_/A vssd1 vssd1 vccd1 vccd1 _16948_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15391__B _15665_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19667_ _19813_/A _19813_/B _19666_/X vssd1 vssd1 vccd1 vccd1 _19670_/A sky130_fd_sc_hd__a21o_1
X_16879_ _16879_/A _16879_/B _17840_/A vssd1 vssd1 vccd1 vccd1 _16879_/X sky130_fd_sc_hd__and3_1
XFILLER_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18618_ _18618_/A _18618_/B vssd1 vssd1 vccd1 vccd1 _18618_/Y sky130_fd_sc_hd__nand2_1
X_19598_ _19684_/A _19684_/B _19684_/C vssd1 vssd1 vccd1 vccd1 _19598_/Y sky130_fd_sc_hd__nand3_1
XFILLER_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18549_ _18519_/Y _18523_/Y _18527_/Y _18557_/A vssd1 vssd1 vccd1 vccd1 _18556_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_127_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22856__CLK _22937_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21560_ _21560_/A _21560_/B vssd1 vssd1 vccd1 vccd1 _21561_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20456__C _20456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20511_ _20511_/A _20511_/B _20511_/C _20511_/D vssd1 vssd1 vccd1 vccd1 _20519_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_127_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21491_ _21467_/A _21467_/B _21323_/Y vssd1 vssd1 vccd1 vccd1 _21504_/A sky130_fd_sc_hd__a21oi_2
XFILLER_20_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11440__A _15633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20442_ _20442_/A _20442_/B vssd1 vssd1 vccd1 vccd1 _20754_/A sky130_fd_sc_hd__nand2_2
XFILLER_146_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20465__A2 _16745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20373_ _20236_/B _20236_/C _20363_/Y vssd1 vssd1 vccd1 vccd1 _20375_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12942__A3 _20584_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22112_ _21853_/X _21970_/X _22111_/Y vssd1 vssd1 vccd1 vccd1 _22113_/C sky130_fd_sc_hd__o21ai_1
XFILLER_161_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15892__A2 _12774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22043_ _21960_/Y _22040_/Y _21963_/A _22042_/Y _22176_/A vssd1 vssd1 vccd1 vccd1
+ _22044_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_47_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22611__A0 _18127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14447__A3 _22967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15644__A2 _15630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13814__B _13814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22945_ _22948_/CLK _22945_/D vssd1 vssd1 vccd1 vccd1 _22945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14629__C _14911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22876_ _22916_/CLK _22876_/D vssd1 vssd1 vccd1 vccd1 _22876_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22619__S _22619_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20928__A _20928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21827_ _21562_/Y _21707_/X _21708_/X vssd1 vssd1 vccd1 vccd1 _21827_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__21750__C _21750_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12560_ _12645_/A _12645_/C vssd1 vssd1 vccd1 vccd1 _12560_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12091__B1 _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21758_ _21758_/A _21758_/B _21758_/C _21758_/D vssd1 vssd1 vccd1 vccd1 _21760_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18117__B _18128_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_1066 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11511_ _11511_/A vssd1 vssd1 vccd1 vccd1 _11511_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__14368__C1 _14367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20709_ _20709_/A _20709_/B _20709_/C vssd1 vssd1 vccd1 vccd1 _20720_/C sky130_fd_sc_hd__nand3_1
XFILLER_196_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12491_ _12358_/X _12488_/Y _12432_/A vssd1 vssd1 vccd1 vccd1 _12508_/A sky130_fd_sc_hd__o21ai_1
XFILLER_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21689_ _21689_/A vssd1 vssd1 vccd1 vccd1 _22167_/A sky130_fd_sc_hd__buf_2
X_14230_ _14230_/A vssd1 vssd1 vccd1 vccd1 _15050_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_137_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11442_ _18682_/C vssd1 vssd1 vccd1 vccd1 _15415_/C sky130_fd_sc_hd__buf_2
XANTENNA__16109__B1 _16613_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18649__A2 _12158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21102__B1 _22942_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19310__A3 _19481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14161_ _14272_/C _14161_/B _14161_/C _14494_/C vssd1 vssd1 vccd1 vccd1 _14161_/X
+ sky130_fd_sc_hd__and4_1
X_11373_ _22784_/Q vssd1 vssd1 vccd1 vccd1 _11450_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input60_A wb_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ _13143_/A _13143_/B _13112_/C _13112_/D vssd1 vssd1 vccd1 vccd1 _13112_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_152_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19059__C1 _19351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15476__B _20133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14092_ _14054_/Y _14055_/X _14089_/Y _14091_/X vssd1 vssd1 vccd1 vccd1 _14094_/A
+ sky130_fd_sc_hd__o31ai_2
XFILLER_153_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22602__A0 _11980_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17920_ _17920_/A vssd1 vssd1 vccd1 vccd1 _17920_/Y sky130_fd_sc_hd__inv_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _20182_/A _13043_/B _20182_/B vssd1 vssd1 vccd1 vccd1 _13044_/B sky130_fd_sc_hd__nand3_1
XFILLER_106_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17851_ _17800_/Y _17849_/Y _18048_/C _22902_/Q vssd1 vssd1 vccd1 vccd1 _17851_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_67_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18821__A2 _19334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16802_ _16544_/Y _16542_/Y _16524_/Y _16512_/Y vssd1 vssd1 vccd1 vccd1 _16908_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17782_ _17704_/B _17780_/X _17781_/Y _17605_/A vssd1 vssd1 vccd1 vccd1 _17787_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14994_ _15004_/D _15115_/A _15115_/B _15062_/A _15050_/B vssd1 vssd1 vccd1 vccd1
+ _14996_/C sky130_fd_sc_hd__a32o_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19521_ _19521_/A _19581_/A _19521_/C _19521_/D vssd1 vssd1 vccd1 vccd1 _19525_/A
+ sky130_fd_sc_hd__nand4_1
X_16733_ _16723_/X _16726_/Y _16732_/Y vssd1 vssd1 vccd1 vccd1 _16733_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _14613_/A vssd1 vssd1 vccd1 vccd1 _15058_/C sky130_fd_sc_hd__buf_2
XFILLER_93_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16100__B _19000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19452_ _19452_/A _19452_/B vssd1 vssd1 vccd1 vccd1 _22897_/D sky130_fd_sc_hd__xor2_1
XANTENNA__22879__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__A _18482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16664_ _16664_/A _16664_/B _16664_/C vssd1 vssd1 vccd1 vccd1 _16665_/A sky130_fd_sc_hd__nand3_2
XANTENNA__21941__B _22062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13876_ _13876_/A _14722_/A vssd1 vssd1 vccd1 vccd1 _13877_/B sky130_fd_sc_hd__nand2_1
XANTENNA__20392__A1 _12500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18403_ _18571_/D _18442_/B _18442_/C vssd1 vssd1 vccd1 vccd1 _18403_/X sky130_fd_sc_hd__and3_1
X_15615_ _18706_/A _16715_/A _20098_/D _16304_/A _18875_/C vssd1 vssd1 vccd1 vccd1
+ _15616_/A sky130_fd_sc_hd__a32oi_4
XFILLER_90_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19383_ _19457_/A _19389_/B _19389_/C vssd1 vssd1 vccd1 vccd1 _19398_/C sky130_fd_sc_hd__a21o_1
X_12827_ _15370_/B vssd1 vssd1 vccd1 vccd1 _12827_/X sky130_fd_sc_hd__buf_4
XFILLER_62_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16595_ _16595_/A _16595_/B vssd1 vssd1 vccd1 vccd1 _16596_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18334_ _11636_/A _11786_/X _15358_/X _18333_/X vssd1 vssd1 vccd1 vccd1 _18529_/A
+ sky130_fd_sc_hd__o22ai_4
X_15546_ _15546_/A vssd1 vssd1 vccd1 vccd1 _15546_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12758_/A vssd1 vssd1 vccd1 vccd1 _12988_/A sky130_fd_sc_hd__buf_4
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18265_ _18088_/Y _18252_/Y _18262_/Y _18268_/A vssd1 vssd1 vccd1 vccd1 _18266_/B
+ sky130_fd_sc_hd__a31o_1
X_11709_ _16257_/B _11709_/B _16257_/A vssd1 vssd1 vccd1 vccd1 _11938_/A sky130_fd_sc_hd__nand3_1
X_15477_ _15477_/A _15477_/B vssd1 vssd1 vccd1 vccd1 _15479_/B sky130_fd_sc_hd__nand2_1
X_12689_ _12689_/A _17401_/B _12689_/C vssd1 vssd1 vccd1 vccd1 _12689_/X sky130_fd_sc_hd__and3_1
XANTENNA__12356__A _15633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17216_ _17370_/A _17370_/B _17215_/Y _17373_/A vssd1 vssd1 vccd1 vccd1 _17219_/A
+ sky130_fd_sc_hd__a22oi_2
X_14428_ _22719_/Q _14418_/X _14351_/A _22751_/Q _14427_/X vssd1 vssd1 vccd1 vccd1
+ _14428_/X sky130_fd_sc_hd__a221o_2
X_18196_ _15530_/X _15531_/X _11634_/A vssd1 vssd1 vccd1 vccd1 _18197_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__14374__A2 _14370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_506 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17147_ _17138_/A _17142_/A _17145_/Y vssd1 vssd1 vccd1 vccd1 _17149_/A sky130_fd_sc_hd__o21ai_1
XFILLER_156_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14359_ _22731_/Q vssd1 vssd1 vccd1 vccd1 _14359_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17078_ _17078_/A _17078_/B vssd1 vssd1 vccd1 vccd1 _17078_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16029_ _16133_/A vssd1 vssd1 vccd1 vccd1 _16093_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18273__B1 _12251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18812__A2 _11503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16498__A _16498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21554__D _21556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18025__B1 _18778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__A2_N _18875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19719_ _19788_/B _19719_/B vssd1 vssd1 vccd1 vccd1 _19719_/X sky130_fd_sc_hd__or2_1
XANTENNA__11648__B1 _11635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20991_ _20892_/A _20908_/Y _20952_/A _20894_/B vssd1 vssd1 vccd1 vccd1 _20992_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_72_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1120 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19773__B1 _19624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22730_ _22731_/CLK _22730_/D vssd1 vssd1 vccd1 vccd1 _22730_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21851__B _22041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22439__S _22439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14598__C1 _13873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22661_ _22661_/A vssd1 vssd1 vccd1 vccd1 _22950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21612_ _21383_/X _21606_/X _21766_/A vssd1 vssd1 vccd1 vccd1 _21645_/C sky130_fd_sc_hd__o21ai_1
XFILLER_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18879__A2 _15905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22592_ _22592_/A vssd1 vssd1 vccd1 vccd1 _22785_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12612__A2 _15569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21543_ _21547_/A _21547_/B _21531_/X _21534_/Y _21546_/A vssd1 vssd1 vccd1 vccd1
+ _21553_/B sky130_fd_sc_hd__o221ai_4
XANTENNA__12266__A _22703_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_856 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15562__A1 _11704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21474_ _21307_/B _21307_/A _21473_/Y vssd1 vssd1 vccd1 vccd1 _21749_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__15562__B2 _16778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19694__D _19694_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12376__A1 _12343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15577__A _19012_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20425_ _20549_/B _20432_/B _20422_/Y _20424_/Y vssd1 vssd1 vccd1 vccd1 _20554_/A
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_146_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20356_ _12721_/A _15412_/A _20370_/D vssd1 vssd1 vccd1 vccd1 _20511_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__16511__B1 _16964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20287_ _20269_/X _20274_/Y _20401_/A _20401_/B vssd1 vssd1 vccd1 vccd1 _20290_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_115_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20930__B _21017_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22026_ _21917_/Y _21836_/Y _22025_/Y vssd1 vssd1 vccd1 vccd1 _22026_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18264__B1 _18088_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22060__A1 _22062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_620 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11991_ _22792_/Q _11783_/A _12107_/C _11783_/C vssd1 vssd1 vccd1 vccd1 _18140_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_60_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19512__A _19512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13730_ _22757_/Q vssd1 vssd1 vccd1 vccd1 _13963_/D sky130_fd_sc_hd__clkinv_2
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22928_ _22949_/CLK _22928_/D vssd1 vssd1 vccd1 vccd1 _22928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20374__A1 _20511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16578__B1 _11845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_639 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13661_ _13660_/A _13659_/B _13624_/B vssd1 vssd1 vccd1 vccd1 _13665_/A sky130_fd_sc_hd__a21bo_1
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22859_ _22916_/CLK _22859_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15400_ _16257_/D vssd1 vssd1 vccd1 vccd1 _20502_/B sky130_fd_sc_hd__buf_2
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12450_/X _15569_/A _12424_/Y _15450_/A _12595_/Y vssd1 vssd1 vccd1 vccd1
+ _12612_/Y sky130_fd_sc_hd__o221ai_4
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _16366_/Y _16370_/Y _16374_/Y vssd1 vssd1 vccd1 vccd1 _16391_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20126__A1 _15355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _13461_/B _13521_/Y _21874_/A _13528_/X _21445_/C vssd1 vssd1 vccd1 vccd1
+ _13597_/B sky130_fd_sc_hd__o2111ai_1
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15331_ _15893_/A _15901_/B _20133_/A _16781_/B vssd1 vssd1 vccd1 vccd1 _15331_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_12_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12543_ _12543_/A _12543_/B _12543_/C _12543_/D vssd1 vssd1 vccd1 vccd1 _12561_/A
+ sky130_fd_sc_hd__nand4_2
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17542__A2 _20870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18050_ _18045_/Y _18048_/X _18049_/Y vssd1 vssd1 vccd1 vccd1 _18051_/C sky130_fd_sc_hd__o21ai_1
X_15262_ _15262_/A _15262_/B vssd1 vssd1 vccd1 vccd1 _15263_/B sky130_fd_sc_hd__nand2_1
XANTENNA__21489__A _21489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19819__A1 _18246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ _12470_/X _12669_/A _12528_/A _16328_/A _16319_/C vssd1 vssd1 vccd1 vccd1
+ _12500_/A sky130_fd_sc_hd__o311a_2
XFILLER_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16750__B1 _16853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17001_ _17001_/A _17001_/B _17001_/C vssd1 vssd1 vccd1 vccd1 _17006_/B sky130_fd_sc_hd__nand3_2
X_14213_ _14765_/A _14779_/A _14765_/C _14595_/B _14222_/A vssd1 vssd1 vccd1 vccd1
+ _14265_/B sky130_fd_sc_hd__a32o_1
XFILLER_172_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ _12170_/A _12171_/A _18682_/C vssd1 vssd1 vccd1 vccd1 _11425_/Y sky130_fd_sc_hd__o21ai_4
X_15193_ _15186_/X _15187_/X _15194_/C _15216_/A vssd1 vssd1 vccd1 vccd1 _15197_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15305__A1 _15298_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ _14085_/A _13808_/A _14619_/A _14143_/X _13829_/Y vssd1 vssd1 vccd1 vccd1
+ _14146_/B sky130_fd_sc_hd__o221ai_1
X_11356_ _11434_/A vssd1 vssd1 vccd1 vccd1 _15484_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_180_550 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12119__A1 _12116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12119__B2 _16016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18952_ _18952_/A _18952_/B _18952_/C vssd1 vssd1 vccd1 vccd1 _18955_/B sky130_fd_sc_hd__nand3_1
XFILLER_140_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14075_ _13819_/Y _13829_/Y _14619_/A _14576_/A vssd1 vssd1 vccd1 vccd1 _14075_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
X_11287_ _22954_/Q vssd1 vssd1 vccd1 vccd1 _11404_/B sky130_fd_sc_hd__buf_2
XFILLER_106_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17903_ _17949_/B vssd1 vssd1 vccd1 vccd1 _17919_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__11743__B1_N _11438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13026_ _16157_/C _13016_/C _13024_/A _13024_/B vssd1 vssd1 vccd1 vccd1 _13026_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18883_ _18883_/A _18883_/B _18883_/C vssd1 vssd1 vccd1 vccd1 _18901_/A sky130_fd_sc_hd__nand3_1
XFILLER_117_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17834_ _19901_/D _17872_/C _17833_/X _17753_/B vssd1 vssd1 vccd1 vccd1 _17871_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_120_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17765_ _17765_/A _17765_/B _17763_/X vssd1 vssd1 vccd1 vccd1 _17768_/C sky130_fd_sc_hd__nor3b_1
XFILLER_19_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14977_ _14977_/A _14977_/B _15035_/A vssd1 vssd1 vccd1 vccd1 _15035_/B sky130_fd_sc_hd__nand3_2
XFILLER_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19504_ _19504_/A _19504_/B _19504_/C _19504_/D vssd1 vssd1 vccd1 vccd1 _19652_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16716_ _20101_/B vssd1 vssd1 vccd1 vccd1 _20781_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__21671__B _21677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13928_ _14069_/A vssd1 vssd1 vccd1 vccd1 _14765_/A sky130_fd_sc_hd__clkbuf_2
X_17696_ _17697_/B _17697_/C _17697_/A vssd1 vssd1 vccd1 vccd1 _17699_/A sky130_fd_sc_hd__a21o_1
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13173__C _13519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19435_ _19418_/A _19418_/C _19418_/B _19419_/X vssd1 vssd1 vccd1 vccd1 _19435_/X
+ sky130_fd_sc_hd__a31o_1
X_16647_ _17039_/C vssd1 vssd1 vccd1 vccd1 _21086_/D sky130_fd_sc_hd__buf_4
X_13859_ _22858_/D vssd1 vssd1 vccd1 vccd1 _13923_/A sky130_fd_sc_hd__inv_2
XFILLER_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19366_ _19200_/B _19195_/Y _19357_/Y vssd1 vssd1 vccd1 vccd1 _19366_/Y sky130_fd_sc_hd__a21oi_1
X_16578_ _16586_/A _16879_/A _11845_/X _17007_/A vssd1 vssd1 vccd1 vccd1 _16578_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18980__B _19771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15529_ _15439_/X _15524_/X _16265_/A _19587_/A _16100_/A vssd1 vssd1 vccd1 vccd1
+ _16253_/B sky130_fd_sc_hd__o2111ai_4
X_18317_ _18319_/A _18313_/Y _18319_/C _22796_/Q vssd1 vssd1 vccd1 vccd1 _18691_/B
+ sky130_fd_sc_hd__o211ai_4
X_19297_ _19043_/X _18023_/A _19265_/X _19065_/X vssd1 vssd1 vccd1 vccd1 _19298_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__15529__D1 _16100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11802__B1 _18665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16781__A _20133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18248_ _18224_/Y _18226_/Y _18230_/Y vssd1 vssd1 vccd1 vccd1 _18772_/B sky130_fd_sc_hd__a21o_1
XANTENNA__21399__A _21399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20734__C _20734_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18179_ _18163_/Y _18174_/A _18177_/X _18178_/Y vssd1 vssd1 vccd1 vccd1 _18181_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__12814__A _15633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20210_ _20210_/A _20210_/B vssd1 vssd1 vccd1 vccd1 _20210_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21190_ _21480_/A vssd1 vssd1 vccd1 vccd1 _21609_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20141_ _12721_/A _12696_/X _12718_/X _16708_/X vssd1 vssd1 vccd1 vccd1 _20142_/C
+ sky130_fd_sc_hd__o22ai_2
XFILLER_143_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20072_ _12522_/A _12522_/B _12767_/A vssd1 vssd1 vccd1 vccd1 _20077_/A sky130_fd_sc_hd__a21o_1
XANTENNA__19316__B _19316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17117__A _20781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20356__A1 _12721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20974_ _21083_/C _21017_/A _21017_/B _20975_/D _20975_/A vssd1 vssd1 vccd1 vccd1
+ _20977_/A sky130_fd_sc_hd__a32o_1
XFILLER_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20478__A _20579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16675__B _22893_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22713_ _22744_/CLK _22713_/D vssd1 vssd1 vccd1 vccd1 _22713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15232__B1 _14552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13380__A _21609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22644_ _22809_/Q input52/X _22652_/S vssd1 vssd1 vccd1 vccd1 _22645_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14195__B _14953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21856__A1 _21220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12597__B2 _15569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22575_ _22575_/A vssd1 vssd1 vccd1 vccd1 _22778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21526_ _21507_/Y _21512_/Y _21464_/X _21465_/Y vssd1 vssd1 vccd1 vccd1 _21529_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_108_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21457_ _21460_/B _21460_/C _21453_/X _21456_/X vssd1 vssd1 vccd1 vccd1 _21666_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_135_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12190_ _12182_/C _12182_/D _12189_/Y vssd1 vssd1 vccd1 vccd1 _18214_/A sky130_fd_sc_hd__a21o_1
X_20408_ _20408_/A vssd1 vssd1 vccd1 vccd1 _20408_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21084__A2 _21083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21388_ _21388_/A vssd1 vssd1 vccd1 vccd1 _21393_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20339_ _20339_/A _20460_/A vssd1 vssd1 vccd1 vccd1 _20339_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__12162__C _19490_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22033__A1 _21683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput88 _14386_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput99 _14415_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[25] sky130_fd_sc_hd__buf_2
XANTENNA__18130__B _19587_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14900_ _14901_/A _14930_/A _14901_/C vssd1 vssd1 vccd1 vccd1 _14904_/B sky130_fd_sc_hd__a21o_1
XFILLER_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22009_ _22013_/A _22013_/B vssd1 vssd1 vccd1 vccd1 _22024_/B sky130_fd_sc_hd__nand2_1
X_15880_ _16209_/A _16403_/A _16402_/B _15879_/X vssd1 vssd1 vccd1 vccd1 _15881_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input23_A wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14831_ _15107_/C vssd1 vssd1 vccd1 vccd1 _15186_/D sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_4_0_bq_clk_i clkbuf_3_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12809__C1 _15352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _17550_/A _17550_/B vssd1 vssd1 vccd1 vccd1 _17550_/Y sky130_fd_sc_hd__nor2_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14762_ _14762_/A _14929_/B vssd1 vssd1 vccd1 vccd1 _22675_/D sky130_fd_sc_hd__xnor2_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ _11974_/A _18338_/C _11974_/C vssd1 vssd1 vccd1 vccd1 _11974_/Y sky130_fd_sc_hd__nand3_2
XFILLER_45_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20388__A _20388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16501_ _16496_/X _16498_/Y _16499_/X _16500_/X vssd1 vssd1 vccd1 vccd1 _16501_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__16585__B _16585_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _14165_/B vssd1 vssd1 vccd1 vccd1 _14054_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17481_ _17475_/X _17476_/Y _17479_/Y _17480_/Y vssd1 vssd1 vccd1 vccd1 _17490_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14693_ _14693_/A _14693_/B _14889_/A _14693_/D vssd1 vssd1 vccd1 vccd1 _14693_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19220_ _19213_/Y _19219_/Y _19208_/A vssd1 vssd1 vccd1 vccd1 _19223_/A sky130_fd_sc_hd__o21ai_1
X_16432_ _16432_/A _16439_/A _16439_/B vssd1 vssd1 vccd1 vccd1 _16432_/Y sky130_fd_sc_hd__nand3_2
XFILLER_147_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13644_ _13643_/A _13643_/B _13643_/C vssd1 vssd1 vccd1 vccd1 _13647_/B sky130_fd_sc_hd__a21oi_1
XFILLER_147_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19151_ _19028_/X _19032_/Y _19085_/Y _19086_/Y vssd1 vssd1 vccd1 vccd1 _19237_/B
+ sky130_fd_sc_hd__o22ai_4
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22917__CLK _22922_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16363_ _16360_/X _16431_/B _15660_/A _15652_/X vssd1 vssd1 vccd1 vccd1 _16369_/C
+ sky130_fd_sc_hd__a31o_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13618_/B _13575_/B vssd1 vssd1 vccd1 vccd1 _13627_/C sky130_fd_sc_hd__nand2_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18102_ _18102_/A _18102_/B vssd1 vssd1 vccd1 vccd1 _18896_/C sky130_fd_sc_hd__nand2_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _15314_/A vssd1 vssd1 vccd1 vccd1 _15911_/A sky130_fd_sc_hd__buf_2
XFILLER_184_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19082_ _19106_/C _19106_/D vssd1 vssd1 vccd1 vccd1 _19082_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15526__A1 _12672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ _15306_/C _12540_/C _12515_/A _12970_/A _22824_/Q vssd1 vssd1 vccd1 vccd1
+ _12526_/X sky130_fd_sc_hd__a32o_1
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16294_ _16294_/A vssd1 vssd1 vccd1 vccd1 _16294_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_173_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18033_ _18033_/A _18065_/A vssd1 vssd1 vccd1 vccd1 _18035_/A sky130_fd_sc_hd__or2b_1
XANTENNA__18305__B _18305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _15244_/B _15245_/B vssd1 vssd1 vccd1 vccd1 _15246_/B sky130_fd_sc_hd__and2b_1
XFILLER_145_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12457_ _12457_/A vssd1 vssd1 vccd1 vccd1 _16477_/C sky130_fd_sc_hd__buf_2
XANTENNA__12634__A _22823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16106__A _16106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _22956_/Q _22955_/Q vssd1 vssd1 vccd1 vccd1 _11712_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15176_ _15176_/A _15180_/B _15180_/A vssd1 vssd1 vccd1 vccd1 _15178_/A sky130_fd_sc_hd__or3_1
X_12388_ _16318_/A _12386_/X _12387_/Y vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__o21ai_2
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16487__C1 _15810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14127_ _14126_/Y _14085_/Y _14071_/Y vssd1 vssd1 vccd1 vccd1 _14128_/C sky130_fd_sc_hd__a21o_1
X_11339_ _11713_/B vssd1 vssd1 vccd1 vccd1 _11720_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19984_ _19419_/B _20012_/B _20012_/C _19901_/B _18028_/A vssd1 vssd1 vccd1 vccd1
+ _19985_/D sky130_fd_sc_hd__a32o_1
XFILLER_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18935_ _18935_/A vssd1 vssd1 vccd1 vccd1 _18935_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14058_ _14061_/A _14061_/D _13923_/X _14057_/X vssd1 vssd1 vccd1 vccd1 _14058_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18678__D _18678_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13009_ _13004_/B _12962_/Y _13004_/A _13012_/A _13012_/B vssd1 vssd1 vccd1 vccd1
+ _13009_/Y sky130_fd_sc_hd__o2111ai_1
X_18866_ _17421_/X _17422_/X _11639_/A vssd1 vssd1 vccd1 vccd1 _18866_/Y sky130_fd_sc_hd__a21oi_2
X_17817_ _17817_/A vssd1 vssd1 vccd1 vccd1 _19839_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18797_ _19351_/B _18797_/B _18797_/C vssd1 vssd1 vccd1 vccd1 _18797_/Y sky130_fd_sc_hd__nand3_4
XFILLER_55_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19152__A _19329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22928__D _22928_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17748_ _17833_/A _19901_/A _20917_/B _19844_/D vssd1 vssd1 vccd1 vccd1 _17752_/B
+ sky130_fd_sc_hd__nand4_1
X_17679_ _17669_/X _17679_/B _17679_/C vssd1 vssd1 vccd1 vccd1 _17681_/A sky130_fd_sc_hd__nand3b_1
XFILLER_165_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19418_ _19418_/A _19418_/B _19418_/C vssd1 vssd1 vccd1 vccd1 _19418_/X sky130_fd_sc_hd__and3_1
XFILLER_126_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20690_ _20793_/A _17833_/B _17833_/C _20936_/B _17530_/A vssd1 vssd1 vccd1 vccd1
+ _20690_/X sky130_fd_sc_hd__a32o_1
XANTENNA__17103__C _17103_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19349_ _19374_/A _19374_/B vssd1 vssd1 vccd1 vccd1 _19371_/A sky130_fd_sc_hd__and2_1
XFILLER_176_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20745__B _21017_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17400__A _17400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22360_ _22341_/B _22338_/A _22338_/B _22816_/Q vssd1 vssd1 vccd1 vccd1 _22360_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21311_ _21185_/A _21187_/A _13519_/B _21480_/A vssd1 vssd1 vccd1 vccd1 _21313_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_11_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22291_ _22206_/C _22206_/A _22682_/Q vssd1 vssd1 vccd1 vccd1 _22291_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16016__A _16016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15558__C _15558_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21242_ _13387_/X _13359_/X _13394_/Y vssd1 vssd1 vccd1 vccd1 _21243_/C sky130_fd_sc_hd__a21boi_1
XFILLER_116_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17809__A3 _21017_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21173_ _21173_/A _21448_/B _21173_/C vssd1 vssd1 vccd1 vccd1 _21173_/Y sky130_fd_sc_hd__nand3_1
XFILLER_85_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20124_ _15504_/X _15546_/A _20123_/X _12792_/C vssd1 vssd1 vccd1 vccd1 _20125_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_172_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15150__C1 _15006_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15574__B _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19967__B1 _22924_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20055_ _20055_/A _20055_/B vssd1 vssd1 vccd1 vccd1 _20055_/Y sky130_fd_sc_hd__nor2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater160 _22751_/CLK vssd1 vssd1 vccd1 vccd1 _22772_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater171 _22690_/CLK vssd1 vssd1 vccd1 vccd1 _22728_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20329__A1 _12721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12806__A2 _15637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20329__B2 _20210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19195__A1 _11786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ _20958_/A _20958_/B _22938_/Q vssd1 vssd1 vccd1 vccd1 _20959_/A sky130_fd_sc_hd__a21o_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12719__A _12719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17745__A2 _20675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19212__D _19587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11644_/X _11646_/Y _11648_/Y vssd1 vssd1 vccd1 vccd1 _11690_/Y sky130_fd_sc_hd__o21ai_2
X_20888_ _20888_/A vssd1 vssd1 vccd1 vccd1 _20894_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22627_ _22627_/A vssd1 vssd1 vccd1 vccd1 _22801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17310__A _17310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ _13423_/A vssd1 vssd1 vccd1 vccd1 _21964_/A sky130_fd_sc_hd__buf_2
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22558_ _22771_/Q input45/X _22558_/S vssd1 vssd1 vccd1 vccd1 _22559_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12311_ _12368_/D _12369_/A vssd1 vssd1 vccd1 vccd1 _12409_/A sky130_fd_sc_hd__nand2_1
XANTENNA__20642__A1_N _20631_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21509_ _21509_/A _21509_/B vssd1 vssd1 vccd1 vccd1 _21509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16181__A1 _15918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ _13087_/A _13300_/A _13139_/B _13322_/A vssd1 vssd1 vccd1 vccd1 _13314_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22489_ _22740_/Q input47/X _22497_/S vssd1 vssd1 vccd1 vccd1 _22490_/A sky130_fd_sc_hd__mux2_1
X_15030_ _15088_/A _15030_/B _15030_/C vssd1 vssd1 vccd1 vccd1 _15088_/B sky130_fd_sc_hd__nand3_1
X_12242_ _18236_/B _18272_/B vssd1 vssd1 vccd1 vccd1 _18249_/B sky130_fd_sc_hd__nand2_1
XANTENNA__21767__A _21767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20804__A2 _15919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12173_ _12156_/X _12162_/Y _12172_/Y vssd1 vssd1 vccd1 vccd1 _12173_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16981_ _16981_/A vssd1 vssd1 vccd1 vccd1 _17188_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18720_ _18722_/A _18722_/B vssd1 vssd1 vccd1 vccd1 _18721_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16299__C _20870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15932_ _15932_/A vssd1 vssd1 vccd1 vccd1 _15932_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15863_ _15864_/C _15864_/D _15862_/Y vssd1 vssd1 vccd1 vccd1 _15952_/B sky130_fd_sc_hd__a21o_1
X_18651_ _11598_/X _16275_/A _18657_/A _18659_/B vssd1 vssd1 vccd1 vccd1 _18654_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__18091__D1 _18093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15402__A2_N _15394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17602_ _17516_/Y _17519_/Y _17605_/B vssd1 vssd1 vccd1 vccd1 _17611_/A sky130_fd_sc_hd__o21bai_2
XFILLER_36_228 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14814_ _14815_/C _14815_/B _14815_/A vssd1 vssd1 vccd1 vccd1 _14816_/A sky130_fd_sc_hd__a21o_1
XFILLER_92_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18582_ _18582_/A _18582_/B _18582_/C vssd1 vssd1 vccd1 vccd1 _18774_/D sky130_fd_sc_hd__nand3_4
X_15794_ _15918_/A _15792_/C _15792_/A _15788_/A _15834_/A vssd1 vssd1 vccd1 vccd1
+ _15794_/X sky130_fd_sc_hd__o311a_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _20870_/A _20870_/B _18303_/A _18303_/B vssd1 vssd1 vccd1 vccd1 _17533_/X
+ sky130_fd_sc_hd__and4_1
X_14745_ _14745_/A _14745_/B _14745_/C vssd1 vssd1 vccd1 vccd1 _14747_/B sky130_fd_sc_hd__nand3_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _11502_/X _11503_/X _16912_/A _11938_/Y _11956_/Y vssd1 vssd1 vccd1 vccd1
+ _11957_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_83_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17464_ _17464_/A _17464_/B vssd1 vssd1 vccd1 vccd1 _17464_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15005__A _15006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13207__C1 _13202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_743 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14676_ _14622_/X _14636_/D _14672_/X vssd1 vssd1 vccd1 vccd1 _14676_/X sky130_fd_sc_hd__a21o_1
XFILLER_177_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16944__B1 _12689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11888_ _15912_/C vssd1 vssd1 vccd1 vccd1 _16103_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_32_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19203_ _12064_/A _18814_/A _19211_/A vssd1 vssd1 vccd1 vccd1 _19203_/X sky130_fd_sc_hd__o21a_1
X_16415_ _16198_/Y _16414_/X _15964_/A _15964_/B vssd1 vssd1 vccd1 vccd1 _16419_/A
+ sky130_fd_sc_hd__o211ai_1
X_13627_ _13627_/A _13627_/B _13627_/C vssd1 vssd1 vccd1 vccd1 _13643_/A sky130_fd_sc_hd__nand3_1
XFILLER_189_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17395_ _17252_/Y _17535_/A _17394_/Y vssd1 vssd1 vccd1 vccd1 _17408_/A sky130_fd_sc_hd__o21ai_1
XFILLER_158_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19489__A2 _17526_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18316__A _18691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19134_ _19134_/A _19134_/B vssd1 vssd1 vccd1 vccd1 _19301_/D sky130_fd_sc_hd__nand2_1
XFILLER_158_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16346_ _15617_/A _16323_/D _16580_/A vssd1 vssd1 vccd1 vccd1 _20357_/C sky130_fd_sc_hd__a21o_1
X_13558_ _13558_/A _13558_/B _13558_/C vssd1 vssd1 vccd1 vccd1 _13612_/A sky130_fd_sc_hd__nand3_1
XFILLER_173_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18161__A2 _12168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19065_ _19065_/A vssd1 vssd1 vccd1 vccd1 _19065_/X sky130_fd_sc_hd__clkbuf_2
X_12509_ _12509_/A vssd1 vssd1 vccd1 vccd1 _12510_/B sky130_fd_sc_hd__clkbuf_2
X_16277_ _16179_/A _17434_/A _16276_/X _16177_/A vssd1 vssd1 vccd1 vccd1 _16277_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__16172__A1 _16124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13489_ _13492_/A _13492_/B vssd1 vssd1 vccd1 vccd1 _13554_/A sky130_fd_sc_hd__xor2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18016_ _18014_/Y _18016_/B vssd1 vssd1 vccd1 vccd1 _18017_/A sky130_fd_sc_hd__and2b_1
XFILLER_173_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15228_ _15197_/X _15210_/X _15227_/X vssd1 vssd1 vccd1 vccd1 _15230_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__21677__A _21677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12733__A1 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17657__D1 _17816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15159_ _15156_/Y _15157_/X _15119_/B _15120_/C vssd1 vssd1 vccd1 vccd1 _15160_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19967_ _19977_/A _19977_/B _22924_/Q vssd1 vssd1 vccd1 vccd1 _19974_/B sky130_fd_sc_hd__a21o_1
XFILLER_45_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18918_ _18713_/A _18713_/B _18836_/A _18725_/A vssd1 vssd1 vccd1 vccd1 _18918_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19898_ _19899_/A _19899_/B _19937_/A _19899_/D vssd1 vssd1 vccd1 vccd1 _19905_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16002__C _16011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18849_ _19504_/A _18850_/A _18849_/C _18849_/D vssd1 vssd1 vccd1 vccd1 _18861_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_68_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16937__C _17128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21860_ _21858_/Y _21859_/X _21857_/A vssd1 vssd1 vccd1 vccd1 _21986_/B sky130_fd_sc_hd__o21bai_2
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19177__A1 _17427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20811_ _20810_/A _20810_/B _20810_/C vssd1 vssd1 vccd1 vccd1 _20812_/D sky130_fd_sc_hd__a21o_1
XANTENNA__17114__B _17311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21791_ _21789_/B _21778_/D _21790_/Y vssd1 vssd1 vccd1 vccd1 _21791_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11443__A _15415_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19610__A _19610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20742_ _20738_/X _20739_/Y _20740_/Y _20741_/Y vssd1 vssd1 vccd1 vccd1 _20748_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12258__B _22909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13749__B1 _13748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_478 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20673_ _15617_/X _12827_/X _20853_/A _17386_/B vssd1 vssd1 vccd1 vccd1 _20782_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22412_ _22412_/A vssd1 vssd1 vccd1 vccd1 _22706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11775__A2 _12165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22343_ _22684_/Q _22289_/B _22324_/B _22342_/Y vssd1 vssd1 vccd1 vccd1 _22343_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_148_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_954 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_998 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22274_ _22301_/A _22301_/B vssd1 vssd1 vccd1 vccd1 _22277_/A sky130_fd_sc_hd__xnor2_1
XFILLER_191_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15910__B2 _15933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21225_ _21216_/A _21216_/B _21183_/X _21212_/Y vssd1 vssd1 vccd1 vccd1 _21227_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16466__A2 _15903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18860__B1 _19313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21156_ _21150_/Y _21151_/X _21154_/B _21155_/X vssd1 vssd1 vccd1 vccd1 _21162_/A
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__18896__A _19329_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20107_ _20107_/A _20107_/B _20107_/C vssd1 vssd1 vccd1 vccd1 _20119_/B sky130_fd_sc_hd__nand3_4
XFILLER_59_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21087_ _21087_/A _21087_/B vssd1 vssd1 vccd1 vccd1 _21088_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20038_ _20018_/A _20018_/B _20016_/A _20037_/X vssd1 vssd1 vccd1 vccd1 _20041_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18612__B1 _19197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19504__B _19504_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12860_ _20120_/A vssd1 vssd1 vccd1 vccd1 _12860_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20970__A1 _17928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _12035_/A _12035_/B _12036_/A vssd1 vssd1 vccd1 vccd1 _11811_/Y sky130_fd_sc_hd__nand3_1
XFILLER_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12788_/B _12788_/C _20241_/A _12929_/A vssd1 vssd1 vccd1 vccd1 _12792_/D
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21989_ _22167_/A _21341_/X _21988_/X vssd1 vssd1 vccd1 vccd1 _21989_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14530_/A _14530_/B vssd1 vssd1 vccd1 vccd1 _14561_/D sky130_fd_sc_hd__nor2_1
X_11742_ _11324_/X _11675_/B _14438_/A _11438_/B vssd1 vssd1 vccd1 vccd1 _11904_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14461_ _14468_/A _14468_/B vssd1 vssd1 vccd1 vccd1 _14461_/Y sky130_fd_sc_hd__nor2_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11673_ _11664_/D _11666_/X _11672_/X _18288_/A _18666_/B vssd1 vssd1 vccd1 vccd1
+ _11673_/X sky130_fd_sc_hd__a32o_2
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17678__C _17678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16200_ _16414_/A _16414_/B _16200_/C _16414_/C vssd1 vssd1 vccd1 vccd1 _16201_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__20385__B _20398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13412_ _21442_/A vssd1 vssd1 vccd1 vccd1 _21268_/A sky130_fd_sc_hd__inv_2
XFILLER_186_269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17180_ _17180_/A _17180_/B _17180_/C vssd1 vssd1 vccd1 vccd1 _17180_/X sky130_fd_sc_hd__and3_1
XANTENNA__22475__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14392_ _22802_/Q _14381_/X _14382_/X _14391_/X _22770_/Q vssd1 vssd1 vccd1 vccd1
+ _14392_/X sky130_fd_sc_hd__a32o_1
XANTENNA__12558__A4 _12672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_995 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18143__A2 _12167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _16131_/A _16131_/B vssd1 vssd1 vccd1 vccd1 _16145_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13343_ _13343_/A vssd1 vssd1 vccd1 vccd1 _13343_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19893__C _22921_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16062_ _16062_/A vssd1 vssd1 vccd1 vccd1 _16586_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_170_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13274_ _13517_/A _13421_/A _13517_/C vssd1 vssd1 vccd1 vccd1 _13274_/Y sky130_fd_sc_hd__nand3_1
XFILLER_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15013_ _15013_/A _15013_/B vssd1 vssd1 vccd1 vccd1 _15015_/B sky130_fd_sc_hd__nand2_1
XFILLER_182_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12225_ _12225_/A vssd1 vssd1 vccd1 vccd1 _18228_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19821_ _19880_/A _19880_/B _19761_/D _19680_/A _19820_/Y vssd1 vssd1 vccd1 vccd1
+ _19822_/C sky130_fd_sc_hd__a311o_1
XFILLER_97_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18851__B1 _18330_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ _12156_/A vssd1 vssd1 vccd1 vccd1 _12156_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19752_ _19680_/A _19761_/D _19751_/Y _19760_/A _19760_/B vssd1 vssd1 vccd1 vccd1
+ _19752_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_150_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16964_ _16964_/A vssd1 vssd1 vccd1 vccd1 _19504_/B sky130_fd_sc_hd__clkbuf_4
X_12087_ _12087_/A _12087_/B _18239_/B vssd1 vssd1 vccd1 vccd1 _12251_/A sky130_fd_sc_hd__nand3_2
XANTENNA__12350__C _20341_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18703_ _18715_/A vssd1 vssd1 vccd1 vccd1 _18722_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15915_ _15915_/A _15915_/B _15915_/C vssd1 vssd1 vccd1 vccd1 _15915_/Y sky130_fd_sc_hd__nand3_1
X_19683_ _19813_/A _19813_/B _19666_/X vssd1 vssd1 vccd1 vccd1 _19683_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16895_ _16895_/A _16895_/B vssd1 vssd1 vccd1 vccd1 _16895_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18634_ _18619_/Y _18835_/A _18633_/Y vssd1 vssd1 vccd1 vccd1 _18634_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _15864_/A _15709_/Y _15734_/X vssd1 vssd1 vccd1 vccd1 _15846_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18565_ _18565_/A _18565_/B vssd1 vssd1 vccd1 vccd1 _18568_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ _11504_/X _11505_/X _11506_/A _15893_/C vssd1 vssd1 vccd1 vccd1 _15779_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12359__A _22821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12989_ _12989_/A _12989_/B _12989_/C vssd1 vssd1 vccd1 vccd1 _12990_/D sky130_fd_sc_hd__nand3_1
XANTENNA__17709__A2 _17227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17516_ _17603_/D _17229_/Y _17515_/X vssd1 vssd1 vccd1 vccd1 _17516_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_33_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14728_ _14727_/B _14727_/C _14624_/A _13905_/Y vssd1 vssd1 vccd1 vccd1 _14728_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_75_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18496_ _19329_/B vssd1 vssd1 vccd1 vccd1 _19694_/D sky130_fd_sc_hd__buf_4
XFILLER_36_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17447_ _19012_/D vssd1 vssd1 vccd1 vccd1 _19619_/D sky130_fd_sc_hd__clkbuf_4
X_14659_ _14758_/A _14758_/B vssd1 vssd1 vccd1 vccd1 _14660_/B sky130_fd_sc_hd__and2_1
XFILLER_178_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15389__B _15389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17378_ _17298_/A _17298_/C _17377_/Y vssd1 vssd1 vccd1 vccd1 _17416_/A sky130_fd_sc_hd__a21oi_1
XFILLER_186_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19117_ _19117_/A _19117_/B _19117_/C vssd1 vssd1 vccd1 vccd1 _19117_/X sky130_fd_sc_hd__and3_2
XFILLER_174_943 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16329_ _16435_/B _16579_/A _22701_/Q vssd1 vssd1 vccd1 vccd1 _20357_/A sky130_fd_sc_hd__o21bai_2
XFILLER_173_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14156__B1 _14147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19048_ _19194_/D _19490_/A _19199_/A _19490_/B vssd1 vssd1 vccd1 vccd1 _19048_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_118_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16448__A2 _11702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21010_ _12671_/X _21048_/B _21048_/C _20514_/X _21082_/C vssd1 vssd1 vccd1 vccd1
+ _21010_/X sky130_fd_sc_hd__o32a_1
XFILLER_88_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21441__A2 _21415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18842__B1 _22798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22961_ _22964_/CLK _22961_/D vssd1 vssd1 vccd1 vccd1 _22961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21912_ _22008_/A _21909_/B _22007_/B vssd1 vssd1 vccd1 vccd1 _21912_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11693__A1 _11561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22892_ _22952_/CLK _22892_/D vssd1 vssd1 vccd1 vccd1 _22892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21843_ _21841_/Y _21733_/A _21842_/X vssd1 vssd1 vccd1 vccd1 _21897_/A sky130_fd_sc_hd__a21oi_1
XFILLER_55_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16964__A _16964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19340__A _19340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21774_ _21736_/Y _21737_/Y _21773_/Y vssd1 vssd1 vccd1 vccd1 _21781_/A sky130_fd_sc_hd__o21ai_1
X_20725_ _20806_/B _17643_/A _20620_/A _20620_/B _20724_/X vssd1 vssd1 vccd1 vccd1
+ _20728_/C sky130_fd_sc_hd__a221oi_4
XANTENNA__15408__A_N _15397_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15299__B _16256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20656_ _20656_/A _20656_/B _20656_/C vssd1 vssd1 vccd1 vccd1 _20660_/A sky130_fd_sc_hd__nand3_4
XFILLER_177_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20587_ _20587_/A _20587_/B vssd1 vssd1 vccd1 vccd1 _20587_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16687__A2 _16670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22326_ _22325_/A _22325_/B _22325_/C vssd1 vssd1 vccd1 vccd1 _22327_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__17884__B2 _20975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22851__D _22863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22257_ _22142_/B _22164_/A _22255_/X _22256_/Y vssd1 vssd1 vccd1 vccd1 _22258_/C
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__15746__C _19772_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _12010_/A vssd1 vssd1 vccd1 vccd1 _19350_/A sky130_fd_sc_hd__clkbuf_4
X_21208_ _21192_/A _21195_/Y _13591_/A _21197_/Y _21615_/A vssd1 vssd1 vccd1 vccd1
+ _21210_/B sky130_fd_sc_hd__o2111ai_1
X_22188_ _22188_/A _22188_/B vssd1 vssd1 vccd1 vccd1 _22231_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21139_ _21066_/X _21137_/Y _21138_/X _21135_/Y _21118_/A vssd1 vssd1 vccd1 vccd1
+ _21141_/B sky130_fd_sc_hd__o311a_1
XFILLER_120_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13961_ _13833_/X _13736_/B _14112_/A vssd1 vssd1 vccd1 vccd1 _14073_/A sky130_fd_sc_hd__o21ai_2
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21196__A1 _21185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15700_ _15707_/B _15700_/B _15700_/C vssd1 vssd1 vccd1 vccd1 _15740_/C sky130_fd_sc_hd__nand3_1
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12912_ _12912_/A _20793_/B _16067_/B _12958_/B vssd1 vssd1 vccd1 vccd1 _12958_/C
+ sky130_fd_sc_hd__nand4_2
X_16680_ _16683_/B _16683_/C _16426_/X vssd1 vssd1 vccd1 vccd1 _16680_/X sky130_fd_sc_hd__a21o_1
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15481__C _22662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13892_ _13892_/A _13892_/B vssd1 vssd1 vccd1 vccd1 _13907_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15631_ _15631_/A _15631_/B _15631_/C vssd1 vssd1 vccd1 vccd1 _15631_/X sky130_fd_sc_hd__and3_4
X_12843_ _20120_/A _12859_/A _12859_/B vssd1 vssd1 vccd1 vccd1 _12843_/X sky130_fd_sc_hd__and3_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15562_ _11704_/X _11705_/X _16779_/A _16778_/A _11707_/A vssd1 vssd1 vccd1 vccd1
+ _15568_/B sky130_fd_sc_hd__o221a_1
X_18350_ _11361_/A _18135_/A _18343_/X _18337_/X _18340_/Y vssd1 vssd1 vccd1 vccd1
+ _18351_/C sky130_fd_sc_hd__o221ai_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12774_/A vssd1 vssd1 vccd1 vccd1 _12774_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17301_/A _17301_/B _17301_/C vssd1 vssd1 vccd1 vccd1 _17334_/A sky130_fd_sc_hd__nand3_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14134_/Y _13968_/Y _14002_/C _14002_/A vssd1 vssd1 vccd1 vccd1 _14515_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11725_ _11718_/A _12210_/A _15481_/A vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__a21o_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20827__C _20827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15493_ _19197_/C _19197_/D _16489_/A vssd1 vssd1 vccd1 vccd1 _15567_/B sky130_fd_sc_hd__and3_1
X_18281_ _11859_/X _11861_/X _18453_/C _19358_/A _19358_/B vssd1 vssd1 vccd1 vccd1
+ _18281_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_159_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12907__A _16129_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17232_ _17200_/A _17331_/A _17231_/Y vssd1 vssd1 vccd1 vccd1 _17485_/A sky130_fd_sc_hd__a21o_1
XFILLER_175_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14444_ _16130_/B vssd1 vssd1 vccd1 vccd1 _16400_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11656_ _11668_/A _16242_/A _15435_/D vssd1 vssd1 vccd1 vccd1 _11656_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_174_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11739__A2 _11626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12936__A1 _12988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17163_ _16760_/X _17138_/X _16949_/Y vssd1 vssd1 vccd1 vccd1 _17163_/X sky130_fd_sc_hd__a21o_1
X_14375_ _22798_/Q _14354_/X _14355_/X _14361_/X _22766_/Q vssd1 vssd1 vccd1 vccd1
+ _14375_/X sky130_fd_sc_hd__a32o_1
XFILLER_31_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16127__B2 _16015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ _11587_/A _11790_/C _11587_/C vssd1 vssd1 vccd1 vccd1 _11793_/A sky130_fd_sc_hd__nand3_2
XFILLER_31_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16114_ _16169_/C vssd1 vssd1 vccd1 vccd1 _16174_/A sky130_fd_sc_hd__inv_2
XANTENNA__14138__B1 _14491_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13326_ _22844_/Q vssd1 vssd1 vccd1 vccd1 _13326_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17094_ _17088_/X _17094_/B _17094_/C vssd1 vssd1 vccd1 vccd1 _17341_/C sky130_fd_sc_hd__nand3b_4
XFILLER_143_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16045_ _16045_/A _16045_/B _16045_/C vssd1 vssd1 vccd1 vccd1 _16047_/A sky130_fd_sc_hd__nand3_4
XANTENNA_clkbuf_3_3_0_bq_clk_i_A clkbuf_3_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ _13257_/A _13257_/B vssd1 vssd1 vccd1 vccd1 _13662_/C sky130_fd_sc_hd__nand2_2
XFILLER_143_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19616__A2 _19624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ _16226_/C _12208_/B vssd1 vssd1 vccd1 vccd1 _12209_/A sky130_fd_sc_hd__nor2_2
XFILLER_123_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13457__B _21498_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13188_ _13161_/C _13161_/A _13157_/A _13131_/X vssd1 vssd1 vccd1 vccd1 _13450_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19804_ _19804_/A _19804_/B vssd1 vssd1 vccd1 vccd1 _19804_/X sky130_fd_sc_hd__and2_1
XFILLER_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15953__A _17525_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _12139_/A vssd1 vssd1 vccd1 vccd1 _18162_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17996_ _17996_/A _17996_/B vssd1 vssd1 vccd1 vccd1 _18020_/D sky130_fd_sc_hd__xnor2_2
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13113__A1 _13112_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19735_ _19735_/A _19735_/B _19735_/C vssd1 vssd1 vccd1 vccd1 _19736_/B sky130_fd_sc_hd__nand3_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16947_ _16947_/A _17139_/A _17140_/A vssd1 vssd1 vccd1 vccd1 _17145_/A sky130_fd_sc_hd__nand3_1
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19666_ _19814_/A _19814_/B vssd1 vssd1 vccd1 vccd1 _19666_/X sky130_fd_sc_hd__or2_1
XFILLER_65_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16878_ _20936_/C vssd1 vssd1 vccd1 vccd1 _17840_/A sky130_fd_sc_hd__clkbuf_2
X_18617_ _17635_/A _12116_/X _18613_/B _18451_/B vssd1 vssd1 vccd1 vccd1 _18618_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15829_ _15829_/A vssd1 vssd1 vccd1 vccd1 _15915_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19597_ _19497_/B _19494_/Y _19500_/X _19359_/X vssd1 vssd1 vccd1 vccd1 _19684_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19160__A _19160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18548_ _18548_/A _18548_/B vssd1 vssd1 vccd1 vccd1 _18557_/A sky130_fd_sc_hd__nand2_1
XFILLER_166_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18479_ _18565_/B vssd1 vssd1 vccd1 vccd1 _18765_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20510_ _20249_/B _17401_/A _17401_/B _20503_/Y _20505_/Y vssd1 vssd1 vccd1 vccd1
+ _20511_/D sky130_fd_sc_hd__a32o_1
XANTENNA__22439__A1 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20456__D _20576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21490_ _21490_/A _21490_/B vssd1 vssd1 vccd1 vccd1 _21490_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12927__A1 _12772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20441_ _20441_/A _20441_/B vssd1 vssd1 vccd1 vccd1 _22912_/D sky130_fd_sc_hd__xor2_4
XFILLER_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20372_ _20349_/A _20366_/C _20371_/Y vssd1 vssd1 vccd1 vccd1 _20375_/A sky130_fd_sc_hd__a21o_1
XFILLER_162_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22111_ _22040_/Y _22108_/Y _22179_/A _22105_/X vssd1 vssd1 vccd1 vccd1 _22111_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_162_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12155__A2 _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1071 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22042_ _22042_/A _22105_/A vssd1 vssd1 vccd1 vccd1 _22042_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__22611__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1052 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1085 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19335__A _19587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16841__A2 _16842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14479__A _14721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22944_ _22944_/CLK _22944_/D vssd1 vssd1 vccd1 vccd1 _22944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22875_ _22916_/CLK _22875_/D vssd1 vssd1 vccd1 vccd1 _22875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14604__A1 _15050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20928__B _20928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21826_ _21825_/A _21825_/B _22677_/Q vssd1 vssd1 vccd1 vccd1 _21831_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21757_ _21757_/A _22058_/A _21877_/A _21757_/D vssd1 vssd1 vccd1 vccd1 _21758_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12727__A _12727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ _18512_/A vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__buf_4
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20708_ _20110_/B _20689_/Y _20690_/X _20796_/B _20797_/A vssd1 vssd1 vccd1 vccd1
+ _20709_/C sky130_fd_sc_hd__o2111ai_2
X_12490_ _12358_/X _12432_/Y _12455_/Y _12480_/X _12489_/Y vssd1 vssd1 vccd1 vccd1
+ _12510_/A sky130_fd_sc_hd__o221ai_4
XFILLER_180_1078 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21688_ _21688_/A _21688_/B _21688_/C vssd1 vssd1 vccd1 vccd1 _21837_/A sky130_fd_sc_hd__nand3_2
XFILLER_196_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22950__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11441_ _15714_/B vssd1 vssd1 vccd1 vccd1 _16711_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__16109__A1 _12500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20639_ _20449_/B _20178_/A _20734_/C _20734_/B vssd1 vssd1 vccd1 vccd1 _20639_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14942__A _14942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14160_ _22870_/Q vssd1 vssd1 vccd1 vccd1 _14494_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_153_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11372_ _11372_/A vssd1 vssd1 vccd1 vccd1 _11911_/A sky130_fd_sc_hd__buf_4
XFILLER_164_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13111_ _22725_/Q _13110_/Y _13234_/C _13057_/C vssd1 vssd1 vccd1 vccd1 _13344_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_152_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19059__B1 _18665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22309_ _22309_/A _22309_/B vssd1 vssd1 vccd1 vccd1 _22310_/B sky130_fd_sc_hd__nand2_1
XFILLER_166_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14091_ _14169_/A _14169_/B _14169_/C _14090_/Y vssd1 vssd1 vccd1 vccd1 _14091_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_124_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15476__C _20133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17609__A1 _17226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A wb_dat_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ _12882_/A _20183_/A _12757_/A _12757_/B vssd1 vssd1 vccd1 vccd1 _13044_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__22602__A1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12551__C1 _12470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17850_ _17800_/Y _18048_/C _17849_/Y vssd1 vssd1 vccd1 vccd1 _17850_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_182_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21494__B _21494_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16801_ _16972_/A _16971_/A _16798_/X _16800_/X vssd1 vssd1 vccd1 vccd1 _16908_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17781_ _17781_/A _17781_/B _17781_/C vssd1 vssd1 vccd1 vccd1 _17781_/Y sky130_fd_sc_hd__nand3_1
XFILLER_8_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14993_ _14792_/A _14792_/B _14942_/A _14942_/C vssd1 vssd1 vccd1 vccd1 _14996_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_59_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19520_ _19510_/Y _19513_/Y _19514_/X _19532_/A vssd1 vssd1 vccd1 vccd1 _19523_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16732_ _16732_/A _16732_/B vssd1 vssd1 vccd1 vccd1 _16732_/Y sky130_fd_sc_hd__nand2_4
XFILLER_47_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13944_ _14613_/A _14181_/C _14181_/A _13935_/X _13931_/X vssd1 vssd1 vccd1 vccd1
+ _13947_/B sky130_fd_sc_hd__a32o_1
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16100__C _16106_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19451_ _19290_/A _19290_/B _19288_/Y _19289_/A vssd1 vssd1 vccd1 vccd1 _19452_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11525__B _18482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16663_ _17064_/C _16660_/Y _22893_/Q vssd1 vssd1 vccd1 vccd1 _16663_/Y sky130_fd_sc_hd__a21oi_1
X_13875_ _13875_/A vssd1 vssd1 vccd1 vccd1 _14722_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__20392__A2 _12501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18402_ _18402_/A _18402_/B vssd1 vssd1 vccd1 vccd1 _18442_/C sky130_fd_sc_hd__nor2_2
XFILLER_179_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15614_ _20101_/B vssd1 vssd1 vccd1 vccd1 _20098_/D sky130_fd_sc_hd__clkbuf_4
X_12826_ _15608_/C _16322_/A vssd1 vssd1 vccd1 vccd1 _15370_/B sky130_fd_sc_hd__nand2_2
X_19382_ _19457_/A _19389_/B _19389_/C vssd1 vssd1 vccd1 vccd1 _19458_/B sky130_fd_sc_hd__nand3_1
X_16594_ _16594_/A _16594_/B _16594_/C vssd1 vssd1 vccd1 vccd1 _16873_/A sky130_fd_sc_hd__nand3_2
XFILLER_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18333_ _18492_/A vssd1 vssd1 vccd1 vccd1 _18333_/X sky130_fd_sc_hd__buf_2
X_15545_ _18203_/C vssd1 vssd1 vccd1 vccd1 _15545_/X sky130_fd_sc_hd__buf_4
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12757_ _12757_/A _12757_/B vssd1 vssd1 vccd1 vccd1 _12891_/A sky130_fd_sc_hd__nor2_1
XFILLER_91_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12637__A _16486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11541__A _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ _11502_/A _11503_/A _11704_/X _11705_/X _15458_/A vssd1 vssd1 vccd1 vccd1
+ _11708_/Y sky130_fd_sc_hd__o221ai_4
X_18264_ _18261_/X _18251_/Y _18088_/Y _18263_/X vssd1 vssd1 vccd1 vccd1 _18268_/A
+ sky130_fd_sc_hd__a211oi_2
X_15476_ _15476_/A _20133_/A _20133_/B vssd1 vssd1 vccd1 vccd1 _15477_/B sky130_fd_sc_hd__and3_1
X_12688_ _15299_/C _15299_/D _20355_/D vssd1 vssd1 vccd1 vccd1 _12689_/C sky130_fd_sc_hd__and3_1
X_17215_ _17215_/A _17215_/B _17215_/C _17215_/D vssd1 vssd1 vccd1 vccd1 _17215_/Y
+ sky130_fd_sc_hd__nand4_4
X_14427_ _22815_/Q _14354_/A _14355_/A _14361_/A _22783_/Q vssd1 vssd1 vccd1 vccd1
+ _14427_/X sky130_fd_sc_hd__a32o_1
X_11639_ _11639_/A vssd1 vssd1 vccd1 vccd1 _11639_/X sky130_fd_sc_hd__buf_2
X_18195_ _11634_/A _15839_/A _18194_/Y vssd1 vssd1 vccd1 vccd1 _18195_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_144_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17146_ _16060_/A _17400_/A _17138_/X _17142_/X _17145_/Y vssd1 vssd1 vccd1 vccd1
+ _17146_/Y sky130_fd_sc_hd__o221ai_4
X_14358_ _22699_/Q vssd1 vssd1 vccd1 vccd1 _16322_/B sky130_fd_sc_hd__buf_2
XFILLER_143_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13309_ _21207_/A _13309_/B _21495_/C _13521_/B vssd1 vssd1 vccd1 vccd1 _13309_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_171_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17077_ _17077_/A _17077_/B vssd1 vssd1 vccd1 vccd1 _17078_/B sky130_fd_sc_hd__nor2_1
XFILLER_170_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12372__A _22817_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14289_ _14289_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14289_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16028_ _15967_/X _15971_/Y _16021_/Y vssd1 vssd1 vccd1 vccd1 _16028_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13187__B _22845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16779__A _16779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17979_ _19899_/B vssd1 vssd1 vccd1 vccd1 _18023_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18025__A1 _21048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19718_ _19864_/B _19799_/B _19788_/B _19719_/B vssd1 vssd1 vccd1 vccd1 _19725_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18025__B2 _21081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22823__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11648__B2 _11641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12845__B1 _12721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20990_ _20990_/A _20990_/B vssd1 vssd1 vccd1 vccd1 _21006_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16036__B1 _15942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19773__A1 _15840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19773__B2 _17636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19649_ _19643_/Y _19649_/B _19649_/C vssd1 vssd1 vccd1 vccd1 _19650_/D sky130_fd_sc_hd__nand3b_1
XFILLER_168_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22666__D _22666_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22660_ _22662_/A _22660_/B vssd1 vssd1 vccd1 vccd1 _22661_/A sky130_fd_sc_hd__and2_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21611_ _21607_/X _21613_/A _21614_/A vssd1 vssd1 vccd1 vccd1 _21766_/A sky130_fd_sc_hd__o21ai_1
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17122__B _17122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22591_ _11395_/A input46/X _22597_/S vssd1 vssd1 vccd1 vccd1 _22592_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11451__A _18303_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17000__A2 _16712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14465__C _14564_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21542_ _21535_/X _21536_/Y _21540_/Y _21541_/X vssd1 vssd1 vccd1 vccd1 _21546_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_193_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_6_0_bq_clk_i clkbuf_4_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _22915_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_119_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21579__B _21580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21473_ _21473_/A _21583_/D vssd1 vssd1 vccd1 vccd1 _21473_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15562__A2 _11705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20424_ _20549_/D vssd1 vssd1 vccd1 vccd1 _20424_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15577__B _17672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18497__D1 _19694_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16511__A1 _15997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20355_ _20355_/A _20582_/C _20582_/A _20355_/D vssd1 vssd1 vccd1 vccd1 _20370_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20286_ _20286_/A _20286_/B _20286_/C vssd1 vssd1 vccd1 vccd1 _20298_/A sky130_fd_sc_hd__nand3_2
XFILLER_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22025_ _21908_/X _21911_/X _22024_/Y vssd1 vssd1 vccd1 vccd1 _22025_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_103_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20071__A1 _13041_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11990_ _22793_/Q vssd1 vssd1 vccd1 vccd1 _12107_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__12836__B1 _16708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22927_ _22949_/CLK _22927_/D vssd1 vssd1 vccd1 vccd1 _22927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16578__B2 _17007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13660_ _13660_/A _13665_/D vssd1 vssd1 vccd1 vccd1 _13660_/X sky130_fd_sc_hd__and2_1
X_22858_ _22943_/CLK _22858_/D vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15250__A1 _15230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _16515_/A _12938_/A _12973_/A _20576_/B vssd1 vssd1 vccd1 vccd1 _12611_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21809_ _21809_/A _21809_/B vssd1 vssd1 vccd1 vccd1 _21814_/D sky130_fd_sc_hd__nand2_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13591_/A vssd1 vssd1 vccd1 vccd1 _21874_/A sky130_fd_sc_hd__buf_2
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17527__B1 _17443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22789_ _22789_/CLK _22789_/D vssd1 vssd1 vccd1 vccd1 _22789_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__20126__A2 _15355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _20130_/B vssd1 vssd1 vccd1 vccd1 _16781_/B sky130_fd_sc_hd__clkbuf_4
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12542_ _20210_/A _12988_/C _12479_/A vssd1 vssd1 vccd1 vccd1 _12543_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__17967__B _22904_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17542__A3 _19768_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15261_ _15230_/A _15247_/X _15205_/B _15249_/Y vssd1 vssd1 vccd1 vccd1 _15262_/B
+ sky130_fd_sc_hd__o211ai_1
X_12473_ _12518_/A vssd1 vssd1 vccd1 vccd1 _12528_/A sky130_fd_sc_hd__buf_2
XFILLER_185_879 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19819__A2 _18246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17000_ _16710_/Y _16712_/X _16711_/Y vssd1 vssd1 vccd1 vccd1 _17001_/C sky130_fd_sc_hd__a21boi_1
X_14212_ _14917_/C _14779_/A _15004_/D _14212_/D vssd1 vssd1 vccd1 vccd1 _14265_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11424_ _12154_/C vssd1 vssd1 vccd1 vccd1 _18682_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_6_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15192_ _15154_/X _15156_/Y _15189_/A _15190_/X vssd1 vssd1 vccd1 vccd1 _15216_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_137_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14143_ _14576_/A vssd1 vssd1 vccd1 vccd1 _14143_/X sky130_fd_sc_hd__buf_2
X_11355_ _22968_/Q vssd1 vssd1 vccd1 vccd1 _11434_/A sky130_fd_sc_hd__inv_2
XFILLER_4_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15305__A2 _15309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16502__B2 _16501_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12119__A2 _16014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18951_ _18955_/A _18951_/B _18951_/C vssd1 vssd1 vccd1 vccd1 _18958_/B sky130_fd_sc_hd__nand3b_2
X_14074_ _14074_/A vssd1 vssd1 vccd1 vccd1 _14576_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_180_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ _11936_/A vssd1 vssd1 vccd1 vccd1 _18107_/A sky130_fd_sc_hd__buf_2
XFILLER_180_595 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17902_ _18020_/A _18020_/B vssd1 vssd1 vccd1 vccd1 _17949_/B sky130_fd_sc_hd__xnor2_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13025_ _12982_/A _12982_/B _13024_/X _13022_/X _20284_/A vssd1 vssd1 vccd1 vccd1
+ _13028_/B sky130_fd_sc_hd__a32o_1
X_18882_ _12009_/X _19313_/A _18493_/A _18875_/Y _18881_/X vssd1 vssd1 vccd1 vccd1
+ _18883_/C sky130_fd_sc_hd__o221ai_1
XANTENNA__22846__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17833_ _17833_/A _17833_/B _17833_/C vssd1 vssd1 vccd1 vccd1 _17833_/X sky130_fd_sc_hd__and3_1
XANTENNA__17463__C1 _21011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11536__A _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19204__B1 _17393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17764_ _17765_/A _17765_/B _17763_/X vssd1 vssd1 vccd1 vccd1 _17768_/B sky130_fd_sc_hd__o21ba_1
XFILLER_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14976_ _14977_/B _15035_/A _14977_/A vssd1 vssd1 vccd1 vccd1 _14980_/A sky130_fd_sc_hd__a21o_1
XFILLER_47_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19503_ _19503_/A _19503_/B _19503_/C vssd1 vssd1 vccd1 vccd1 _19580_/A sky130_fd_sc_hd__nand3_2
XANTENNA__18558__A2 _18407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16715_ _16715_/A vssd1 vssd1 vccd1 vccd1 _20781_/A sky130_fd_sc_hd__buf_2
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16569__A1 _11800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13927_ _13814_/A _13814_/B _14502_/A vssd1 vssd1 vccd1 vccd1 _13927_/X sky130_fd_sc_hd__a21o_1
X_17695_ _17695_/A vssd1 vssd1 vccd1 vccd1 _17697_/A sky130_fd_sc_hd__inv_2
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19434_ _19434_/A _19434_/B vssd1 vssd1 vccd1 vccd1 _19434_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16646_ _16444_/Y _16445_/X _16644_/Y _16645_/X vssd1 vssd1 vccd1 vccd1 _17076_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_35_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _14571_/A _13857_/X _13725_/A vssd1 vssd1 vccd1 vccd1 _13930_/B sky130_fd_sc_hd__o21ai_4
XFILLER_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19365_ _16940_/X _18718_/X _19350_/A _18282_/X vssd1 vssd1 vccd1 vccd1 _19365_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_16_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12809_ _12804_/Y _15409_/A _20346_/C _15352_/A _12808_/Y vssd1 vssd1 vccd1 vccd1
+ _12810_/C sky130_fd_sc_hd__o2111ai_4
X_16577_ _20697_/C vssd1 vssd1 vccd1 vccd1 _17007_/A sky130_fd_sc_hd__buf_2
XANTENNA__19884__B1_N _22922_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13789_ _14212_/D vssd1 vssd1 vccd1 vccd1 _14273_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18980__C _18980_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18316_ _18691_/A vssd1 vssd1 vccd1 vccd1 _19322_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__15529__C1 _19587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15528_ _15528_/A vssd1 vssd1 vccd1 vccd1 _19587_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19296_ _19296_/A _19434_/A vssd1 vssd1 vccd1 vccd1 _19298_/A sky130_fd_sc_hd__nand2_1
XFILLER_187_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16781__B _16781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18247_ _18247_/A vssd1 vssd1 vccd1 vccd1 _19443_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15459_ _11324_/X _11675_/B _15482_/B _11737_/X vssd1 vssd1 vccd1 vccd1 _15810_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_175_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20734__D _20928_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18178_ _18184_/A _18184_/B vssd1 vssd1 vccd1 vccd1 _18178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12814__B _16450_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17129_ _17234_/A _17129_/B _20323_/B vssd1 vssd1 vccd1 vccd1 _17129_/Y sky130_fd_sc_hd__nand3_4
XFILLER_143_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18494__A1 _11541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20140_ _20129_/Y _20131_/Y _20134_/X vssd1 vssd1 vccd1 vccd1 _20143_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__14504__B1 _14503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11869__A1 _11308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20071_ _13041_/Y _20064_/Y _20314_/B _13046_/Y vssd1 vssd1 vccd1 vccd1 _20189_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_170_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1096 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14807__A1 _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20759__A _20759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19332__B _19512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20973_ _20972_/D _21083_/A _21083_/B _21011_/B _20972_/B vssd1 vssd1 vccd1 vccd1
+ _20975_/A sky130_fd_sc_hd__a32o_1
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20478__B _20579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17133__A _17133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22712_ _22744_/CLK _22712_/D vssd1 vssd1 vccd1 vccd1 _22712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16965__D1 _19504_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22643_ _22643_/A vssd1 vssd1 vccd1 vccd1 _22652_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22574_ _22778_/Q input53/X _22580_/S vssd1 vssd1 vccd1 vccd1 _22575_/A sky130_fd_sc_hd__mux2_1
XANTENNA__21856__A2 _21853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21525_ _21539_/A _21539_/B vssd1 vssd1 vccd1 vccd1 _21531_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21456_ _22034_/A _21866_/C _13326_/Y _21455_/X vssd1 vssd1 vccd1 vccd1 _21456_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_181_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20407_ _20427_/A _20427_/B _20407_/C vssd1 vssd1 vccd1 vccd1 _20420_/A sky130_fd_sc_hd__nand3_2
XFILLER_147_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21387_ _21387_/A _21387_/B vssd1 vssd1 vccd1 vccd1 _21387_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__22869__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21084__A3 _21083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20338_ _20341_/A _20341_/B _20338_/C vssd1 vssd1 vccd1 vccd1 _20460_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19507__B _19507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12162__D _19490_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22033__A2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20269_ _20408_/A vssd1 vssd1 vccd1 vccd1 _20269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput89 _14388_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18130__C _18130_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22008_ _22008_/A _22008_/B _22008_/C _22008_/D vssd1 vssd1 vccd1 vccd1 _22013_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14830_ _14963_/C vssd1 vssd1 vccd1 vccd1 _15107_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19737__A1 _19689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A wb_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11973_ _11361_/A _11639_/A _11793_/B _11793_/A vssd1 vssd1 vccd1 vccd1 _11976_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_57_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14761_ _14761_/A _14761_/B vssd1 vssd1 vccd1 vccd1 _14929_/B sky130_fd_sc_hd__xnor2_4
XFILLER_91_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_730 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _16241_/D _15536_/X _16240_/X _12716_/A vssd1 vssd1 vccd1 vccd1 _16500_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13712_ _14212_/D _15114_/C _15115_/C _14273_/C vssd1 vssd1 vccd1 vccd1 _14165_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_72_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17480_ _17479_/A _17479_/B _17469_/A _17469_/B vssd1 vssd1 vccd1 vccd1 _17480_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _14270_/A _15056_/A _14785_/A _14688_/Y _14685_/Y vssd1 vssd1 vccd1 vccd1
+ _14695_/B sky130_fd_sc_hd__a32o_1
XFILLER_72_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16431_ _16431_/A _16431_/B _16431_/C _16444_/A vssd1 vssd1 vccd1 vccd1 _16439_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17978__A _19896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13643_ _13643_/A _13643_/B _13643_/C vssd1 vssd1 vccd1 vccd1 _13647_/C sky130_fd_sc_hd__and3_1
XFILLER_188_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19150_ _19254_/A _19254_/B _19149_/X vssd1 vssd1 vccd1 vccd1 _19150_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__13785__A1 _14079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16362_ _15646_/X _15645_/X _20793_/C _16586_/B _16400_/A vssd1 vssd1 vccd1 vccd1
+ _16431_/B sky130_fd_sc_hd__o2111ai_4
X_13574_ _13401_/A _21848_/B _13618_/A _13573_/A vssd1 vssd1 vccd1 vccd1 _13575_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18101_ _18128_/A _18127_/B vssd1 vssd1 vccd1 vccd1 _18102_/B sky130_fd_sc_hd__nand2_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _15313_/A _15313_/B _15313_/C vssd1 vssd1 vccd1 vccd1 _15386_/A sky130_fd_sc_hd__nand3_1
X_12525_ _12525_/A _12525_/B vssd1 vssd1 vccd1 vccd1 _12970_/A sky130_fd_sc_hd__nand2_2
X_19081_ _19254_/A _19254_/B _19104_/A _19096_/A vssd1 vssd1 vccd1 vccd1 _19106_/D
+ sky130_fd_sc_hd__nand4_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16293_ _16293_/A vssd1 vssd1 vccd1 vccd1 _16293_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18032_ _18030_/C _18030_/Y _18025_/X _18029_/X vssd1 vssd1 vccd1 vccd1 _18065_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18305__C _18305_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15244_ _15245_/B _15244_/B vssd1 vssd1 vccd1 vccd1 _15259_/A sky130_fd_sc_hd__and2b_1
XANTENNA__20554__D _20554_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ _12448_/Y _12449_/Y _12322_/X vssd1 vssd1 vccd1 vccd1 _12456_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_184_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16106__B _16106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11407_ _11727_/C _11407_/B vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18476__A1 _18305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15010__B _15115_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15175_ _15101_/B _15175_/B _15175_/C _15175_/D vssd1 vssd1 vccd1 vccd1 _15180_/A
+ sky130_fd_sc_hd__and4b_1
XANTENNA__19673__B1 _22919_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12387_ _12387_/A _12387_/B vssd1 vssd1 vccd1 vccd1 _12387_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16487__B1 _16964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ _14126_/A _14126_/B _14693_/B vssd1 vssd1 vccd1 vccd1 _14126_/Y sky130_fd_sc_hd__nand3_1
X_11338_ _11334_/X _11423_/A _15539_/A vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__20283__B2 _20429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19983_ _19983_/A _19983_/B _19987_/B _19987_/C vssd1 vssd1 vccd1 vccd1 _19985_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_154_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13168__D _21595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15695__D1 _16100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18934_ _18646_/A _18646_/C _18933_/X vssd1 vssd1 vccd1 vccd1 _18935_/A sky130_fd_sc_hd__a21oi_2
XFILLER_141_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14057_ _14057_/A vssd1 vssd1 vccd1 vccd1 _14057_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13008_ _13007_/B _13007_/C _12749_/A _12749_/B vssd1 vssd1 vccd1 vccd1 _13012_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__21963__A _21963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18865_ _18865_/A _19013_/C _19602_/C vssd1 vssd1 vccd1 vccd1 _18865_/X sky130_fd_sc_hd__and3_1
XANTENNA__13465__B _13465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15383__D _15665_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17816_ _17816_/A _17816_/B _19842_/D _19896_/B vssd1 vssd1 vccd1 vccd1 _17886_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__15961__A _17645_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18796_ _11474_/X _15545_/X _18795_/X _12216_/X vssd1 vssd1 vccd1 vccd1 _18796_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20579__A _20579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17747_ _19774_/D vssd1 vssd1 vccd1 vccd1 _19901_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19152__B _19694_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14959_ _14959_/A _14959_/B _14959_/C vssd1 vssd1 vccd1 vccd1 _14960_/B sky130_fd_sc_hd__nand3_1
XANTENNA__14577__A _14684_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17678_ _17678_/A _17678_/B _17678_/C _17678_/D vssd1 vssd1 vccd1 vccd1 _17679_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19417_ _19306_/X _19203_/X _19411_/X _19555_/A vssd1 vssd1 vccd1 vccd1 _19417_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_51_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16629_ _15653_/Y _16628_/X _15660_/C _16369_/A vssd1 vssd1 vccd1 vccd1 _16630_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_23_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16962__A1 _16179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16501__A1_N _16496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19348_ _19455_/A _19346_/Y _18795_/X _18814_/X vssd1 vssd1 vccd1 vccd1 _19374_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_149_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20745__C _20745_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19279_ _19279_/A _19279_/B vssd1 vssd1 vccd1 vccd1 _19301_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20510__A2 _17401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21310_ _21482_/A vssd1 vssd1 vccd1 vccd1 _21466_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22290_ _22290_/A _22290_/B _22290_/C _22290_/D vssd1 vssd1 vccd1 vccd1 _22290_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_163_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15558__D _20133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21241_ _21231_/A _21247_/C _21240_/A vssd1 vssd1 vccd1 vccd1 _21243_/B sky130_fd_sc_hd__a21o_1
XFILLER_105_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18512__A _18512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21172_ _13337_/C _13329_/X _21216_/A _13346_/X vssd1 vssd1 vccd1 vccd1 _21179_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_116_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20123_ _20123_/A vssd1 vssd1 vccd1 vccd1 _20123_/X sky130_fd_sc_hd__buf_2
XFILLER_77_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17128__A _19694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19046__C _19046_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22969__A input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20054_ _20025_/X _20059_/B _22928_/Q vssd1 vssd1 vccd1 vccd1 _20055_/B sky130_fd_sc_hd__o21a_1
XFILLER_98_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input8_A wb_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16245__A3 _19507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater150 _22804_/CLK vssd1 vssd1 vccd1 vccd1 _22807_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15453__A1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater161 _22771_/CLK vssd1 vssd1 vccd1 vccd1 _22751_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater172 _22725_/CLK vssd1 vssd1 vccd1 vccd1 _22690_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20329__A2 _15718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11904__A _11904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20956_ _20834_/X _20835_/X _20906_/Y _21007_/B vssd1 vssd1 vccd1 vccd1 _20958_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17745__A3 _18305_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__A1 _12018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16953__A1 _12727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _20887_/A _20887_/B _20887_/C vssd1 vssd1 vccd1 vccd1 _20888_/A sky130_fd_sc_hd__or3_1
XFILLER_42_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22626_ _22801_/Q input43/X _22630_/S vssd1 vssd1 vccd1 vccd1 _22627_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22854__D _22866_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14964__B1 _14670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14809__A2_N _14808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22557_ _22557_/A vssd1 vssd1 vccd1 vccd1 _22770_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12735__A _15450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12310_ _12340_/A vssd1 vssd1 vccd1 vccd1 _12401_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21508_ _21508_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21508_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13290_ _13484_/A _13290_/B vssd1 vssd1 vccd1 vccd1 _13392_/A sky130_fd_sc_hd__nand2_1
XFILLER_155_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16181__A2 _20449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22488_ _22499_/A vssd1 vssd1 vccd1 vccd1 _22497_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_166_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12241_ _12241_/A _12241_/B _12241_/C vssd1 vssd1 vccd1 vccd1 _18272_/B sky130_fd_sc_hd__nand3_2
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21439_ _22675_/Q vssd1 vssd1 vccd1 vccd1 _21568_/A sky130_fd_sc_hd__inv_2
XFILLER_182_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12172_ _12170_/X _12171_/X _18716_/A vssd1 vssd1 vccd1 vccd1 _12172_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_150_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17130__A1 _16039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20390__C _20390_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16980_ _16980_/A _16980_/B _16980_/C vssd1 vssd1 vccd1 vccd1 _16981_/A sky130_fd_sc_hd__nand3_1
XFILLER_123_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15692__A1 _11935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15931_ _15883_/Y _15856_/Y _16043_/A _15930_/X vssd1 vssd1 vccd1 vccd1 _15949_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__15692__B2 _15691_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_822 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16299__D _18130_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16877__A _20972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18650_ _18657_/A _18659_/B _18649_/X vssd1 vssd1 vccd1 vccd1 _18654_/A sky130_fd_sc_hd__a21o_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15862_ _15862_/A vssd1 vssd1 vccd1 vccd1 _15862_/Y sky130_fd_sc_hd__inv_2
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17601_ _17781_/A _17781_/B vssd1 vssd1 vccd1 vccd1 _17605_/B sky130_fd_sc_hd__nand2_2
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14813_ _14813_/A _14813_/B vssd1 vssd1 vccd1 vccd1 _14815_/A sky130_fd_sc_hd__nand2_1
X_18581_ _18576_/Y _18411_/B _18219_/B _18417_/C vssd1 vssd1 vccd1 vccd1 _18582_/C
+ sky130_fd_sc_hd__a22oi_2
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15793_ _15921_/A _15834_/A _15792_/X vssd1 vssd1 vccd1 vccd1 _15793_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_92_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17532_ _17532_/A _17532_/B _17532_/C _17532_/D vssd1 vssd1 vccd1 vccd1 _17532_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14744_ _14745_/A _14741_/Y _14743_/Y vssd1 vssd1 vccd1 vccd1 _14836_/A sky130_fd_sc_hd__o21ai_2
XFILLER_91_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _19016_/A _18093_/C _11956_/C _18093_/D vssd1 vssd1 vccd1 vccd1 _11956_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_83_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17463_ _11904_/X _11905_/X _16579_/X _16580_/X _21011_/A vssd1 vssd1 vccd1 vccd1
+ _17463_/X sky130_fd_sc_hd__o221a_1
XANTENNA__13207__B1 _21580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16944__A1 _15325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11887_ _19202_/D vssd1 vssd1 vccd1 vccd1 _19455_/C sky130_fd_sc_hd__buf_2
X_14675_ _14670_/A _13924_/X _14622_/X _14636_/D vssd1 vssd1 vccd1 vccd1 _14675_/Y
+ sky130_fd_sc_hd__o211ai_2
X_19202_ _19346_/A _19507_/B _19504_/C _19202_/D vssd1 vssd1 vccd1 vccd1 _19211_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16414_ _16414_/A _16414_/B _16414_/C vssd1 vssd1 vccd1 vccd1 _16414_/X sky130_fd_sc_hd__and3_1
X_13626_ _13576_/X _13578_/X _13587_/Y _13588_/X vssd1 vssd1 vccd1 vccd1 _13627_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17394_ _16040_/A _17393_/X _17247_/X vssd1 vssd1 vccd1 vccd1 _17394_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_160_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14844__B _14929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19133_ _18958_/B _19132_/Y _19131_/B vssd1 vssd1 vccd1 vccd1 _19134_/B sky130_fd_sc_hd__a21o_1
XFILLER_160_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ _16316_/Y _16351_/A _15978_/C _20793_/D vssd1 vssd1 vccd1 vccd1 _16345_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13557_ _13558_/A _13558_/B vssd1 vssd1 vccd1 vccd1 _13557_/X sky130_fd_sc_hd__and2_1
XFILLER_185_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19064_ _19044_/X _19046_/X _19074_/A _19074_/B vssd1 vssd1 vccd1 vccd1 _19149_/B
+ sky130_fd_sc_hd__o211ai_2
X_12508_ _12508_/A _12508_/B _12508_/C vssd1 vssd1 vccd1 vccd1 _12509_/A sky130_fd_sc_hd__nand3_1
XFILLER_157_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16276_ _16276_/A vssd1 vssd1 vccd1 vccd1 _16276_/X sky130_fd_sc_hd__buf_2
X_13488_ _13237_/X _13601_/A _13546_/B _13440_/A vssd1 vssd1 vccd1 vccd1 _13492_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_173_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16172__A2 _12876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18015_ _18015_/A _18053_/C _18015_/C vssd1 vssd1 vccd1 vccd1 _18016_/B sky130_fd_sc_hd__nand3_1
XANTENNA__18449__A1 _18795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15227_ _15227_/A _15227_/B vssd1 vssd1 vccd1 vccd1 _15227_/X sky130_fd_sc_hd__xor2_2
X_12439_ _12802_/C vssd1 vssd1 vccd1 vccd1 _12610_/A sky130_fd_sc_hd__buf_2
XANTENNA__21677__B _21677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18332__A _18691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17657__C1 _18305_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12733__A2 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17121__A1 _17732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15158_ _15119_/B _15120_/C _15156_/Y _15157_/X vssd1 vssd1 vccd1 vccd1 _15160_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14109_ _14231_/A _14231_/B _15115_/C _15010_/C _14222_/A vssd1 vssd1 vccd1 vccd1
+ _14115_/B sky130_fd_sc_hd__a32o_1
X_19966_ _20025_/A _19926_/A _19928_/B _19963_/A _19963_/B vssd1 vssd1 vccd1 vccd1
+ _19977_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_113_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15089_ _15089_/A _15089_/B vssd1 vssd1 vccd1 vccd1 _15092_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12380__A _22817_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18917_ _18915_/Y _18916_/Y _18836_/A _18713_/A vssd1 vssd1 vccd1 vccd1 _18917_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_171_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19897_ _19941_/B _18889_/X _18890_/X _19941_/D _19839_/B vssd1 vssd1 vccd1 vccd1
+ _19899_/D sky130_fd_sc_hd__o32a_1
XFILLER_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18848_ _19194_/A _19351_/A _18848_/C _18848_/D vssd1 vssd1 vccd1 vccd1 _18849_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__16002__D _16011_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16937__D _19496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18779_ _18779_/A _18779_/B vssd1 vssd1 vccd1 vccd1 _18779_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19177__A2 _19176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20810_ _20810_/A _20810_/B _20810_/C vssd1 vssd1 vccd1 vccd1 _20812_/C sky130_fd_sc_hd__nand3_1
X_21790_ _21790_/A _21790_/B vssd1 vssd1 vccd1 vccd1 _21790_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_763 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17114__C _17311_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20741_ _20818_/B _20730_/B _20731_/A vssd1 vssd1 vccd1 vccd1 _20741_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14150__A2_N _14147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13749__A1 _13737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20672_ _15941_/A _20611_/Y _20609_/X _20671_/Y vssd1 vssd1 vccd1 vccd1 _20717_/B
+ sky130_fd_sc_hd__o22a_2
X_22411_ _22706_/Q input44/X _22413_/S vssd1 vssd1 vccd1 vccd1 _22412_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_996 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22342_ _22685_/Q _22340_/X _22341_/Y _22289_/B _22684_/Q vssd1 vssd1 vccd1 vccd1
+ _22342_/Y sky130_fd_sc_hd__o32ai_1
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22273_ _22273_/A _22314_/A vssd1 vssd1 vccd1 vccd1 _22301_/B sky130_fd_sc_hd__or2_1
XANTENNA__20247__A1 _15326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21224_ _21621_/C vssd1 vssd1 vccd1 vccd1 _22057_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17112__B2 _17732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18860__A1 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16466__A3 _20255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21155_ _22945_/Q _22946_/Q _21149_/A vssd1 vssd1 vccd1 vccd1 _21155_/X sky130_fd_sc_hd__o21a_1
XFILLER_144_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18860__B2 _11845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20106_ _12329_/X _12803_/X _20086_/Y _20087_/Y vssd1 vssd1 vccd1 vccd1 _20107_/C
+ sky130_fd_sc_hd__a22oi_4
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21086_ _21086_/A _21086_/B _21086_/C _21086_/D vssd1 vssd1 vccd1 vccd1 _21087_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_98_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20037_ _19988_/X _20037_/B _20037_/C vssd1 vssd1 vccd1 vccd1 _20037_/X sky130_fd_sc_hd__and3b_1
XANTENNA__18612__A1 _12170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22849__D _22861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19504__C _19504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14929__B _14929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13437__B1 _21383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20012__A _20012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11634__A _11634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11814_/B _12024_/A _11810_/C vssd1 vssd1 vccd1 vccd1 _12036_/A sky130_fd_sc_hd__nand3_2
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12790_ _12790_/A vssd1 vssd1 vccd1 vccd1 _12929_/A sky130_fd_sc_hd__buf_4
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21988_ _22034_/A _21522_/D _21986_/C _21986_/B vssd1 vssd1 vccd1 vccd1 _21988_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11999__B1 _15633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _18203_/A _17427_/A _11755_/A vssd1 vssd1 vccd1 vccd1 _11741_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_109_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ _20935_/Y _20938_/Y _20933_/Y vssd1 vssd1 vccd1 vccd1 _20939_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17959__C _17959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11672_/A vssd1 vssd1 vccd1 vccd1 _11672_/X sky130_fd_sc_hd__buf_2
X_14460_ _14465_/A _14465_/B _14693_/D vssd1 vssd1 vccd1 vccd1 _14468_/B sky130_fd_sc_hd__nand3_2
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13411_ _13405_/Y _13406_/Y _21665_/D _21299_/B vssd1 vssd1 vccd1 vccd1 _13416_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14391_ _14413_/A vssd1 vssd1 vccd1 vccd1 _14391_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22609_ _22609_/A vssd1 vssd1 vccd1 vccd1 _22793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12465__A _20086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16130_ _16130_/A _16130_/B _20745_/C vssd1 vssd1 vccd1 vccd1 _16131_/B sky130_fd_sc_hd__and3_1
X_13342_ _21173_/C _21173_/A vssd1 vssd1 vccd1 vccd1 _13343_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16154__A2 _16130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15776__A _15776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16061_ _16080_/A _16080_/C _11845_/X _16177_/A vssd1 vssd1 vccd1 vccd1 _16064_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_13273_ _13273_/A _13273_/B vssd1 vssd1 vccd1 vccd1 _13361_/A sky130_fd_sc_hd__nand2_1
XFILLER_154_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12224_ _12054_/X _12056_/Y _12039_/Y _12081_/A vssd1 vssd1 vccd1 vccd1 _12227_/B
+ sky130_fd_sc_hd__a2bb2oi_1
X_15012_ _15080_/A _15080_/B vssd1 vssd1 vccd1 vccd1 _15013_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12912__B _20793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19820_ _19880_/C vssd1 vssd1 vccd1 vccd1 _19820_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12155_ _11585_/A _11415_/A _12154_/Y vssd1 vssd1 vccd1 vccd1 _12156_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11809__A _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18851__B2 _17434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11931__A1_N _11693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19751_ _19569_/A _19669_/Y _19750_/X vssd1 vssd1 vccd1 vccd1 _19751_/Y sky130_fd_sc_hd__o21ai_1
X_16963_ _16773_/B _16954_/A _16760_/X _16494_/X vssd1 vssd1 vccd1 vccd1 _16967_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_12086_ _12086_/A _12086_/B _12086_/C vssd1 vssd1 vccd1 vccd1 _18239_/B sky130_fd_sc_hd__nand3_2
XANTENNA__11528__B _18691_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18702_ _18702_/A _18702_/B _18702_/C vssd1 vssd1 vccd1 vccd1 _18715_/A sky130_fd_sc_hd__nand3_1
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18603__A1 _19443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15914_ _15914_/A _16414_/B vssd1 vssd1 vccd1 vccd1 _15915_/C sky130_fd_sc_hd__nand2_1
X_19682_ _19682_/A _19682_/B vssd1 vssd1 vccd1 vccd1 _19761_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16894_ _16397_/X _15630_/X _16652_/A vssd1 vssd1 vccd1 vccd1 _16894_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16400__A _16400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20410__A1 _20378_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18633_ _18633_/A _18633_/B vssd1 vssd1 vccd1 vccd1 _18633_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _15752_/X _15753_/Y _15864_/A _15709_/Y vssd1 vssd1 vccd1 vccd1 _15845_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11544__A _15624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18564_ _18564_/A _18564_/B _18564_/C vssd1 vssd1 vccd1 vccd1 _18761_/A sky130_fd_sc_hd__nand3_2
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _15776_/A _15776_/B _20134_/A _15776_/D vssd1 vssd1 vccd1 vccd1 _15780_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _12988_/A _12988_/B _12988_/C vssd1 vssd1 vccd1 vccd1 _13036_/A sky130_fd_sc_hd__or3_2
XFILLER_33_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17515_ _17494_/A _17375_/A _17514_/Y vssd1 vssd1 vccd1 vccd1 _17515_/X sky130_fd_sc_hd__a21o_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14727_ _14727_/A _14727_/B _14727_/C _14892_/D vssd1 vssd1 vccd1 vccd1 _14727_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__16917__A1 _15580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18495_ _18495_/A _18495_/B vssd1 vssd1 vccd1 vccd1 _19329_/B sky130_fd_sc_hd__nand2_1
X_11939_ _12111_/A _11936_/Y _11938_/Y vssd1 vssd1 vccd1 vccd1 _11943_/A sky130_fd_sc_hd__o21ai_1
XFILLER_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20576__B _20576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17446_ _17523_/B _17449_/C _17441_/X _17445_/X vssd1 vssd1 vccd1 vccd1 _17457_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_21_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14658_ _14530_/A _14530_/B _14541_/B _14655_/Y _14752_/A vssd1 vssd1 vccd1 vccd1
+ _14758_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_162_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ _13608_/A _13608_/C _13608_/B vssd1 vssd1 vccd1 vccd1 _13609_/Y sky130_fd_sc_hd__a21oi_1
X_17377_ _17260_/B _17260_/C _17260_/A vssd1 vssd1 vccd1 vccd1 _17377_/Y sky130_fd_sc_hd__a21oi_1
X_14589_ _14785_/A vssd1 vssd1 vccd1 vccd1 _15056_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12375__A _12519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19116_ _19116_/A _19116_/B vssd1 vssd1 vccd1 vccd1 _19303_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16328_ _16328_/A _22701_/Q vssd1 vssd1 vccd1 vccd1 _16580_/A sky130_fd_sc_hd__nand2_2
XFILLER_119_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12094__B _19358_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_955 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19047_ _19507_/A _19047_/B vssd1 vssd1 vccd1 vccd1 _19357_/A sky130_fd_sc_hd__nand2_1
X_16259_ _19016_/A vssd1 vssd1 vccd1 vccd1 _18848_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_173_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18842__A1 _18259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11390__A1 _15484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11438__B _11438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19949_ _19949_/A _19949_/B vssd1 vssd1 vccd1 vccd1 _20037_/C sky130_fd_sc_hd__nor2_1
XANTENNA__19605__B _19605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21729__A1 _21853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22960_ _22964_/CLK _22960_/D vssd1 vssd1 vccd1 vccd1 _22960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_983 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21911_ _21911_/A vssd1 vssd1 vccd1 vccd1 _21911_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22891_ _22952_/CLK _22891_/D vssd1 vssd1 vccd1 vccd1 _22891_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11693__A2 _11563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15813__D1 _11779_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21842_ _21269_/A _21341_/X _21841_/B _21841_/C vssd1 vssd1 vccd1 vccd1 _21842_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19340__B _19340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21773_ _21789_/B _21778_/D vssd1 vssd1 vccd1 vccd1 _21773_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14765__A _14765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17141__A _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20724_ _20479_/Y _20614_/Y _20615_/Y _20616_/X vssd1 vssd1 vccd1 vccd1 _20724_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_928 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20655_ _20454_/B _20449_/Y _20650_/A _20650_/B _20454_/C vssd1 vssd1 vccd1 vccd1
+ _20656_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20468__A1 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20586_ _20586_/A _20586_/B _20586_/C vssd1 vssd1 vccd1 vccd1 _20596_/A sky130_fd_sc_hd__nand3_1
XANTENNA__18530__B1 _19316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22325_ _22325_/A _22325_/B _22325_/C vssd1 vssd1 vccd1 vccd1 _22327_/A sky130_fd_sc_hd__and3_1
XFILLER_165_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22256_ _22142_/A _22142_/B _22143_/X vssd1 vssd1 vccd1 vccd1 _22256_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21207_ _21207_/A vssd1 vssd1 vccd1 vccd1 _21615_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22187_ _22220_/A _22265_/C _22186_/X _22183_/Y vssd1 vssd1 vccd1 vccd1 _22188_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_78_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21138_ _21138_/A _21138_/B _21138_/C vssd1 vssd1 vccd1 vccd1 _21138_/X sky130_fd_sc_hd__and3_1
XFILLER_94_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13960_ _14510_/C vssd1 vssd1 vccd1 vccd1 _14911_/A sky130_fd_sc_hd__clkbuf_2
X_21069_ _21066_/X _21067_/X _21079_/B vssd1 vssd1 vccd1 vccd1 _21070_/B sky130_fd_sc_hd__o21ai_1
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12911_ _15988_/B _16078_/B _12680_/X _16498_/A _20593_/C vssd1 vssd1 vccd1 vccd1
+ _12912_/A sky130_fd_sc_hd__a32o_1
XFILLER_171_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13891_ _13891_/A vssd1 vssd1 vccd1 vccd1 _14021_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15630_ _15647_/A _16431_/A _15912_/C _16361_/A vssd1 vssd1 vccd1 vccd1 _15630_/X
+ sky130_fd_sc_hd__and4_4
XFILLER_34_508 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _12855_/A _12855_/B vssd1 vssd1 vccd1 vccd1 _12859_/B sky130_fd_sc_hd__nand2_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _12111_/A _15569_/A _15568_/A vssd1 vssd1 vccd1 vccd1 _15565_/C sky130_fd_sc_hd__o21ai_2
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12773_/A vssd1 vssd1 vccd1 vccd1 _12774_/A sky130_fd_sc_hd__buf_4
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17273_/A _17307_/C _17304_/B vssd1 vssd1 vccd1 vccd1 _17301_/C sky130_fd_sc_hd__a21o_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_552 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14512_/A _14512_/B _14512_/C _15058_/C vssd1 vssd1 vccd1 vccd1 _14515_/C
+ sky130_fd_sc_hd__nand4_2
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _11859_/X _11861_/X _19358_/A _19358_/B vssd1 vssd1 vccd1 vccd1 _18451_/A
+ sky130_fd_sc_hd__o211ai_4
X_11724_ _11708_/Y _11935_/C _19320_/A _11664_/D vssd1 vssd1 vccd1 vccd1 _11724_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_9_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _12758_/A _16786_/A _15439_/A vssd1 vssd1 vccd1 vccd1 _15567_/A sky130_fd_sc_hd__o21ai_2
XFILLER_15_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12907__B _16078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17231_ _17184_/A _17184_/B _17184_/C vssd1 vssd1 vccd1 vccd1 _17231_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14386__A1 _20069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14443_ _22658_/A vssd1 vssd1 vccd1 vccd1 _14443_/X sky130_fd_sc_hd__clkbuf_2
X_11655_ _22960_/Q vssd1 vssd1 vccd1 vccd1 _15435_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_187_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14386__B2 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17162_ _16954_/A _16954_/B _16959_/B _16959_/A vssd1 vssd1 vccd1 vccd1 _17162_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_156_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12936__A2 _12721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11586_ _11589_/A _11583_/Y _11361_/A _18156_/A vssd1 vssd1 vccd1 vccd1 _11591_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_14374_ _14369_/X _14370_/X _14351_/X _21580_/B _14373_/X vssd1 vssd1 vccd1 vccd1
+ _14374_/X sky130_fd_sc_hd__a221o_1
XFILLER_10_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16603__B1_N _16600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16113_ _16069_/X _16113_/B _16113_/C _16150_/B vssd1 vssd1 vccd1 vccd1 _16169_/C
+ sky130_fd_sc_hd__nand4b_2
XFILLER_6_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13325_ _13318_/Y _13321_/X _13322_/Y _13324_/Y vssd1 vssd1 vccd1 vccd1 _13354_/B
+ sky130_fd_sc_hd__o211ai_4
X_17093_ _17087_/B _17083_/X _17460_/A _17085_/Y _17520_/A vssd1 vssd1 vccd1 vccd1
+ _17094_/C sky130_fd_sc_hd__o311ai_4
XFILLER_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16044_ _16200_/C _16414_/C vssd1 vssd1 vccd1 vccd1 _16044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13256_ _13230_/X _13623_/A _21584_/C _13240_/A vssd1 vssd1 vccd1 vccd1 _13662_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _16940_/A vssd1 vssd1 vccd1 vccd1 _12207_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11539__A _15357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ _21495_/B _22845_/Q vssd1 vssd1 vccd1 vccd1 _13192_/B sky130_fd_sc_hd__and2_1
XANTENNA__13457__C _21498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19803_ _19735_/C _19736_/B _19804_/A _19804_/B vssd1 vssd1 vccd1 vccd1 _19872_/A
+ sky130_fd_sc_hd__a22o_1
X_12138_ _12138_/A _12138_/B _12138_/C vssd1 vssd1 vccd1 vccd1 _12139_/A sky130_fd_sc_hd__nand3_1
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17995_ _17945_/A _17945_/B _17899_/B _18020_/C vssd1 vssd1 vccd1 vccd1 _17996_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13649__B1 _21195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17226__A _17226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19734_ _19735_/B _19726_/A _19735_/A vssd1 vssd1 vccd1 vccd1 _19736_/A sky130_fd_sc_hd__a21o_1
X_16946_ _16946_/A vssd1 vssd1 vccd1 vccd1 _16946_/X sky130_fd_sc_hd__clkbuf_2
X_12069_ _11918_/B _12069_/B _16130_/B _19046_/C vssd1 vssd1 vccd1 vccd1 _12069_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19665_ _19814_/A _19814_/B _19813_/B _19813_/A vssd1 vssd1 vccd1 vccd1 _19670_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_93_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16877_ _20972_/A vssd1 vssd1 vccd1 vccd1 _20936_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18616_ _18616_/A _18616_/B vssd1 vssd1 vccd1 vccd1 _18616_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11274__A _22799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _15828_/A vssd1 vssd1 vccd1 vccd1 _15828_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19596_ _19842_/A _19596_/B _19596_/C _19774_/D vssd1 vssd1 vccd1 vccd1 _19684_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18547_ _18553_/A _18553_/B _18546_/C vssd1 vssd1 vccd1 vccd1 _18548_/B sky130_fd_sc_hd__a21o_1
XANTENNA__19001__A1 _19000_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15759_ _15758_/A _15758_/B _15758_/C vssd1 vssd1 vccd1 vccd1 _15759_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_178_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18478_ _18765_/A _18478_/B _18478_/C vssd1 vssd1 vccd1 vccd1 _18565_/B sky130_fd_sc_hd__nand3_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17429_ _17427_/X _17111_/A _17564_/A vssd1 vssd1 vccd1 vccd1 _17431_/D sky130_fd_sc_hd__o21ai_2
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20440_ _20563_/A _20562_/C vssd1 vssd1 vccd1 vccd1 _20441_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12927__A2 _12774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22952__D _22952_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20371_ _20371_/A _20371_/B vssd1 vssd1 vccd1 vccd1 _20371_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22110_ _22105_/X _22179_/A _22220_/A _22173_/B _22109_/Y vssd1 vssd1 vccd1 vccd1
+ _22113_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12552__B _12567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22041_ _22041_/A _22041_/B _22041_/C vssd1 vssd1 vccd1 vccd1 _22105_/A sky130_fd_sc_hd__nand3_1
XFILLER_88_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16826__B1 _16452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21584__C _21584_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1097 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16040__A _16040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22943_ _22943_/CLK _22943_/D vssd1 vssd1 vccd1 vccd1 _22943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19351__A _19351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22874_ _22915_/CLK _22874_/D vssd1 vssd1 vccd1 vccd1 _22874_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20928__C _20928_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21825_ _21825_/A _21825_/B _22677_/Q vssd1 vssd1 vccd1 vccd1 _21922_/A sky130_fd_sc_hd__nand3_1
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14495__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_658 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11912__A _11912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21756_ _21755_/Y _21582_/B _21937_/A vssd1 vssd1 vccd1 vccd1 _22058_/A sky130_fd_sc_hd__a21boi_2
XFILLER_196_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14368__A1 _22700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20707_ _20706_/X _20690_/X _20796_/B _20699_/A vssd1 vssd1 vccd1 vccd1 _20709_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21687_ _21809_/A _21814_/A _21687_/C vssd1 vssd1 vccd1 vccd1 _21688_/C sky130_fd_sc_hd__nand3_1
XFILLER_138_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11440_ _15633_/A vssd1 vssd1 vccd1 vccd1 _15714_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22862__D _22874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20638_ _12606_/X _12607_/X _20734_/B _20734_/C _20178_/A vssd1 vssd1 vccd1 vccd1
+ _20638_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16109__A2 _12501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14942__B _14942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11371_ _11371_/A _11371_/B _15357_/A vssd1 vssd1 vccd1 vccd1 _11371_/X sky130_fd_sc_hd__and3_1
XANTENNA__15317__B1 _12577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20569_ _20511_/A _20511_/B _20511_/C _20511_/D vssd1 vssd1 vccd1 vccd1 _20569_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_152_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22308_ _22308_/A _22308_/B _22308_/C _22309_/B vssd1 vssd1 vccd1 vccd1 _22310_/A
+ sky130_fd_sc_hd__or4_1
X_13110_ _13143_/A _13143_/B _13112_/D vssd1 vssd1 vccd1 vccd1 _13110_/Y sky130_fd_sc_hd__nand3_2
XFILLER_192_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14090_ _14167_/A _14167_/C vssd1 vssd1 vccd1 vccd1 _14090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13879__B1 _13873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ _13045_/A _13045_/B vssd1 vssd1 vccd1 vccd1 _13041_/Y sky130_fd_sc_hd__nand2_4
XFILLER_65_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17609__A2 _17227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22239_ _22240_/B _22240_/C _22240_/A vssd1 vssd1 vccd1 vccd1 _22241_/A sky130_fd_sc_hd__a21oi_1
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12551__B1 _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input46_A wb_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16800_ _16177_/A _16799_/X _16782_/X _16787_/Y _16792_/B vssd1 vssd1 vccd1 vccd1
+ _16800_/X sky130_fd_sc_hd__o311a_1
XFILLER_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17780_ _17600_/A _17600_/B _17704_/A vssd1 vssd1 vccd1 vccd1 _17780_/X sky130_fd_sc_hd__o21a_1
X_14992_ _14961_/B _14961_/A _14971_/Y vssd1 vssd1 vccd1 vccd1 _15031_/A sky130_fd_sc_hd__o21ai_1
XFILLER_115_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16731_ _16564_/B _20792_/A _20792_/B _20793_/D _16106_/B vssd1 vssd1 vccd1 vccd1
+ _16732_/B sky130_fd_sc_hd__a32o_2
X_13943_ _13911_/X _13942_/Y _13903_/Y vssd1 vssd1 vccd1 vccd1 _13947_/A sky130_fd_sc_hd__o21a_1
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_655 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19450_ _19442_/Y _19445_/Y _19449_/Y vssd1 vssd1 vccd1 vccd1 _19452_/A sky130_fd_sc_hd__o21a_1
XFILLER_90_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16662_ _16426_/X _16664_/B _16664_/C _16438_/A vssd1 vssd1 vccd1 vccd1 _17064_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__16100__D _16100_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13874_ _13745_/B _13745_/C _13736_/C _14122_/A vssd1 vssd1 vccd1 vccd1 _13876_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_47_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18401_ _18309_/B _18442_/B _18402_/A _18402_/B vssd1 vssd1 vccd1 vccd1 _18401_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_90_945 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15613_ _20101_/A vssd1 vssd1 vccd1 vccd1 _16715_/A sky130_fd_sc_hd__clkbuf_4
X_19381_ _19206_/Y _19211_/X _19209_/Y _19208_/A vssd1 vssd1 vccd1 vccd1 _19389_/C
+ sky130_fd_sc_hd__o31a_1
X_12825_ _22698_/Q vssd1 vssd1 vccd1 vccd1 _16322_/A sky130_fd_sc_hd__buf_2
XFILLER_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16593_ _16598_/A _16598_/B _16599_/C _16599_/B vssd1 vssd1 vccd1 vccd1 _16594_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18332_ _18691_/A _18691_/B vssd1 vssd1 vccd1 vccd1 _18492_/A sky130_fd_sc_hd__nand2_1
XFILLER_188_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15544_ _15838_/A vssd1 vssd1 vccd1 vccd1 _18203_/C sky130_fd_sc_hd__buf_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _15746_/B _20390_/B vssd1 vssd1 vccd1 vccd1 _12757_/A sky130_fd_sc_hd__nand2_1
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18263_ _18257_/B _18598_/B _12258_/A _18247_/A _18257_/Y vssd1 vssd1 vccd1 vccd1
+ _18263_/X sky130_fd_sc_hd__o221a_1
X_11707_ _11707_/A vssd1 vssd1 vccd1 vccd1 _15458_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15475_ _12202_/A _12202_/B _12672_/A _15755_/A vssd1 vssd1 vccd1 vccd1 _15479_/A
+ sky130_fd_sc_hd__a211o_2
X_12687_ _20357_/B _12687_/B vssd1 vssd1 vccd1 vccd1 _20355_/D sky130_fd_sc_hd__and2_2
XANTENNA__20854__B _20854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17214_ _16889_/B _16673_/A _16665_/X vssd1 vssd1 vccd1 vccd1 _17215_/A sky130_fd_sc_hd__a21oi_1
X_14426_ _22718_/Q _14418_/X _14351_/A _22750_/Q _14425_/X vssd1 vssd1 vccd1 vccd1
+ _14426_/X sky130_fd_sc_hd__a221o_1
X_18194_ _11502_/X _11503_/X _17380_/A _17381_/X _18200_/A vssd1 vssd1 vccd1 vccd1
+ _18194_/Y sky130_fd_sc_hd__o221ai_4
X_11638_ _18330_/A vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__buf_2
XFILLER_129_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18324__B _22796_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17145_ _17145_/A _17145_/B vssd1 vssd1 vccd1 vccd1 _17145_/Y sky130_fd_sc_hd__nand2_2
X_14357_ _16322_/A _14344_/X _14351_/X _21329_/B _14356_/X vssd1 vssd1 vccd1 vccd1
+ _14357_/X sky130_fd_sc_hd__a221o_1
X_11569_ _15476_/A vssd1 vssd1 vccd1 vccd1 _19318_/A sky130_fd_sc_hd__buf_4
XANTENNA__12653__A _16498_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1042 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13308_ _21312_/B vssd1 vssd1 vccd1 vccd1 _13521_/B sky130_fd_sc_hd__buf_2
XFILLER_7_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20852__A1 _12671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17076_ _17076_/A _17076_/B _17076_/C vssd1 vssd1 vccd1 vccd1 _17077_/B sky130_fd_sc_hd__nand3_1
XFILLER_170_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20870__A _20870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14288_ _14288_/A _14288_/B _14288_/C vssd1 vssd1 vccd1 vccd1 _14289_/B sky130_fd_sc_hd__nand3_1
X_16027_ _15945_/A _15945_/B _15917_/X _16026_/Y vssd1 vssd1 vccd1 vccd1 _16043_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_143_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13239_ _13234_/A _13234_/B _13157_/A vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__o21ai_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17978_ _19896_/A vssd1 vssd1 vccd1 vccd1 _19419_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18025__A2 _18023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16929_ _16930_/A _17341_/A _16930_/C vssd1 vssd1 vccd1 vccd1 _16988_/A sky130_fd_sc_hd__a21o_1
X_19717_ _16015_/X _19838_/A _19793_/A _19621_/Y _19715_/X vssd1 vssd1 vccd1 vccd1
+ _19719_/B sky130_fd_sc_hd__o311a_1
XFILLER_133_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12845__B2 _16178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16036__B2 _15937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19773__A2 _19517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19648_ _19488_/A _19636_/X _19637_/Y _19635_/A _19724_/B vssd1 vssd1 vccd1 vccd1
+ _19649_/C sky130_fd_sc_hd__o2111ai_2
XANTENNA__19602__C _19602_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22109__A1 _21376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20748__C _20748_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19579_ _19682_/A _19682_/B _19569_/A vssd1 vssd1 vccd1 vccd1 _19880_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__15795__B1 _15891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21610_ _21610_/A _21610_/B vssd1 vssd1 vccd1 vccd1 _21614_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13650__C _21195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22590_ _22590_/A vssd1 vssd1 vccd1 vccd1 _22784_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17122__C _17122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21541_ _21531_/A _21531_/C _21539_/Y vssd1 vssd1 vccd1 vccd1 _21541_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21472_ _22733_/Q vssd1 vssd1 vccd1 vccd1 _21583_/D sky130_fd_sc_hd__clkinv_2
XFILLER_53_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14762__B _14929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20423_ _20423_/A _20423_/B _20423_/C vssd1 vssd1 vccd1 vccd1 _20549_/D sky130_fd_sc_hd__nand3_4
XANTENNA__18497__C1 _16564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15577__C _20390_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20354_ _12988_/B _16566_/A _16568_/A _20358_/A vssd1 vssd1 vccd1 vccd1 _20354_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__20780__A _21019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19346__A _19346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21595__B _21595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20285_ _20401_/A _20401_/B _20269_/X _20274_/Y vssd1 vssd1 vccd1 vccd1 _20286_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_161_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22024_ _22024_/A _22024_/B vssd1 vssd1 vccd1 vccd1 _22024_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20071__A2 _20064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13089__A1 _13050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22857__D _22869_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22926_ _22948_/CLK _22926_/D vssd1 vssd1 vccd1 vccd1 _22926_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17313__B _17313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22857_ _22943_/CLK _22869_/Q vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15250__A2 _15247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12610_ _12610_/A vssd1 vssd1 vccd1 vccd1 _20576_/B sky130_fd_sc_hd__buf_2
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21808_ _21805_/X _21677_/A _21797_/Y _21913_/A vssd1 vssd1 vccd1 vccd1 _21808_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18128__C _18128_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17527__A1 _15940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13590_ _21445_/C _21489_/A _13586_/Y _13528_/X vssd1 vssd1 vccd1 vccd1 _13597_/A
+ sky130_fd_sc_hd__a22o_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17527__B2 _17636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22788_ _22797_/CLK _22788_/D vssd1 vssd1 vccd1 vccd1 _22788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_680 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _12553_/A _12789_/A _12536_/Y _12540_/X vssd1 vssd1 vccd1 vccd1 _12543_/C
+ sky130_fd_sc_hd__o22ai_4
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16735__C1 _16842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21739_ _22041_/A _21739_/B _21739_/C vssd1 vssd1 vccd1 vccd1 _21868_/A sky130_fd_sc_hd__nand3_1
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14953__A _14953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15260_ _15260_/A _15260_/B vssd1 vssd1 vccd1 vccd1 _15263_/A sky130_fd_sc_hd__or2_1
XFILLER_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12472_ _12520_/A vssd1 vssd1 vccd1 vccd1 _12669_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_61_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16750__A2 _16740_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14211_ _14595_/B vssd1 vssd1 vccd1 vccd1 _15004_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_137_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11423_ _11423_/A vssd1 vssd1 vccd1 vccd1 _12154_/C sky130_fd_sc_hd__buf_2
XANTENNA__13569__A _21621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15191_ _15238_/B _15190_/X _15154_/X _15156_/Y vssd1 vssd1 vccd1 vccd1 _15194_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11354_ _11334_/X _11423_/A _11720_/A vssd1 vssd1 vccd1 vccd1 _11593_/A sky130_fd_sc_hd__and3b_1
X_14142_ _13819_/Y _13829_/Y _13824_/X vssd1 vssd1 vccd1 vccd1 _14146_/A sky130_fd_sc_hd__a21o_1
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18950_ _18950_/A _18952_/A vssd1 vssd1 vccd1 vccd1 _18951_/C sky130_fd_sc_hd__nand2_1
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11285_ _11285_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__nand2_2
X_14073_ _14073_/A vssd1 vssd1 vccd1 vccd1 _14619_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12524__B1 _12493_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17901_ _17842_/A _17842_/B _17900_/X vssd1 vssd1 vccd1 vccd1 _18020_/B sky130_fd_sc_hd__a21oi_2
XFILLER_152_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13024_ _13024_/A _13024_/B _15746_/B vssd1 vssd1 vccd1 vccd1 _13024_/X sky130_fd_sc_hd__and3_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18881_ _18881_/A vssd1 vssd1 vccd1 vccd1 _18881_/X sky130_fd_sc_hd__buf_2
XFILLER_126_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17832_ _17871_/A _17897_/A vssd1 vssd1 vccd1 vccd1 _17835_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17463__B1 _16579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17763_ _17687_/A _17687_/B _17687_/C vssd1 vssd1 vccd1 vccd1 _17763_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__19204__A1 _18371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19204__B2 _12018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14975_ _14912_/A _14912_/B _14909_/Y vssd1 vssd1 vccd1 vccd1 _14977_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__16018__A1 _15812_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19502_ _19368_/B _19355_/Y _19352_/X _19215_/X vssd1 vssd1 vccd1 vccd1 _19503_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_16714_ _16714_/A vssd1 vssd1 vccd1 vccd1 _16714_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13926_ _13857_/X _13725_/Y _22859_/D _13728_/A vssd1 vssd1 vccd1 vccd1 _13926_/Y
+ sky130_fd_sc_hd__o211ai_4
X_17694_ _17626_/B _17626_/A _17627_/X vssd1 vssd1 vccd1 vccd1 _17695_/A sky130_fd_sc_hd__o21a_1
XANTENNA__17766__A1 _17669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16569__A2 _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19433_ _19429_/Y _19131_/A _19432_/Y vssd1 vssd1 vccd1 vccd1 _19439_/A sky130_fd_sc_hd__o21bai_1
X_16645_ _16895_/A _16895_/B _16644_/C vssd1 vssd1 vccd1 vccd1 _16645_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15777__B1 _11506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13857_ _13963_/A vssd1 vssd1 vccd1 vccd1 _13857_/X sky130_fd_sc_hd__buf_4
XFILLER_16_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19364_ _11639_/X _17526_/X _19215_/X _19352_/X vssd1 vssd1 vccd1 vccd1 _19364_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_16_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ _12701_/A _15335_/A _12803_/A vssd1 vssd1 vccd1 vccd1 _12808_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16576_ _20584_/A _20584_/B vssd1 vssd1 vccd1 vccd1 _20697_/C sky130_fd_sc_hd__nand2_1
X_13788_ _14054_/A _14055_/B _14165_/A vssd1 vssd1 vccd1 vccd1 _14049_/B sky130_fd_sc_hd__o21a_1
XFILLER_188_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18315_ _18678_/C _18324_/A vssd1 vssd1 vccd1 vccd1 _18691_/A sky130_fd_sc_hd__nand2_2
X_15527_ _15527_/A vssd1 vssd1 vccd1 vccd1 _16265_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19295_ _19295_/A _19295_/B vssd1 vssd1 vccd1 vccd1 _19301_/B sky130_fd_sc_hd__nand2_1
XFILLER_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ _12739_/A _12739_/B _12739_/C vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__nand3_2
XFILLER_148_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16781__C _18192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18246_ _18246_/A _18246_/B vssd1 vssd1 vccd1 vccd1 _18247_/A sky130_fd_sc_hd__nand2_1
XFILLER_187_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15458_ _15458_/A vssd1 vssd1 vccd1 vccd1 _15810_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__14201__B1 _14786_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16741__A2 _16842_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14409_ _22712_/Q _14403_/X _14396_/X _22744_/Q _14408_/X vssd1 vssd1 vccd1 vccd1
+ _14409_/X sky130_fd_sc_hd__a221o_1
X_18177_ _18184_/A _18184_/B vssd1 vssd1 vccd1 vccd1 _18177_/X sky130_fd_sc_hd__and2_1
XFILLER_190_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15389_ _15389_/A _15389_/B _15389_/C vssd1 vssd1 vccd1 vccd1 _15389_/X sky130_fd_sc_hd__and3_1
XANTENNA__12383__A _15352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17128_ _19694_/B _17128_/B _17407_/A _19496_/A vssd1 vssd1 vccd1 vccd1 _17128_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__20825__A1 _20759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12814__C _20341_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13198__B _21609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18494__A2 _19624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15694__A _15694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14504__A1 _14818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17059_ _17213_/B vssd1 vssd1 vccd1 vccd1 _17060_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__19166__A _19168_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14504__B2 _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20070_ _20834_/A _20835_/A vssd1 vssd1 vccd1 vccd1 _20314_/B sky130_fd_sc_hd__or2_1
XANTENNA__11869__A2 _11308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22940__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20759__B _20759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20972_ _20972_/A _20972_/B _21011_/B _20972_/D vssd1 vssd1 vccd1 vccd1 _20975_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_39_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22711_ _22743_/CLK _22711_/D vssd1 vssd1 vccd1 vccd1 _22711_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__20478__C _20478_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17133__B _17631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16965__C1 _20249_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11462__A _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15232__A2 _15205_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22642_ _22642_/A vssd1 vssd1 vccd1 vccd1 _22808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15869__A _17739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22573_ _22573_/A vssd1 vssd1 vccd1 vccd1 _22777_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14991__A1 _14990_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18245__A _18259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21524_ _21524_/A _21524_/B vssd1 vssd1 vccd1 vccd1 _21539_/B sky130_fd_sc_hd__nand2_2
XFILLER_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21455_ _21606_/A vssd1 vssd1 vccd1 vccd1 _21455_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20406_ _20395_/A _20395_/B _20388_/Y _20405_/Y vssd1 vssd1 vccd1 vccd1 _20407_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_181_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21386_ _21386_/A _21386_/B _21386_/C vssd1 vssd1 vccd1 vccd1 _21386_/X sky130_fd_sc_hd__and3_1
XFILLER_162_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20337_ _20337_/A vssd1 vssd1 vccd1 vccd1 _20403_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19507__C _19507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20268_ _20268_/A _20268_/B _20268_/C vssd1 vssd1 vccd1 vccd1 _20408_/A sky130_fd_sc_hd__nand3_1
XFILLER_103_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22033__A3 _21724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22007_ _22007_/A _22007_/B vssd1 vssd1 vccd1 vccd1 _22008_/B sky130_fd_sc_hd__nand2_1
XFILLER_163_67 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17445__B1 _16016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14013__A _14013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20199_ _20077_/B _20293_/A _20077_/A vssd1 vssd1 vccd1 vccd1 _20199_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_193_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13852__A _22869_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _14758_/C _14660_/B _14759_/Y vssd1 vssd1 vccd1 vccd1 _14761_/B sky130_fd_sc_hd__o21a_1
XFILLER_91_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ _12137_/A _11970_/Y _11984_/B vssd1 vssd1 vccd1 vccd1 _11972_/Y sky130_fd_sc_hd__a21oi_4
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20388__C _20388_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ _14191_/B vssd1 vssd1 vccd1 vccd1 _14273_/C sky130_fd_sc_hd__buf_2
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22909_ _22915_/CLK _22909_/D vssd1 vssd1 vccd1 vccd1 _22909_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _14568_/B _14793_/A _14685_/Y _14686_/X vssd1 vssd1 vccd1 vccd1 _14695_/A
+ sky130_fd_sc_hd__o211ai_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12468__A _20210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__A _11372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16430_ _16652_/A _16444_/A _16400_/X _16397_/X vssd1 vssd1 vccd1 vccd1 _16439_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_13642_ _13637_/Y _13640_/Y _13641_/Y vssd1 vssd1 vccd1 vccd1 _13643_/C sky130_fd_sc_hd__a21o_1
XFILLER_32_628 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20685__A _20685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16361_/A vssd1 vssd1 vccd1 vccd1 _20793_/C sky130_fd_sc_hd__clkbuf_4
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13785__A2 _14489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13573_ _13573_/A _21944_/A _13664_/B _13618_/A vssd1 vssd1 vccd1 vccd1 _13618_/B
+ sky130_fd_sc_hd__nand4_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18100_ _12146_/Y _12148_/Y _18841_/B _18116_/D vssd1 vssd1 vccd1 vccd1 _18102_/A
+ sky130_fd_sc_hd__o211ai_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _11935_/B _16178_/A _15461_/A vssd1 vssd1 vccd1 vccd1 _15313_/C sky130_fd_sc_hd__o21ai_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19080_ _19080_/A vssd1 vssd1 vccd1 vccd1 _19254_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ _12421_/A _12550_/A _12493_/Y vssd1 vssd1 vccd1 vccd1 _12540_/C sky130_fd_sc_hd__a21o_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16292_ _16286_/Y _16287_/Y _16288_/Y _16291_/Y vssd1 vssd1 vccd1 vccd1 _16370_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__15498__B _15498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18031_ _18025_/X _18029_/X _18030_/C _18030_/Y vssd1 vssd1 vccd1 vccd1 _18033_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__22108__C _22108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15243_ _15243_/A _15243_/B vssd1 vssd1 vccd1 vccd1 _15244_/B sky130_fd_sc_hd__xor2_1
XANTENNA__18305__D _18305_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ _12455_/A vssd1 vssd1 vccd1 vccd1 _12455_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20807__A1 _20178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11406_ _22957_/Q vssd1 vssd1 vccd1 vccd1 _11407_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16106__C _16106_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18476__A2 _18459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15174_ _15174_/A _15174_/B vssd1 vssd1 vccd1 vccd1 _15180_/B sky130_fd_sc_hd__nand2_2
XFILLER_67_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12386_ _12421_/A _12550_/A _16319_/C _12387_/B vssd1 vssd1 vccd1 vccd1 _12386_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__16487__A1 _16100_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14125_ _14184_/C vssd1 vssd1 vccd1 vccd1 _14693_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_181_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11337_ _12210_/A vssd1 vssd1 vccd1 vccd1 _15539_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_125_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19982_ _19983_/A _18778_/D _19941_/D _19987_/B _19946_/C vssd1 vssd1 vccd1 vccd1
+ _19995_/A sky130_fd_sc_hd__o41a_1
XFILLER_126_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15695__C1 _19012_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18933_ _18933_/A _18933_/B _18933_/C vssd1 vssd1 vccd1 vccd1 _18933_/X sky130_fd_sc_hd__and3_1
XFILLER_140_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14056_ _13807_/Y _13808_/Y _13830_/Y _13837_/Y vssd1 vssd1 vccd1 vccd1 _14169_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22963__CLK _22964_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13007_ _13007_/A _13007_/B _13007_/C _13007_/D vssd1 vssd1 vccd1 vccd1 _13012_/A
+ sky130_fd_sc_hd__nand4_1
X_18864_ _19507_/D vssd1 vssd1 vccd1 vccd1 _19602_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_67_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17815_ _19768_/D vssd1 vssd1 vccd1 vccd1 _19896_/B sky130_fd_sc_hd__clkbuf_2
X_18795_ _18795_/A vssd1 vssd1 vccd1 vccd1 _18795_/X sky130_fd_sc_hd__buf_2
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13762__A _13948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20579__B _20579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17746_ _17745_/X _17826_/B _17744_/A vssd1 vssd1 vccd1 vccd1 _17746_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17234__A _17234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14958_ _14959_/B _14959_/C _14959_/A vssd1 vssd1 vccd1 vccd1 _14960_/A sky130_fd_sc_hd__a21o_1
XFILLER_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13909_ _14465_/A _14465_/B _13975_/D vssd1 vssd1 vccd1 vccd1 _13909_/Y sky130_fd_sc_hd__nand3_1
XFILLER_78_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17677_ _17678_/B _17678_/C _17678_/D _17678_/A vssd1 vssd1 vccd1 vccd1 _17679_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14889_ _14889_/A _15006_/B _15005_/B _14889_/D vssd1 vssd1 vccd1 vccd1 _14955_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12378__A _12378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19416_ _19556_/A vssd1 vssd1 vccd1 vccd1 _19555_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16628_ _15616_/X _15657_/Y _15658_/Y vssd1 vssd1 vccd1 vccd1 _16628_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13225__A1 _21383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16962__A2 _16758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19347_ _18795_/X _18814_/X _19455_/A _19346_/Y vssd1 vssd1 vccd1 vccd1 _19374_/A
+ sky130_fd_sc_hd__o211ai_2
X_16559_ _15797_/X _15378_/A _16554_/A vssd1 vssd1 vccd1 vccd1 _16561_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12433__C1 _16318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18164__A1 _12173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19361__B1 _19350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19278_ _19268_/Y _19271_/Y _19274_/Y _19295_/B vssd1 vssd1 vccd1 vccd1 _19284_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__17911__A1 _17226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20510__A3 _17401_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18229_ _18228_/Y _12230_/C _12231_/A vssd1 vssd1 vccd1 vccd1 _18229_/X sky130_fd_sc_hd__a21o_1
XFILLER_164_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19113__B1 _19983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21240_ _21240_/A _21247_/B _21247_/C vssd1 vssd1 vccd1 vccd1 _21243_/A sky130_fd_sc_hd__nand3_1
XFILLER_191_658 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16478__A1 _15455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18512__B _18512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17675__B1 _16016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21171_ _13434_/X _13364_/Y _13385_/B vssd1 vssd1 vccd1 vccd1 _21245_/A sky130_fd_sc_hd__o21a_1
XFILLER_117_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16313__A _20092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20122_ _20154_/A _20154_/B vssd1 vssd1 vccd1 vccd1 _20147_/A sky130_fd_sc_hd__nand2_1
XFILLER_172_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17128__B _17128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19046__D _19689_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20053_ _20032_/B _20042_/Y _20044_/Y _20025_/X _22928_/Q vssd1 vssd1 vccd1 vccd1
+ _20055_/A sky130_fd_sc_hd__a311oi_1
XANTENNA__19624__A _19624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater140 _22761_/CLK vssd1 vssd1 vccd1 vccd1 _22757_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15453__A2 _15450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater151 _22772_/CLK vssd1 vssd1 vccd1 vccd1 _22804_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_27_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17144__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater162 _22738_/CLK vssd1 vssd1 vccd1 vccd1 _22771_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater173 input33/X vssd1 vssd1 vccd1 vccd1 _22725_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20955_ _20906_/Y _21037_/D _21007_/B vssd1 vssd1 vccd1 vccd1 _20958_/A sky130_fd_sc_hd__a21o_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__A2 _15888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20887_/C _20887_/B _20887_/A vssd1 vssd1 vccd1 vccd1 _20894_/C sky130_fd_sc_hd__o21ai_1
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20936__C _20936_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22625_ _22625_/A vssd1 vssd1 vccd1 vccd1 _22800_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14964__A1 _13737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22836__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22556_ _22770_/Q input44/X _22558_/S vssd1 vssd1 vccd1 vccd1 _22557_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21507_ _21658_/A _21658_/B _21658_/C vssd1 vssd1 vccd1 vccd1 _21507_/Y sky130_fd_sc_hd__nand3_2
XFILLER_182_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15913__B1 _16011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22487_ _22487_/A vssd1 vssd1 vccd1 vccd1 _22739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12240_ _12240_/A _12240_/B vssd1 vssd1 vccd1 vccd1 _12241_/B sky130_fd_sc_hd__nor2_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21438_ _21438_/A vssd1 vssd1 vccd1 vccd1 _22931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12171_ _12171_/A vssd1 vssd1 vccd1 vccd1 _12171_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17319__A _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21369_ _21369_/A _21369_/B _21369_/C _21369_/D vssd1 vssd1 vccd1 vccd1 _21374_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17130__A2 _17634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15930_ _15883_/A _15875_/A _15883_/B vssd1 vssd1 vccd1 vccd1 _15930_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15692__A2 _12930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15861_ _15861_/A _15861_/B _15861_/C vssd1 vssd1 vccd1 vccd1 _15864_/C sky130_fd_sc_hd__nand3_1
XFILLER_49_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _17600_/A _17600_/B _17600_/C vssd1 vssd1 vccd1 vccd1 _17781_/B sky130_fd_sc_hd__or3_2
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14812_ _14624_/A _14619_/X _14808_/Y _14809_/Y vssd1 vssd1 vccd1 vccd1 _14813_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _18442_/C _18572_/X _18761_/A _18575_/B _18571_/D vssd1 vssd1 vccd1 vccd1
+ _18582_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _15792_/A _15792_/B _15792_/C vssd1 vssd1 vccd1 vccd1 _15792_/X sky130_fd_sc_hd__or3_1
XFILLER_149_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17531_ _19772_/D _17531_/B _17833_/A _17531_/D vssd1 vssd1 vccd1 vccd1 _17531_/X
+ sky130_fd_sc_hd__and4_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14743_ _14745_/A _14741_/Y _14747_/A vssd1 vssd1 vccd1 vccd1 _14743_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _11285_/A _11285_/B _11633_/A vssd1 vssd1 vccd1 vccd1 _11956_/C sky130_fd_sc_hd__a21oi_1
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17462_ _17462_/A vssd1 vssd1 vccd1 vccd1 _21011_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_189_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14674_ _14622_/X _14636_/D _14672_/X _14057_/X _14560_/A vssd1 vssd1 vccd1 vccd1
+ _14674_/X sky130_fd_sc_hd__a311o_1
XFILLER_33_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15005__C _15006_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11886_ _11896_/C _11886_/B _11886_/C vssd1 vssd1 vccd1 vccd1 _11909_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__16944__A2 _15326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19201_ _19201_/A _19201_/B _19201_/C vssd1 vssd1 vccd1 vccd1 _19208_/A sky130_fd_sc_hd__nand3_2
X_16413_ _16035_/C _16408_/Y _16211_/Y _16204_/Y vssd1 vssd1 vccd1 vccd1 _16686_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__22478__A0 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13625_ _13625_/A vssd1 vssd1 vccd1 vccd1 _13647_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17393_ _17403_/A vssd1 vssd1 vccd1 vccd1 _17393_/X sky130_fd_sc_hd__buf_4
XFILLER_60_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19132_ _19132_/A _19132_/B _19132_/C vssd1 vssd1 vccd1 vccd1 _19132_/Y sky130_fd_sc_hd__nand3_1
X_16344_ _16344_/A vssd1 vssd1 vccd1 vccd1 _20793_/D sky130_fd_sc_hd__clkbuf_2
X_13556_ _13556_/A _13556_/B _13556_/C vssd1 vssd1 vccd1 vccd1 _13558_/B sky130_fd_sc_hd__nand3_1
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19063_ _19063_/A _19063_/B _19063_/C vssd1 vssd1 vccd1 vccd1 _19074_/B sky130_fd_sc_hd__nand3_4
XANTENNA__14707__A1 _14494_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ _12484_/Y _12487_/X _12506_/Y _12432_/B vssd1 vssd1 vccd1 vccd1 _12508_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_160_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16275_ _16275_/A vssd1 vssd1 vccd1 vccd1 _17434_/A sky130_fd_sc_hd__buf_4
XFILLER_185_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13487_ _13487_/A vssd1 vssd1 vccd1 vccd1 _13601_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18014_ _18053_/C _18015_/C _18015_/A vssd1 vssd1 vccd1 vccd1 _18014_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_172_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15226_ _15242_/A _15223_/Y _15225_/Y vssd1 vssd1 vccd1 vccd1 _15227_/B sky130_fd_sc_hd__o21ba_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12438_ _12904_/A vssd1 vssd1 vccd1 vccd1 _20130_/B sky130_fd_sc_hd__buf_2
XANTENNA__18332__B _18691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21453__A1 _21767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15157_ _15188_/A _15185_/B _15154_/X _15155_/X vssd1 vssd1 vccd1 vccd1 _15157_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12661__A _15810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12369_ _12369_/A _12378_/C vssd1 vssd1 vccd1 vccd1 _16293_/A sky130_fd_sc_hd__nand2_2
XFILLER_141_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14108_ _14808_/B vssd1 vssd1 vccd1 vccd1 _15010_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_141_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19965_ _19965_/A _19965_/B vssd1 vssd1 vccd1 vccd1 _19977_/A sky130_fd_sc_hd__nand2_1
X_15088_ _15088_/A _15088_/B vssd1 vssd1 vccd1 vccd1 _15089_/B sky130_fd_sc_hd__and2_1
XFILLER_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22402__A0 _22702_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18916_ _18916_/A _18916_/B vssd1 vssd1 vccd1 vccd1 _18916_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14039_ _14039_/A vssd1 vssd1 vccd1 vccd1 _14099_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_141_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19896_ _19896_/A _19896_/B _19945_/C _19985_/C vssd1 vssd1 vccd1 vccd1 _19937_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18847_ _11702_/X _12010_/A _19014_/A vssd1 vssd1 vccd1 vccd1 _18850_/A sky130_fd_sc_hd__o21ai_1
XFILLER_41_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18778_ _18778_/A _18778_/B _19983_/A _18778_/D vssd1 vssd1 vccd1 vccd1 _18779_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_55_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17729_ _17806_/D _11672_/X _11666_/X _17442_/X _17922_/A vssd1 vssd1 vccd1 vccd1
+ _17736_/A sky130_fd_sc_hd__a311o_1
XFILLER_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22859__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20740_ _20778_/A _20778_/B _20812_/A vssd1 vssd1 vccd1 vccd1 _20740_/Y sky130_fd_sc_hd__nand3_1
XFILLER_24_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20671_ _15940_/A _20611_/Y _20606_/Y vssd1 vssd1 vccd1 vccd1 _20671_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13749__A2 _13746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22410_ _22410_/A vssd1 vssd1 vccd1 vccd1 _22705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16699__A1 _16685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22341_ _22341_/A _22341_/B _22341_/C vssd1 vssd1 vccd1 vccd1 _22341_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__19619__A _19792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22272_ _22309_/A _22272_/B _22272_/C vssd1 vssd1 vccd1 vccd1 _22314_/A sky130_fd_sc_hd__and3_1
XFILLER_117_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17648__B1 _17817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20247__A2 _15325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21223_ _21238_/C _21238_/B _21219_/X _21222_/X vssd1 vssd1 vccd1 vccd1 _21230_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_89_1081 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17139__A _17139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12571__A _12571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21154_ _21154_/A _21154_/B vssd1 vssd1 vccd1 vccd1 _22926_/D sky130_fd_sc_hd__xor2_1
XANTENNA__18860__A2 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20105_ _12803_/X _20214_/A _20471_/C _20090_/Y _16304_/A vssd1 vssd1 vccd1 vccd1
+ _20107_/B sky130_fd_sc_hd__o2111ai_4
XANTENNA__18896__C _18896_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21085_ _21086_/C _17839_/B _17839_/C _21086_/A _21086_/B vssd1 vssd1 vccd1 vccd1
+ _21087_/A sky130_fd_sc_hd__a32o_1
X_20036_ _20035_/A _20058_/C _20033_/A vssd1 vssd1 vccd1 vccd1 _20049_/A sky130_fd_sc_hd__a21oi_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18612__A2 _12171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19504__D _19504_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14929__C _14929_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20012__B _20012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21987_ _21987_/A vssd1 vssd1 vccd1 vccd1 _21987_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11736_/Y _11739_/Y _11935_/C _11708_/Y vssd1 vssd1 vccd1 vccd1 _11755_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22865__D _22877_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _20924_/X _20980_/A _20938_/C vssd1 vssd1 vccd1 vccd1 _20938_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_187_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ _16257_/B vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__buf_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20869_ _20869_/A _20869_/B _20869_/C _20869_/D vssd1 vssd1 vccd1 vccd1 _20879_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ _13664_/D vssd1 vssd1 vccd1 vccd1 _21299_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21668__D1 _21990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22608_ _12107_/C input66/X _22608_/S vssd1 vssd1 vccd1 vccd1 _22609_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17040__C _17040_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14390_ _22769_/Q _14330_/X _14379_/X _22737_/Q _14389_/X vssd1 vssd1 vccd1 vccd1
+ _14390_/X sky130_fd_sc_hd__a221o_1
XFILLER_168_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22654__S _22656_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12465__B _20207_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13341_ _13223_/Y _13225_/X _13286_/B vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__o21a_1
XFILLER_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22539_ _13973_/B input36/X _22547_/S vssd1 vssd1 vccd1 vccd1 _22540_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16060_ _16060_/A vssd1 vssd1 vccd1 vccd1 _16177_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15776__B _15776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ _13272_/A _13272_/B vssd1 vssd1 vccd1 vccd1 _13272_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_input76_A x[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12176__A1 _12173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15268__S _15268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15011_ _15007_/Y _15010_/Y _15008_/X vssd1 vssd1 vccd1 vccd1 _15080_/B sky130_fd_sc_hd__a21oi_1
XFILLER_120_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12223_ _12225_/A _18228_/B _18227_/C vssd1 vssd1 vccd1 vccd1 _12227_/A sky130_fd_sc_hd__a21o_1
XFILLER_68_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18300__A1 _18305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12912__C _16067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16311__B1 _15938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ _19016_/B _19016_/C _12154_/C vssd1 vssd1 vccd1 vccd1 _12154_/Y sky130_fd_sc_hd__nand3_1
XFILLER_29_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11809__B _11809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15792__A _15792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19750_ _19750_/A vssd1 vssd1 vccd1 vccd1 _19750_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16103__D _16103_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16962_ _16179_/A _16758_/X _16959_/A vssd1 vssd1 vccd1 vccd1 _16967_/A sky130_fd_sc_hd__o21ai_1
X_12085_ _12054_/X _12056_/Y _12039_/Y _12081_/Y vssd1 vssd1 vccd1 vccd1 _12086_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_96_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11528__C _12003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14873__B1 _14575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18701_ _18705_/A _18487_/B _18340_/B _18482_/Y vssd1 vssd1 vccd1 vccd1 _18702_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_15913_ _15924_/A _15924_/B _15924_/C _16011_/A _16011_/B vssd1 vssd1 vccd1 vccd1
+ _15913_/Y sky130_fd_sc_hd__a32oi_4
X_19681_ _19681_/A _19681_/B _19681_/C vssd1 vssd1 vccd1 vccd1 _19761_/A sky130_fd_sc_hd__and3_1
X_16893_ _16890_/X _16672_/A _16889_/C vssd1 vssd1 vccd1 vccd1 _17215_/B sky130_fd_sc_hd__o21ai_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16400__B _21050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18632_ _12204_/X _17400_/X _18626_/Y _18629_/Y _18953_/A vssd1 vssd1 vccd1 vccd1
+ _18633_/B sky130_fd_sc_hd__o311ai_1
X_15844_ _15756_/X _15750_/Y _15864_/B _15854_/A vssd1 vssd1 vccd1 vccd1 _15844_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__20410__A2 _20381_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14625__B1 _15188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18563_ _18565_/A _18765_/B _18568_/B _18568_/C vssd1 vssd1 vccd1 vccd1 _18564_/C
+ sky130_fd_sc_hd__a22o_1
X_15775_ _16191_/A _15775_/B _15775_/C _17085_/C vssd1 vssd1 vccd1 vccd1 _15783_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _20452_/A _20452_/B _12711_/X _20793_/A _16153_/A vssd1 vssd1 vccd1 vccd1
+ _12990_/B sky130_fd_sc_hd__a32o_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12100__A1 _11381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17514_ _17514_/A _17600_/A vssd1 vssd1 vccd1 vccd1 _17514_/Y sky130_fd_sc_hd__nand2_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14729_/A _14729_/B _14726_/C _14726_/D vssd1 vssd1 vccd1 vccd1 _14731_/B
+ sky130_fd_sc_hd__nand4_1
X_11938_ _11938_/A _11938_/B vssd1 vssd1 vccd1 vccd1 _11938_/Y sky130_fd_sc_hd__nand2_2
X_18494_ _11541_/X _19624_/A _18487_/A vssd1 vssd1 vccd1 vccd1 _18499_/A sky130_fd_sc_hd__o21ai_1
XFILLER_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16917__A2 _17443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _17442_/X _17731_/A _16016_/X _17439_/X vssd1 vssd1 vccd1 vccd1 _17445_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14657_ _14561_/D _14561_/Y _14655_/Y _14752_/A vssd1 vssd1 vccd1 vccd1 _14758_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_11869_ _11308_/A _11308_/B _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11869_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12939__B1 _15696_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ _13608_/A _13608_/B _13608_/C vssd1 vssd1 vccd1 vccd1 _13617_/A sky130_fd_sc_hd__nand3_1
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17376_ _17060_/B _17229_/Y _17353_/X vssd1 vssd1 vccd1 vccd1 _17376_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14588_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14729_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19115_ _19122_/A _19122_/B _19122_/C _19114_/X vssd1 vssd1 vccd1 vccd1 _19121_/A
+ sky130_fd_sc_hd__a31oi_2
X_16327_ _15645_/X _16332_/B _16996_/A _16062_/A vssd1 vssd1 vccd1 vccd1 _16327_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15338__D1 _16809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13539_ _13539_/A vssd1 vssd1 vccd1 vccd1 _13614_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_145_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21688__B _21688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20331__D1 _20129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12094__C _19358_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19046_ _19046_/A _19065_/A _19046_/C _19689_/C vssd1 vssd1 vccd1 vccd1 _19046_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_174_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16258_ _16059_/A _16274_/A _16257_/Y vssd1 vssd1 vccd1 vccd1 _16258_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__16550__B1 _11779_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15209_ _15209_/A _15209_/B vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__nor2_2
XFILLER_126_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16189_ _16043_/C _16090_/Y _16188_/Y vssd1 vssd1 vccd1 vccd1 _16190_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12391__A _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16838__D1 _16452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18842__A2 _18678_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15656__A2 _15630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19948_ _19948_/A _19948_/B vssd1 vssd1 vccd1 vccd1 _19949_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14864__B1 _14366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19879_ _19293_/X _19294_/X _19820_/Y _19761_/Y _19878_/Y vssd1 vssd1 vccd1 vccd1
+ _19885_/B sky130_fd_sc_hd__o221ai_2
XFILLER_96_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_995 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11735__A _15559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22681__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21910_ _21909_/Y _21906_/A _21913_/A _21913_/B vssd1 vssd1 vccd1 vccd1 _21911_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22890_ _22952_/CLK _22890_/D vssd1 vssd1 vccd1 vccd1 _22890_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15813__C1 _11506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21841_ _21841_/A _21841_/B _21841_/C vssd1 vssd1 vccd1 vccd1 _21841_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__18358__A1 _18156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17422__A _17422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21772_ _21846_/B _21846_/C _21770_/Y _21771_/X vssd1 vssd1 vccd1 vccd1 _21778_/D
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_130_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20486__C _20486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17141__B _17532_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20723_ _20723_/A vssd1 vssd1 vccd1 vccd1 _20806_/B sky130_fd_sc_hd__buf_2
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20654_ _20650_/A _20650_/B _20648_/A vssd1 vssd1 vccd1 vccd1 _20656_/B sky130_fd_sc_hd__a21o_1
XFILLER_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20468__A2 _16708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20585_ _20464_/B _20697_/B _20695_/A _20584_/Y vssd1 vssd1 vccd1 vccd1 _20586_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_165_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18530__A1 _18156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22324_ _22324_/A _22324_/B vssd1 vssd1 vccd1 vccd1 _22325_/C sky130_fd_sc_hd__nor2_1
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22255_ _22080_/B _22163_/Y _22140_/A _22140_/B vssd1 vssd1 vccd1 vccd1 _22255_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21206_ _21201_/Y _21202_/Y _21203_/X vssd1 vssd1 vccd1 vccd1 _21210_/A sky130_fd_sc_hd__o21ai_1
XFILLER_132_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22186_ _22186_/A _22186_/B vssd1 vssd1 vccd1 vccd1 _22186_/X sky130_fd_sc_hd__or2_1
XANTENNA__18833__A2 _18619_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_918 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21137_ _21138_/A _21138_/B _21138_/C vssd1 vssd1 vccd1 vccd1 _21137_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_132_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14855__B1 _13904_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11669__B1 _11667_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21068_ _21068_/A _21068_/B vssd1 vssd1 vccd1 vccd1 _21079_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_962 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20019_ _19995_/A _19995_/B _19992_/C _19992_/B vssd1 vssd1 vccd1 vccd1 _20020_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_12910_ _20481_/C vssd1 vssd1 vccd1 vccd1 _20593_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13890_ _13881_/Y _13887_/X _13888_/Y _13889_/Y vssd1 vssd1 vccd1 vccd1 _13891_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_104_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_bq_clk_i clkbuf_2_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_73_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12841_ _20255_/B _12921_/A _12718_/X _16300_/A _20142_/A vssd1 vssd1 vccd1 vccd1
+ _12855_/B sky130_fd_sc_hd__o221ai_4
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15472_/X _15557_/Y _15558_/Y _15559_/Y vssd1 vssd1 vccd1 vccd1 _15568_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12772_/A vssd1 vssd1 vccd1 vccd1 _12772_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _15008_/C _14834_/C _14834_/A _14512_/B _14512_/C vssd1 vssd1 vccd1 vccd1
+ _14515_/B sky130_fd_sc_hd__a32o_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _16447_/A vssd1 vssd1 vccd1 vccd1 _19320_/A sky130_fd_sc_hd__buf_2
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _12209_/A _12211_/A _15586_/C _17234_/A vssd1 vssd1 vccd1 vccd1 _15498_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_9_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_564 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17058_/A _17058_/B _17229_/Y vssd1 vssd1 vccd1 vccd1 _17230_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__11380__A _11380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _22662_/A vssd1 vssd1 vccd1 vccd1 _22658_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12907__C _15804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11654_ _12210_/A vssd1 vssd1 vccd1 vccd1 _16242_/A sky130_fd_sc_hd__buf_2
XFILLER_120_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14386__A2 _14370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17161_ _17181_/A _17181_/B _17161_/C vssd1 vssd1 vccd1 vccd1 _17173_/C sky130_fd_sc_hd__nand3_1
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14373_ _18698_/A _14354_/X _14355_/X _14361_/X _22765_/Q vssd1 vssd1 vccd1 vccd1
+ _14373_/X sky130_fd_sc_hd__a32o_1
X_11585_ _11585_/A vssd1 vssd1 vccd1 vccd1 _18156_/A sky130_fd_sc_hd__buf_2
XFILLER_156_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16112_ _15901_/A _15901_/B _12913_/A _16106_/D _16554_/C vssd1 vssd1 vccd1 vccd1
+ _16113_/B sky130_fd_sc_hd__a32o_1
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13324_ _13324_/A _13324_/B vssd1 vssd1 vccd1 vccd1 _13324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17092_ _15888_/X _17435_/A _17591_/B vssd1 vssd1 vccd1 vccd1 _17520_/A sky130_fd_sc_hd__o21ai_4
XFILLER_10_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13346__B1 _13326_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16043_ _16043_/A _16043_/B _16043_/C vssd1 vssd1 vccd1 vccd1 _16414_/C sky130_fd_sc_hd__nand3_1
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13255_ _13623_/A vssd1 vssd1 vccd1 vccd1 _13401_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater130_A _22870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12206_ _15838_/A vssd1 vssd1 vccd1 vccd1 _16940_/A sky130_fd_sc_hd__buf_2
XANTENNA__18285__B1 _15530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13186_ _13430_/A vssd1 vssd1 vccd1 vccd1 _13581_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19802_ _19864_/A _19864_/B _19866_/A _19865_/B vssd1 vssd1 vccd1 vccd1 _19804_/B
+ sky130_fd_sc_hd__nand4_1
X_12137_ _12137_/A _12137_/B vssd1 vssd1 vccd1 vccd1 _12138_/C sky130_fd_sc_hd__nand2_1
XFILLER_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17994_ _17994_/A _17994_/B vssd1 vssd1 vccd1 vccd1 _17996_/A sky130_fd_sc_hd__or2_2
XFILLER_150_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14846__B1 _14845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19733_ _19728_/Y _19731_/Y _19736_/C vssd1 vssd1 vccd1 vccd1 _19742_/B sky130_fd_sc_hd__o21bai_1
X_16945_ _16940_/X _15723_/X _16941_/X _16944_/Y _16934_/A vssd1 vssd1 vccd1 vccd1
+ _16945_/X sky130_fd_sc_hd__o221a_1
X_12068_ _18810_/D vssd1 vssd1 vccd1 vccd1 _19046_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__18588__A1 _19443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16130__B _16130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__A _22957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19664_ _19664_/A _19664_/B _19664_/C vssd1 vssd1 vccd1 vccd1 _19813_/A sky130_fd_sc_hd__nand3_2
X_16876_ _17006_/A vssd1 vssd1 vccd1 vccd1 _20972_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18615_ _18810_/A _19353_/B _19353_/C vssd1 vssd1 vccd1 vccd1 _18616_/B sky130_fd_sc_hd__and3_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _15784_/Y _15803_/Y _15828_/A _15826_/Y vssd1 vssd1 vccd1 vccd1 _15853_/B
+ sky130_fd_sc_hd__o211a_2
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19595_ _19596_/B _19596_/C _19176_/X _17730_/A vssd1 vssd1 vccd1 vccd1 _19684_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_18_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15758_ _15758_/A _15758_/B _15758_/C vssd1 vssd1 vccd1 vccd1 _15864_/D sky130_fd_sc_hd__nand3_2
X_18546_ _18553_/A _18553_/B _18546_/C vssd1 vssd1 vccd1 vccd1 _18548_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19001__A2 _18986_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17012__A1 _16732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14709_ _14711_/C _14711_/D vssd1 vssd1 vccd1 vccd1 _14716_/C sky130_fd_sc_hd__nand2_1
XFILLER_178_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18477_ _18765_/A _18478_/B _18478_/C vssd1 vssd1 vccd1 vccd1 _18565_/A sky130_fd_sc_hd__a21o_1
X_15689_ _12968_/B _16921_/A _12719_/A _12118_/A vssd1 vssd1 vccd1 vccd1 _15693_/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11290__A _22955_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17428_ _14432_/A _15808_/X _11672_/X _20854_/A _20854_/B vssd1 vssd1 vccd1 vccd1
+ _17564_/A sky130_fd_sc_hd__o2111ai_4
XANTENNA__11721__C _11721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12388__A1 _16318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17359_ _16672_/X _16673_/Y _16892_/B _16892_/C vssd1 vssd1 vccd1 vccd1 _17361_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20370_ _20511_/A _20593_/D _20608_/A _20370_/D vssd1 vssd1 vccd1 vccd1 _20371_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_174_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19029_ _19029_/A vssd1 vssd1 vccd1 vccd1 _19037_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22040_ _22041_/A _22106_/A _22041_/C vssd1 vssd1 vccd1 vccd1 _22040_/Y sky130_fd_sc_hd__nand3_1
XFILLER_86_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18815__A2 _12204_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16826__A1 _16451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11465__A _15776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22942_ _22943_/CLK _22942_/D vssd1 vssd1 vccd1 vccd1 _22942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19351__B _19351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22873_ _22915_/CLK _22873_/D vssd1 vssd1 vccd1 vccd1 _22873_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21824_ _21930_/A _21834_/A _21822_/Y _21823_/Y vssd1 vssd1 vccd1 vccd1 _21825_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_93_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17003__A1 _16098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14495__B _14611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21755_ _21579_/A _14380_/A _22734_/Q vssd1 vssd1 vccd1 vccd1 _21755_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20706_ _17423_/X _17424_/X _20210_/B _12928_/X vssd1 vssd1 vccd1 vccd1 _20706_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21686_ _21686_/A vssd1 vssd1 vccd1 vccd1 _21814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20637_ _20637_/A vssd1 vssd1 vccd1 vccd1 _20734_/C sky130_fd_sc_hd__buf_2
XFILLER_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14942__C _14942_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20846__C1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ _11796_/A vssd1 vssd1 vccd1 vccd1 _15357_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__20310__A1 _20553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20568_ _20568_/A _20568_/B vssd1 vssd1 vccd1 vccd1 _20568_/X sky130_fd_sc_hd__and2_1
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22307_ _22307_/A _22307_/B vssd1 vssd1 vccd1 vccd1 _22309_/B sky130_fd_sc_hd__nand2_1
XFILLER_166_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20499_ _20499_/A _20499_/B _20629_/A _20499_/D vssd1 vssd1 vccd1 vccd1 _20500_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_180_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13040_ _13040_/A _13040_/B _13040_/C vssd1 vssd1 vccd1 vccd1 _13045_/B sky130_fd_sc_hd__nand3_4
XFILLER_180_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22238_ _22238_/A _22238_/B vssd1 vssd1 vccd1 vccd1 _22240_/A sky130_fd_sc_hd__nand2_1
XFILLER_191_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18806__A2 _16799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22233__A _22233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12551__A1 _12669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22169_ _22168_/X _22102_/Y _22102_/B vssd1 vssd1 vccd1 vccd1 _22195_/A sky130_fd_sc_hd__o21ai_2
XFILLER_120_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19180__A2_N _19015_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input39_A wb_dat_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ _14990_/X _14494_/D _14969_/B _14968_/B vssd1 vssd1 vccd1 vccd1 _15034_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_94_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19767__B1 _17817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13942_ _14770_/A _14771_/A _14210_/A _13978_/A _14489_/C vssd1 vssd1 vccd1 vccd1
+ _13942_/Y sky130_fd_sc_hd__a32oi_4
X_16730_ _20584_/B vssd1 vssd1 vccd1 vccd1 _20792_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20688__A _20793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ _16664_/C _16426_/X _16664_/B _17502_/A _16660_/Y vssd1 vssd1 vccd1 vccd1
+ _16702_/B sky130_fd_sc_hd__a311o_1
XFILLER_47_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15789__D1 _15960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13873_ _13873_/A vssd1 vssd1 vccd1 vccd1 _13873_/X sky130_fd_sc_hd__buf_2
XFILLER_62_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18400_ _18308_/Y _18309_/X _18394_/Y _18399_/Y vssd1 vssd1 vccd1 vccd1 _18411_/B
+ sky130_fd_sc_hd__o22ai_2
X_15612_ _16611_/A vssd1 vssd1 vccd1 vccd1 _16737_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12067__B1 _18305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ _12824_/A _16320_/A vssd1 vssd1 vccd1 vccd1 _15617_/A sky130_fd_sc_hd__nor2_4
X_19380_ _19372_/X _19377_/Y _19378_/Y _19379_/Y vssd1 vssd1 vccd1 vccd1 _19389_/B
+ sky130_fd_sc_hd__o211ai_4
X_16592_ _15936_/A _16745_/A _16332_/B _16590_/X _16570_/A vssd1 vssd1 vccd1 vccd1
+ _16598_/B sky130_fd_sc_hd__o311a_2
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15543_ _15532_/X _16215_/A _15542_/X vssd1 vssd1 vccd1 vccd1 _15543_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18331_ _16241_/A _11988_/X _15901_/A _19322_/B _19322_/C vssd1 vssd1 vccd1 vccd1
+ _18980_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12755_ _12755_/A _12755_/B _12755_/C vssd1 vssd1 vccd1 vccd1 _12755_/X sky130_fd_sc_hd__and3_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18262_ _18257_/B _18598_/B _18257_/Y _18261_/X vssd1 vssd1 vccd1 vccd1 _18262_/Y
+ sky130_fd_sc_hd__o211ai_1
X_11706_ _11706_/A vssd1 vssd1 vccd1 vccd1 _11707_/A sky130_fd_sc_hd__buf_2
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15556__A1 _15838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15474_ _15474_/A _15474_/B _15474_/C vssd1 vssd1 vccd1 vccd1 _15501_/A sky130_fd_sc_hd__nand3_1
XFILLER_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15556__B2 _15498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _22817_/Q vssd1 vssd1 vccd1 vccd1 _20357_/B sky130_fd_sc_hd__buf_2
XFILLER_187_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17213_ _17518_/C _17213_/B _17213_/C vssd1 vssd1 vccd1 vccd1 _17370_/B sky130_fd_sc_hd__nand3_2
X_14425_ _22814_/Q _14354_/A _14355_/A _14361_/A _22782_/Q vssd1 vssd1 vccd1 vccd1
+ _14425_/X sky130_fd_sc_hd__a32o_1
X_18193_ _18193_/A vssd1 vssd1 vccd1 vccd1 _19353_/C sky130_fd_sc_hd__clkbuf_2
X_11637_ _18328_/B _18328_/C vssd1 vssd1 vccd1 vccd1 _18330_/A sky130_fd_sc_hd__nand2_2
XFILLER_24_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12934__A _15988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17144_ _17144_/A _17401_/C _17144_/C vssd1 vssd1 vccd1 vccd1 _17145_/B sky130_fd_sc_hd__nand3_2
XFILLER_128_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14356_ _18127_/B _14354_/X _14355_/X _14334_/X _13973_/B vssd1 vssd1 vccd1 vccd1
+ _14356_/X sky130_fd_sc_hd__a32o_1
XFILLER_196_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11568_ _11568_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _15476_/A sky130_fd_sc_hd__nand2_1
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20640__A1_N _20631_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ _13311_/C vssd1 vssd1 vccd1 vccd1 _21495_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_196_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17075_ _17049_/A _17049_/B _16886_/B vssd1 vssd1 vccd1 vccd1 _17077_/A sky130_fd_sc_hd__a21oi_1
XFILLER_116_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20852__A2 _17444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14287_ _14250_/A _14250_/B _14250_/C _14253_/Y _14243_/A vssd1 vssd1 vccd1 vccd1
+ _14288_/C sky130_fd_sc_hd__a32o_1
X_11499_ _12154_/C vssd1 vssd1 vccd1 vccd1 _18507_/C sky130_fd_sc_hd__buf_2
XANTENNA__20870__B _20870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16026_ _16026_/A vssd1 vssd1 vccd1 vccd1 _16026_/Y sky130_fd_sc_hd__inv_2
X_13238_ _22722_/Q vssd1 vssd1 vccd1 vccd1 _13240_/A sky130_fd_sc_hd__inv_2
XANTENNA__20065__B1 _13041_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__A1 _20210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16808__A1 _16275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17237__A _20608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ _13147_/A _13147_/B _13176_/A vssd1 vssd1 vccd1 vccd1 _13169_/X sky130_fd_sc_hd__a21o_1
XFILLER_151_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16498__D _16498_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17977_ _21050_/D _17882_/A _18028_/A _17932_/B _17932_/A vssd1 vssd1 vccd1 vccd1
+ _17988_/A sky130_fd_sc_hd__a32o_1
XFILLER_111_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11285__A _11285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19716_ _19621_/B _19621_/Y _19715_/X vssd1 vssd1 vccd1 vccd1 _19788_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__14299__C input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16928_ _16015_/A _15940_/A _16815_/Y _16810_/D vssd1 vssd1 vccd1 vccd1 _16930_/C
+ sky130_fd_sc_hd__o31a_2
XFILLER_78_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18025__A3 _21048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19647_ _19641_/X _19643_/Y _19649_/B vssd1 vssd1 vccd1 vccd1 _19650_/C sky130_fd_sc_hd__o21bai_1
XFILLER_66_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16859_ _16860_/A _16860_/B _16860_/C _16869_/B vssd1 vssd1 vccd1 vccd1 _16859_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22109__A2 _21594_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19602__D _19769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12058__B1 _11897_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19578_ _19561_/A _19561_/B _19663_/B vssd1 vssd1 vccd1 vccd1 _19682_/B sky130_fd_sc_hd__a21o_1
XFILLER_164_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15795__A1 _12606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20110__B _20110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18529_ _18529_/A _18529_/B vssd1 vssd1 vccd1 vccd1 _18529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18194__C1 _18200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13650__D _21195_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15547__A1 _15545_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21540_ _21537_/Y _21538_/Y _21531_/C _21539_/Y vssd1 vssd1 vccd1 vccd1 _21540_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_194_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16744__B1 _16732_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15547__B2 _15524_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20540__A1 _20843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_2_0_bq_clk_i_A clkbuf_2_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11744__A2_N _11905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21471_ _21476_/A vssd1 vssd1 vccd1 vccd1 _21876_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12844__A _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20422_ _20423_/A _20423_/B _20423_/C vssd1 vssd1 vccd1 vccd1 _20422_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_181_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15577__D _15577_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20353_ _20353_/A _20353_/B _20353_/C vssd1 vssd1 vccd1 vccd1 _20366_/C sky130_fd_sc_hd__nand3_2
XFILLER_134_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20780__B _21019_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20284_ _20284_/A _20284_/B _20284_/C _20452_/C vssd1 vssd1 vccd1 vccd1 _20401_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__19346__B _19504_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22023_ _22011_/X _22013_/B _22013_/A vssd1 vssd1 vccd1 vccd1 _22084_/A sky130_fd_sc_hd__a21boi_2
XANTENNA__16051__A _20745_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15890__A _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17224__A1 _22895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22925_ _22948_/CLK _22925_/D vssd1 vssd1 vccd1 vccd1 _22925_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22856_ _22937_/CLK _22868_/Q vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17313__C _19482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21859__A1 _21964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21807_ _21797_/Y _21913_/A _21806_/X vssd1 vssd1 vccd1 vccd1 _21807_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22787_ _22787_/CLK _22787_/D vssd1 vssd1 vccd1 vccd1 _22787_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17527__A2 _17526_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18706__A _18706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12540_ _20611_/B _12970_/A _12540_/C _15306_/C vssd1 vssd1 vccd1 vccd1 _12540_/X
+ sky130_fd_sc_hd__and4_2
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21738_ _21738_/A vssd1 vssd1 vccd1 vccd1 _22041_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _22688_/Q vssd1 vssd1 vccd1 vccd1 _12520_/A sky130_fd_sc_hd__buf_2
X_21669_ _21651_/X _21665_/Y _21667_/Y vssd1 vssd1 vccd1 vccd1 _21669_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14210_ _14210_/A vssd1 vssd1 vccd1 vccd1 _14779_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11422_ _11428_/B _18319_/C _11418_/A vssd1 vssd1 vccd1 vccd1 _12171_/A sky130_fd_sc_hd__a21boi_4
XFILLER_177_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15190_ _15050_/A _15154_/A _15050_/C _15215_/A _15119_/D vssd1 vssd1 vccd1 vccd1
+ _15190_/X sky130_fd_sc_hd__a32o_1
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16499__C1 _18258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14141_ _14238_/A _14141_/B vssd1 vssd1 vccd1 vccd1 _14151_/A sky130_fd_sc_hd__nand2_1
X_11353_ _11319_/Y _11333_/X _11352_/X vssd1 vssd1 vccd1 vccd1 _11477_/B sky130_fd_sc_hd__a21o_1
XFILLER_165_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14072_ _14085_/A _14085_/B _14071_/Y vssd1 vssd1 vccd1 vccd1 _14072_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14513__A2 _13968_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11284_ _11860_/A _11860_/B _11860_/C vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__nand3_2
XFILLER_4_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17900_ _17900_/A _17900_/B vssd1 vssd1 vccd1 vccd1 _17900_/X sky130_fd_sc_hd__and2_1
XANTENNA__13585__A _21195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ _13018_/X _13019_/Y _20284_/A _13022_/X vssd1 vssd1 vccd1 vccd1 _13028_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16599__C _16599_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18880_ _18880_/A _18880_/B vssd1 vssd1 vccd1 vccd1 _18883_/B sky130_fd_sc_hd__nand2_1
XANTENNA__20598__A1 _20697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17463__A1 _11904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17831_ _17831_/A _17890_/B _17831_/C vssd1 vssd1 vccd1 vccd1 _17897_/A sky130_fd_sc_hd__nand3_2
XANTENNA__17463__B2 _16580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17762_ _17761_/B _17761_/C _17736_/X vssd1 vssd1 vccd1 vccd1 _17765_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__19204__A2 _17400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15008__C _15008_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14974_ _14914_/C _14972_/Y _14970_/X _14971_/Y vssd1 vssd1 vccd1 vccd1 _15035_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_86_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19501_ _19359_/X _19500_/X _19497_/B _19494_/Y vssd1 vssd1 vccd1 vccd1 _19503_/B
+ sky130_fd_sc_hd__o211ai_1
X_16713_ _16710_/Y _16711_/Y _16712_/X vssd1 vssd1 vccd1 vccd1 _16743_/A sky130_fd_sc_hd__a21o_2
X_13925_ _13923_/X _13924_/X _13903_/Y vssd1 vssd1 vccd1 vccd1 _13937_/B sky130_fd_sc_hd__o21ai_1
X_17693_ _17693_/A _17693_/B _17693_/C vssd1 vssd1 vccd1 vccd1 _17701_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12929__A _12929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16569__A3 _17875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19432_ _19147_/A _19299_/Y _19302_/Y vssd1 vssd1 vccd1 vccd1 _19432_/Y sky130_fd_sc_hd__a21oi_2
X_16644_ _16895_/A _16895_/B _16644_/C vssd1 vssd1 vccd1 vccd1 _16644_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__15777__A1 _11504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856_ _13856_/A vssd1 vssd1 vccd1 vccd1 _14571_/A sky130_fd_sc_hd__buf_2
XFILLER_179_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12807_ _12314_/Y _12329_/X _12428_/Y _12334_/A vssd1 vssd1 vccd1 vccd1 _12810_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_19363_ _19357_/Y _19218_/A _19368_/B _19362_/Y vssd1 vssd1 vccd1 vccd1 _19363_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_76_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13787_ _14165_/A _14165_/C vssd1 vssd1 vccd1 vccd1 _14055_/B sky130_fd_sc_hd__nand2_1
X_16575_ _20579_/B vssd1 vssd1 vccd1 vccd1 _20584_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1031 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17520__A _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22892__CLK _22952_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18314_ _11783_/A _18313_/Y _11377_/A vssd1 vssd1 vccd1 vccd1 _18324_/A sky130_fd_sc_hd__o21bai_1
XFILLER_176_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15526_ _12672_/A _16786_/A _15589_/A vssd1 vssd1 vccd1 vccd1 _15527_/A sky130_fd_sc_hd__o21ai_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_692 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12738_ _12933_/B _12933_/C _12933_/D _12710_/Y vssd1 vssd1 vccd1 vccd1 _12739_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_187_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19294_ _19294_/A vssd1 vssd1 vccd1 vccd1 _19294_/X sky130_fd_sc_hd__buf_2
XANTENNA__15959__B _16400_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20584__C _20584_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18245_ _18259_/A _18258_/B vssd1 vssd1 vccd1 vccd1 _18246_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16781__D _18193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15457_ _15457_/A _15457_/B vssd1 vssd1 vccd1 vccd1 _15457_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ _12669_/A vssd1 vssd1 vccd1 vccd1 _12758_/A sky130_fd_sc_hd__inv_2
XFILLER_129_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14201__B2 _14199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14408_ _22808_/Q _14397_/X _14398_/X _14391_/X _22776_/Q vssd1 vssd1 vccd1 vccd1
+ _14408_/X sky130_fd_sc_hd__a32o_1
XFILLER_191_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15388_ _15389_/B _15389_/C _15389_/A vssd1 vssd1 vccd1 vccd1 _15388_/Y sky130_fd_sc_hd__a21oi_1
X_18176_ _18279_/A _18278_/A vssd1 vssd1 vccd1 vccd1 _18184_/A sky130_fd_sc_hd__nand2_1
X_17127_ _17127_/A _17323_/A vssd1 vssd1 vccd1 vccd1 _17178_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14339_ _14355_/A vssd1 vssd1 vccd1 vccd1 _14339_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__20825__A2 _20759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17058_ _17058_/A _17058_/B vssd1 vssd1 vccd1 vccd1 _17213_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14504__A2 _14057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16009_ _16010_/A _16010_/B _16009_/C vssd1 vssd1 vccd1 vccd1 _16009_/Y sky130_fd_sc_hd__nand3_1
XFILLER_98_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20589__A1 _13022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15465__B1 _11667_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20971_ _15355_/A _15355_/B _20967_/Y _20843_/X _20969_/Y vssd1 vssd1 vccd1 vccd1
+ _20982_/B sky130_fd_sc_hd__a2111oi_1
XFILLER_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12839__A _16708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18954__B2 _18627_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22710_ _22743_/CLK _22710_/D vssd1 vssd1 vccd1 vccd1 _22710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15232__A3 _15180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22641_ _22808_/Q input51/X _22641_/S vssd1 vssd1 vccd1 vccd1 _22642_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22572_ _22777_/Q input52/X _22580_/S vssd1 vssd1 vccd1 vccd1 _22573_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12451__B1 _12450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18245__B _18258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21523_ _21665_/D _21522_/A _21522_/C _21522_/B vssd1 vssd1 vccd1 vccd1 _21524_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16193__A1 _16192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21454_ _21454_/A vssd1 vssd1 vccd1 vccd1 _22034_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20405_ _20379_/X _20380_/Y _20403_/X _20404_/Y vssd1 vssd1 vccd1 vccd1 _20405_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_193_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21385_ _21385_/A _21385_/B vssd1 vssd1 vccd1 vccd1 _21386_/C sky130_fd_sc_hd__nand2_1
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_851 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20336_ _20336_/A _20336_/B vssd1 vssd1 vccd1 vccd1 _20337_/A sky130_fd_sc_hd__nor2_2
XFILLER_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19507__D _19507_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20267_ _20264_/A _20390_/D _20260_/A _20234_/A _20397_/B vssd1 vssd1 vccd1 vccd1
+ _20268_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_163_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17445__A1 _17442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22006_ _22008_/C _22008_/D _22005_/Y vssd1 vssd1 vccd1 vccd1 _22013_/A sky130_fd_sc_hd__a21o_1
XFILLER_49_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18642__B1 _18619_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21241__A2 _21247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20198_ _20147_/A _20197_/Y _20150_/B vssd1 vssd1 vccd1 vccd1 _20198_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_163_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14013__B _14013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19737__A3 _19419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _15904_/A _15905_/A _12127_/A _18325_/A vssd1 vssd1 vccd1 vccd1 _11984_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11653__A _15694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13710_ _14203_/B vssd1 vssd1 vccd1 vccd1 _14191_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_72_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22908_ _22968_/CLK _22908_/D vssd1 vssd1 vccd1 vccd1 _22908_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _14681_/X _14682_/X _14687_/X _14689_/Y vssd1 vssd1 vccd1 vccd1 _14716_/A
+ sky130_fd_sc_hd__o22ai_4
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13641_ _13666_/A _13666_/B _13666_/C vssd1 vssd1 vccd1 vccd1 _13641_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22839_ _22850_/CLK _22851_/Q vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_787 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16586_/B _17833_/B _17833_/C _16400_/A _16431_/A vssd1 vssd1 vccd1 vccd1
+ _16360_/X sky130_fd_sc_hd__a32o_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12978__D1 _12930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20504__A1 _15723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ _13572_/A _13572_/B _21866_/C _21938_/B vssd1 vssd1 vccd1 vccd1 _13618_/A
+ sky130_fd_sc_hd__nand4_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15311_ _15302_/B _15306_/Y _15502_/A vssd1 vssd1 vccd1 vccd1 _15461_/A sky130_fd_sc_hd__o21ai_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12523_/A vssd1 vssd1 vccd1 vccd1 _16488_/A sky130_fd_sc_hd__clkbuf_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16291_ _16289_/Y _16290_/X _16282_/A vssd1 vssd1 vccd1 vccd1 _16291_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_9_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18030_ _18030_/A _18030_/B _18030_/C _18030_/D vssd1 vssd1 vccd1 vccd1 _18030_/Y
+ sky130_fd_sc_hd__nand4_1
X_15242_ _15242_/A _15242_/B vssd1 vssd1 vccd1 vccd1 _15243_/B sky130_fd_sc_hd__xnor2_2
X_12454_ _12454_/A _12454_/B _12454_/C vssd1 vssd1 vccd1 vccd1 _12455_/A sky130_fd_sc_hd__nand3_2
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11405_ _16481_/A vssd1 vssd1 vccd1 vccd1 _15482_/A sky130_fd_sc_hd__buf_2
XFILLER_126_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19267__A _19272_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16106__D _16106_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15173_ _15173_/A _15173_/B _15173_/C vssd1 vssd1 vccd1 vccd1 _15174_/B sky130_fd_sc_hd__or3_1
XANTENNA__20807__A2 _15935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12385_ _12385_/A vssd1 vssd1 vccd1 vccd1 _16319_/C sky130_fd_sc_hd__buf_2
XFILLER_153_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14124_ _14576_/A _13905_/Y _13829_/A _14123_/X _14085_/Y vssd1 vssd1 vccd1 vccd1
+ _14128_/B sky130_fd_sc_hd__o221ai_2
XFILLER_67_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11336_ _11411_/A vssd1 vssd1 vccd1 vccd1 _12210_/A sky130_fd_sc_hd__clkbuf_2
X_19981_ _19981_/A vssd1 vssd1 vccd1 vccd1 _19987_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18932_ _18932_/A _18932_/B _18932_/C vssd1 vssd1 vccd1 vccd1 _18932_/Y sky130_fd_sc_hd__nand3_2
XFILLER_97_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14055_ _14165_/B _14055_/B vssd1 vssd1 vccd1 vccd1 _14055_/X sky130_fd_sc_hd__and2_1
XFILLER_140_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13006_ _13006_/A _13006_/B vssd1 vssd1 vccd1 vccd1 _13039_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18863_ _18863_/A _18869_/D _18869_/A _19091_/B vssd1 vssd1 vccd1 vccd1 _18863_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_79_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17814_ _19769_/B vssd1 vssd1 vccd1 vccd1 _19842_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_39_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18794_ _18748_/B _18737_/X _18743_/A vssd1 vssd1 vccd1 vccd1 _18938_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__15998__B2 _15983_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20579__C _20579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17745_ _17386_/B _20675_/B _18305_/C _17826_/A _17743_/D vssd1 vssd1 vccd1 vccd1
+ _17745_/X sky130_fd_sc_hd__a32o_1
XANTENNA__13762__B _13949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14957_ _14952_/Y _14954_/X _14955_/Y _14956_/Y _14955_/B vssd1 vssd1 vccd1 vccd1
+ _14959_/A sky130_fd_sc_hd__a32oi_4
XFILLER_48_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12659__A _16157_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19152__D _19329_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__A _11568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13908_ _13820_/X _13907_/X _22761_/Q _14383_/A vssd1 vssd1 vccd1 vccd1 _14465_/B
+ sky130_fd_sc_hd__o211ai_4
X_17676_ _15840_/X _17439_/X _17531_/D vssd1 vssd1 vccd1 vccd1 _17678_/D sky130_fd_sc_hd__o21ai_1
XFILLER_78_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14888_ _14884_/X _14885_/Y _14886_/Y _14887_/Y vssd1 vssd1 vccd1 vccd1 _14930_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12378__B _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19415_ _19261_/Y _19412_/Y _19413_/X _19414_/Y vssd1 vssd1 vccd1 vccd1 _19556_/A
+ sky130_fd_sc_hd__o22ai_4
X_16627_ _16627_/A vssd1 vssd1 vccd1 vccd1 _16630_/A sky130_fd_sc_hd__inv_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13839_ _22759_/Q _22758_/Q vssd1 vssd1 vccd1 vccd1 _13892_/A sky130_fd_sc_hd__nor2_2
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13225__A2 _13162_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19346_ _19346_/A _19504_/B _19504_/C _19504_/D vssd1 vssd1 vccd1 vccd1 _19346_/Y
+ sky130_fd_sc_hd__nand4_1
X_16558_ _15638_/X _16552_/A _16313_/X _16296_/Y vssd1 vssd1 vccd1 vccd1 _16561_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12433__B1 _12413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19361__A1 _12234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18164__A2 _12174_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11787__A2 _12165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15509_ _15500_/A _15500_/B _15506_/Y _15508_/X vssd1 vssd1 vccd1 vccd1 _15510_/C
+ sky130_fd_sc_hd__o211ai_2
X_19277_ _19131_/B _19131_/A _19147_/X vssd1 vssd1 vccd1 vccd1 _19295_/B sky130_fd_sc_hd__o21ai_1
XFILLER_148_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16489_ _16489_/A _16770_/A _16771_/A vssd1 vssd1 vccd1 vccd1 _16489_/X sky130_fd_sc_hd__and3_2
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17911__A2 _17227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18228_ _18228_/A _18228_/B vssd1 vssd1 vccd1 vccd1 _18228_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14725__A2 _14911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19113__A1 _12064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12736__A1 _12734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17124__B1 _17123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18159_ _15888_/X _18156_/X _18365_/A _18158_/X _18125_/X vssd1 vssd1 vccd1 vccd1
+ _18159_/X sky130_fd_sc_hd__o221a_1
XFILLER_11_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17675__A1 _16585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18512__C _18512_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21170_ _21700_/A _21701_/A vssd1 vssd1 vccd1 vccd1 _21820_/A sky130_fd_sc_hd__or2_2
XANTENNA__16313__B _20092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20121_ _20121_/A _20121_/B _20121_/C vssd1 vssd1 vccd1 vccd1 _20154_/B sky130_fd_sc_hd__nand3_2
XFILLER_89_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17128__C _17407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20052_ _20059_/A _20059_/B _22927_/Q vssd1 vssd1 vccd1 vccd1 _20052_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15989__A1 _11912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1111 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater130 _22870_/Q vssd1 vssd1 vccd1 vccd1 _22858_/D sky130_fd_sc_hd__clkbuf_2
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater141 _22765_/CLK vssd1 vssd1 vccd1 vccd1 _22761_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_86_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater152 _22747_/CLK vssd1 vssd1 vccd1 vccd1 _22813_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__17144__B _17401_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater163 _22738_/CLK vssd1 vssd1 vccd1 vccd1 _22802_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11475__A1 _11818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11475__B2 _11474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20954_ _20990_/A _20954_/B vssd1 vssd1 vccd1 vccd1 _21007_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20885_ _20816_/B _20816_/A _20812_/Y _20818_/X vssd1 vssd1 vccd1 vccd1 _20887_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22624_ _22800_/Q input42/X _22630_/S vssd1 vssd1 vccd1 vccd1 _22625_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14964__A2 _13746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_111 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22555_ _22555_/A vssd1 vssd1 vccd1 vccd1 _22769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21506_ _21332_/A _21332_/B _21332_/C _21386_/A _21386_/C vssd1 vssd1 vccd1 vccd1
+ _21658_/C sky130_fd_sc_hd__a32oi_4
XFILLER_155_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22486_ _22739_/Q input45/X _22486_/S vssd1 vssd1 vccd1 vccd1 _22487_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15913__B2 _16011_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21437_ _21437_/A _21437_/B vssd1 vssd1 vccd1 vccd1 _21438_/A sky130_fd_sc_hd__or2_1
XANTENNA__14192__A3 _14911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12170_ _12170_/A vssd1 vssd1 vccd1 vccd1 _12170_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__17319__B _17523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21368_ _21173_/Y _21449_/A _21638_/B _21372_/B _13630_/A vssd1 vssd1 vccd1 vccd1
+ _21369_/D sky130_fd_sc_hd__o2111ai_1
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20319_ _20319_/A _20319_/B vssd1 vssd1 vccd1 vccd1 _20319_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21299_ _21299_/A _21299_/B _21683_/A vssd1 vssd1 vccd1 vccd1 _21299_/X sky130_fd_sc_hd__and3_1
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _15860_/A _15860_/B vssd1 vssd1 vccd1 vccd1 _15861_/C sky130_fd_sc_hd__nand2_1
XFILLER_77_857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20973__A1 _20972_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20973__B2 _20972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input21_A wb_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14811_ _14808_/Y _14809_/Y _14810_/X vssd1 vssd1 vccd1 vccd1 _14813_/A sky130_fd_sc_hd__a21o_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _20359_/C vssd1 vssd1 vccd1 vccd1 _15792_/C sky130_fd_sc_hd__buf_2
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _17530_/A vssd1 vssd1 vccd1 vccd1 _17833_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11954_ _15476_/A vssd1 vssd1 vccd1 vccd1 _19016_/A sky130_fd_sc_hd__buf_4
X_14742_ _14651_/Y _14638_/Y _14649_/B vssd1 vssd1 vccd1 vccd1 _14747_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__16929__B1 _16930_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20725__A1 _20806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17461_ _15887_/X _17981_/D _20972_/A _19482_/A _17591_/A vssd1 vssd1 vccd1 vccd1
+ _17466_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_17_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14673_ _14622_/X _14636_/D _14672_/X vssd1 vssd1 vccd1 vccd1 _14673_/Y sky130_fd_sc_hd__a21oi_1
X_11885_ _11894_/A _11894_/B _11895_/B _11895_/C vssd1 vssd1 vccd1 vccd1 _11886_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19200_ _19200_/A _19200_/B vssd1 vssd1 vccd1 vccd1 _19201_/C sky130_fd_sc_hd__nand2_1
XANTENNA__19328__D1 _18896_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16412_ _16657_/B _16412_/B _16657_/C vssd1 vssd1 vccd1 vccd1 _16686_/A sky130_fd_sc_hd__nand3_2
X_13624_ _13633_/B _13624_/B _13633_/C _21866_/C vssd1 vssd1 vccd1 vccd1 _13625_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_189_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22478__A1 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17392_ _16778_/X _16779_/X _17532_/C _17532_/D vssd1 vssd1 vccd1 vccd1 _17535_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_186_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19131_ _19131_/A _19131_/B vssd1 vssd1 vccd1 vccd1 _19134_/A sky130_fd_sc_hd__nand2_1
X_16343_ _16336_/Y _16337_/X _15566_/X vssd1 vssd1 vccd1 vccd1 _16355_/A sky130_fd_sc_hd__o21a_1
X_13555_ _13556_/A _13556_/C _13556_/B vssd1 vssd1 vccd1 vccd1 _13558_/A sky130_fd_sc_hd__a21o_1
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13103__A _22842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12506_ _12299_/X _12323_/Y _12346_/Y _12357_/Y vssd1 vssd1 vccd1 vccd1 _12506_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_173_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19062_ _19062_/A _19062_/B vssd1 vssd1 vccd1 vccd1 _19063_/C sky130_fd_sc_hd__nand2_1
X_16274_ _16274_/A vssd1 vssd1 vccd1 vccd1 _16275_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13486_ _13659_/C _21665_/D vssd1 vssd1 vccd1 vccd1 _13492_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18013_ _18053_/A _18053_/B vssd1 vssd1 vccd1 vccd1 _18015_/A sky130_fd_sc_hd__nand2_1
XFILLER_185_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15225_ _15223_/B _15224_/X _15223_/A vssd1 vssd1 vccd1 vccd1 _15225_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12437_ _12437_/A vssd1 vssd1 vccd1 vccd1 _15558_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_66_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15156_ _14865_/A _14865_/B _15188_/A _15154_/X _15155_/X vssd1 vssd1 vccd1 vccd1
+ _15156_/Y sky130_fd_sc_hd__a2111oi_4
XFILLER_153_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12368_ _22695_/Q _22693_/Q _22692_/Q _12368_/D vssd1 vssd1 vccd1 vccd1 _16323_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_126_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _14107_/A vssd1 vssd1 vccd1 vccd1 _14808_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11558__A _15435_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11319_ _18107_/A _18985_/C _11936_/C _16308_/C vssd1 vssd1 vccd1 vccd1 _11319_/Y
+ sky130_fd_sc_hd__nand4_4
X_19964_ _20025_/A _19926_/A _19928_/B vssd1 vssd1 vccd1 vccd1 _19965_/B sky130_fd_sc_hd__o21ai_1
XFILLER_114_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15087_ _15088_/A _15088_/B _15089_/A vssd1 vssd1 vccd1 vccd1 _15092_/A sky130_fd_sc_hd__a21o_1
X_12299_ _12457_/A _20323_/A _20694_/A vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__and3_1
XFILLER_141_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18915_ _18915_/A vssd1 vssd1 vccd1 vccd1 _18915_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22402__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14038_ _14033_/X _14523_/B _14036_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 _14039_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_80_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19895_ _19768_/B _18030_/A _18029_/D _19945_/C _19909_/B vssd1 vssd1 vccd1 vccd1
+ _19917_/A sky130_fd_sc_hd__a41o_2
XFILLER_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14891__A1 _15058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18846_ _11704_/X _11738_/X _15458_/A _19358_/C _19358_/D vssd1 vssd1 vccd1 vccd1
+ _19014_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_95_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18777_ _19941_/A vssd1 vssd1 vccd1 vccd1 _19983_/A sky130_fd_sc_hd__clkbuf_2
X_15989_ _11912_/A _15450_/X _15988_/Y vssd1 vssd1 vccd1 vccd1 _16049_/A sky130_fd_sc_hd__o21ai_2
XFILLER_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11293__A _22955_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19031__B1 _19012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17728_ _17728_/A vssd1 vssd1 vccd1 vccd1 _17922_/A sky130_fd_sc_hd__buf_2
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17659_ _17661_/A _17661_/B _17660_/A _17660_/B vssd1 vssd1 vccd1 vccd1 _17665_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__17593__B1 _17591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22469__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20670_ _20670_/A _20670_/B vssd1 vssd1 vccd1 vccd1 _22914_/D sky130_fd_sc_hd__nor2_2
XFILLER_195_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19329_ _19329_/A _19329_/B _19329_/C _19329_/D vssd1 vssd1 vccd1 vccd1 _19330_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__16148__A1 _16131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22340_ _22336_/A _22341_/A _22341_/C vssd1 vssd1 vccd1 vccd1 _22340_/X sky130_fd_sc_hd__o21a_1
XFILLER_164_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19619__B _19619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_3_0_bq_clk_i clkbuf_3_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_136_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13906__B1 _22761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13948__A _13948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22271_ _22271_/A _22271_/B vssd1 vssd1 vccd1 vccd1 _22272_/B sky130_fd_sc_hd__nor2_1
XFILLER_191_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21222_ _21212_/Y _21220_/X _21237_/A _21369_/A vssd1 vssd1 vccd1 vccd1 _21222_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17648__B2 _15919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16305__D1 _20593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12571__B _12571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__A _15901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21153_ _22946_/Q _21157_/B vssd1 vssd1 vccd1 vccd1 _21154_/B sky130_fd_sc_hd__xnor2_2
XFILLER_171_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20104_ _12697_/A _16300_/A _20093_/A vssd1 vssd1 vccd1 vccd1 _20107_/A sky130_fd_sc_hd__o21ai_2
XFILLER_160_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18896__D _19587_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21084_ _21017_/C _21083_/A _21083_/B _21081_/C _21083_/X vssd1 vssd1 vccd1 vccd1
+ _21086_/B sky130_fd_sc_hd__a32o_2
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20035_ _20035_/A _20035_/B vssd1 vssd1 vccd1 vccd1 _22906_/D sky130_fd_sc_hd__xor2_1
XFILLER_101_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17820__A1 _17731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17820__B2 _15941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20012__C _20012_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ _22034_/A _21986_/B _21986_/C _22172_/A vssd1 vssd1 vccd1 vccd1 _21987_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_54_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16387__A1 _15339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20937_ _20937_/A vssd1 vssd1 vccd1 vccd1 _20938_/C sky130_fd_sc_hd__inv_2
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11734_/A vssd1 vssd1 vccd1 vccd1 _16257_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_187_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ _20869_/A _20869_/B _20869_/C _20869_/D vssd1 vssd1 vccd1 vccd1 _20941_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19325__A1 _18980_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22953__CLK _22964_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21668__C1 _13630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22607_ _22607_/A vssd1 vssd1 vccd1 vccd1 _22792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20799_ _20799_/A _20799_/B _20869_/A _20799_/D vssd1 vssd1 vccd1 vccd1 _20869_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_128_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13340_ _13340_/A vssd1 vssd1 vccd1 vccd1 _13340_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12465__C _20478_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22538_ _22584_/S vssd1 vssd1 vccd1 vccd1 _22547_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_167_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13271_ _13271_/A vssd1 vssd1 vccd1 vccd1 _21853_/A sky130_fd_sc_hd__buf_2
XFILLER_154_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22469_ _14359_/X input37/X _22475_/S vssd1 vssd1 vccd1 vccd1 _22470_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15010_ _15010_/A _15115_/C _15010_/C _15069_/A vssd1 vssd1 vccd1 vccd1 _15010_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12176__A2 _12174_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12222_ _12230_/C vssd1 vssd1 vccd1 vccd1 _18227_/C sky130_fd_sc_hd__inv_2
XFILLER_108_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input69_A x[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18300__A2 _18305_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12153_ _18339_/B vssd1 vssd1 vccd1 vccd1 _19016_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_29_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16311__A1 _15888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16311__B2 _15887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16961_ _16939_/Y _16945_/X _16978_/B vssd1 vssd1 vccd1 vccd1 _16961_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__15792__B _15792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ _12084_/A _12084_/B vssd1 vssd1 vccd1 vccd1 _12086_/B sky130_fd_sc_hd__nand2_1
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22396__A0 _16322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18700_ _18695_/X _18696_/X _19329_/A _18692_/Y _15991_/D vssd1 vssd1 vccd1 vccd1
+ _18702_/B sky130_fd_sc_hd__o2111ai_1
X_15912_ _15978_/A _15978_/B _15912_/C _17407_/A vssd1 vssd1 vccd1 vccd1 _16011_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19680_ _19680_/A vssd1 vssd1 vccd1 vccd1 _20025_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16892_ _16892_/A _16892_/B _16892_/C _17065_/A vssd1 vssd1 vccd1 vccd1 _16899_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_134_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16400__C _16400_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18631_ _18810_/D _18303_/A _18303_/B _19504_/C _18459_/C vssd1 vssd1 vccd1 vccd1
+ _18953_/A sky130_fd_sc_hd__a32o_2
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15843_ _15944_/A _15944_/C vssd1 vssd1 vccd1 vccd1 _15843_/Y sky130_fd_sc_hd__nand2_2
XFILLER_49_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14625__B2 _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11439__A1 _14429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18562_ _18565_/A _18765_/B _18568_/B _18568_/C vssd1 vssd1 vccd1 vccd1 _18564_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _18328_/A _15774_/B _15774_/C _15774_/D vssd1 vssd1 vccd1 vccd1 _15775_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12986_ _20593_/C vssd1 vssd1 vccd1 vccd1 _20793_/A sky130_fd_sc_hd__buf_2
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _17513_/A _17513_/B _17513_/C vssd1 vssd1 vccd1 vccd1 _17603_/D sky130_fd_sc_hd__nand3_1
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14725_ _14892_/D _14911_/C _14911_/A _14727_/B _14727_/C vssd1 vssd1 vccd1 vccd1
+ _14726_/D sky130_fd_sc_hd__a32o_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _18493_/A vssd1 vssd1 vccd1 vccd1 _19624_/A sky130_fd_sc_hd__clkbuf_4
X_11937_ _11704_/X _11705_/X _11936_/A _11707_/A vssd1 vssd1 vccd1 vccd1 _11938_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _17444_/A vssd1 vssd1 vccd1 vccd1 _17731_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11868_ _18459_/C _17085_/C _16106_/B _12050_/B vssd1 vssd1 vccd1 vccd1 _11868_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_33_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14656_ _14655_/B _14656_/B _14656_/C vssd1 vssd1 vccd1 vccd1 _14752_/A sky130_fd_sc_hd__nand3b_1
XFILLER_21_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12939__A1 _20576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11560__B _15539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13607_ _13552_/A _13512_/B _13614_/B _13614_/A vssd1 vssd1 vccd1 vccd1 _13608_/C
+ sky130_fd_sc_hd__o211ai_1
X_17375_ _17375_/A vssd1 vssd1 vccd1 vccd1 _17375_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11799_ _11799_/A _11799_/B _11799_/C vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__nand3_2
X_14587_ _14777_/C _14808_/A _14590_/B _14785_/A vssd1 vssd1 vccd1 vccd1 _14605_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18624__A _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19114_ _18778_/B _18023_/A _19113_/X _18830_/B vssd1 vssd1 vccd1 vccd1 _19114_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_192_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16326_ _16344_/A vssd1 vssd1 vccd1 vccd1 _16996_/A sky130_fd_sc_hd__clkbuf_2
X_13538_ _13538_/A _13538_/B _13538_/C vssd1 vssd1 vccd1 vccd1 _13539_/A sky130_fd_sc_hd__nand3_1
XFILLER_173_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15889__B1 _12968_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19045_ _19045_/A vssd1 vssd1 vccd1 vccd1 _19046_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12094__D _12094_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16257_ _16257_/A _16257_/B _16257_/C _16257_/D vssd1 vssd1 vccd1 vccd1 _16257_/Y
+ sky130_fd_sc_hd__nand4_4
X_13469_ _13469_/A vssd1 vssd1 vccd1 vccd1 _13550_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12672__A _12672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16550__A1 _12827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15208_ _15181_/A _15181_/B _15200_/B vssd1 vssd1 vccd1 vccd1 _15209_/A sky130_fd_sc_hd__o21ba_1
X_16188_ _16024_/A _16090_/B _16092_/Y _16093_/X vssd1 vssd1 vccd1 vccd1 _16188_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_114_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11288__A _22953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15139_ _15173_/A _15139_/B vssd1 vssd1 vccd1 vccd1 _15139_/Y sky130_fd_sc_hd__nor2_1
X_19947_ _19946_/C _19946_/A _19946_/B vssd1 vssd1 vccd1 vccd1 _19948_/B sky130_fd_sc_hd__a21o_1
XFILLER_141_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22387__A0 _12320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19878_ _19878_/A _19878_/B vssd1 vssd1 vccd1 vccd1 _19878_/Y sky130_fd_sc_hd__nand2_2
XFILLER_110_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22826__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12875__B1 _16160_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18829_ _18830_/B _18830_/C _18778_/B _18814_/X vssd1 vssd1 vccd1 vccd1 _18829_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21288__A_N _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21840_ _21730_/C _21730_/D _21775_/Y vssd1 vssd1 vccd1 vccd1 _21841_/B sky130_fd_sc_hd__a21oi_1
XFILLER_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13824__C1 _13823_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18358__A2 _12111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21771_ _21771_/A _21771_/B _21771_/C vssd1 vssd1 vccd1 vccd1 _21771_/X sky130_fd_sc_hd__and3_1
XFILLER_64_882 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14765__C _14765_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20722_ _20778_/B _20812_/A vssd1 vssd1 vccd1 vccd1 _20731_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17141__C _17532_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20653_ _20653_/A _20658_/A vssd1 vssd1 vccd1 vccd1 _20656_/A sky130_fd_sc_hd__nand2_1
XFILLER_177_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20584_ _20584_/A _20584_/B _20584_/C vssd1 vssd1 vccd1 vccd1 _20584_/Y sky130_fd_sc_hd__nand3_1
XFILLER_176_272 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14781__B _14857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18530__A2 _11702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22323_ _22323_/A _22323_/B _22685_/Q vssd1 vssd1 vccd1 vccd1 _22324_/B sky130_fd_sc_hd__and3_1
XANTENNA__20873__B1 _12761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_743 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16054__A _18984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22254_ _22245_/X _22246_/Y _22146_/A vssd1 vssd1 vccd1 vccd1 _22258_/A sky130_fd_sc_hd__a21oi_1
XFILLER_164_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15893__A _15893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21205_ _13321_/X _21184_/X _21198_/Y _21204_/Y vssd1 vssd1 vccd1 vccd1 _21238_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__18294__A1 _11818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22185_ _22108_/Y _22181_/Y _22220_/A _22183_/Y _22265_/C vssd1 vssd1 vccd1 vccd1
+ _22188_/A sky130_fd_sc_hd__o2111a_1
XFILLER_144_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21136_ _21118_/A _21133_/Y _21135_/Y vssd1 vssd1 vccd1 vccd1 _21141_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__22378__A0 _12493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14855__A1 _14942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14855__B2 _14942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11669__A1 _15484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21067_ _21067_/A _21067_/B _21067_/C _21067_/D vssd1 vssd1 vccd1 vccd1 _21067_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_59_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16220__C _16947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20018_ _20018_/A _20018_/B vssd1 vssd1 vccd1 vccd1 _20021_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11645__B _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12840_ _12574_/A _16708_/A _12820_/Y vssd1 vssd1 vccd1 vccd1 _20142_/A sky130_fd_sc_hd__o21ai_4
XFILLER_74_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12771_/A vssd1 vssd1 vccd1 vccd1 _12772_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_15_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21969_ _21972_/B _21972_/C _21967_/X _21968_/Y vssd1 vssd1 vccd1 vccd1 _22031_/B
+ sky130_fd_sc_hd__o2bb2ai_4
XANTENNA__22550__A0 _14863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21353__A1 _13326_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11749_/A _11750_/A vssd1 vssd1 vccd1 vccd1 _16447_/A sky130_fd_sc_hd__nand2_2
X_14510_ _14510_/A _14629_/B _14510_/C _14808_/B vssd1 vssd1 vccd1 vccd1 _14512_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_70_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _16786_/A vssd1 vssd1 vccd1 vccd1 _17379_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__B _11380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14441_ _18259_/B _16481_/C _14435_/Y _22952_/D vssd1 vssd1 vccd1 vccd1 _22662_/A
+ sky130_fd_sc_hd__a31o_1
X_11653_ _15694_/A vssd1 vssd1 vccd1 vccd1 _18666_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_120_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12907__D _20355_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17160_ _17270_/A _17270_/B _17180_/B _17180_/C vssd1 vssd1 vccd1 vccd1 _17161_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18476__B1_N _18305_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14372_ _22797_/Q vssd1 vssd1 vccd1 vccd1 _18698_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11584_ _11792_/A _11792_/B vssd1 vssd1 vccd1 vccd1 _11585_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16111_ _16111_/A _16111_/B vssd1 vssd1 vccd1 vccd1 _16169_/D sky130_fd_sc_hd__nand2_1
X_13323_ _13316_/X _13317_/X _13300_/Y vssd1 vssd1 vccd1 vccd1 _13324_/A sky130_fd_sc_hd__o21ai_1
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17091_ _17091_/A vssd1 vssd1 vccd1 vccd1 _17460_/A sky130_fd_sc_hd__buf_2
XFILLER_128_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16042_ _15967_/X _15971_/Y _16020_/Y _16021_/Y vssd1 vssd1 vccd1 vccd1 _16043_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13254_ _22849_/Q vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12205_ _16477_/A _16477_/B vssd1 vssd1 vccd1 vccd1 _15838_/A sky130_fd_sc_hd__nand2_2
XANTENNA__20616__B1 _15938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18285__A1 _11308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17088__A2 _17431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18285__B2 _15531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185_ _13185_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13430_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22849__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19801_ _19864_/A _19864_/B _19866_/A _19865_/B vssd1 vssd1 vccd1 vccd1 _19804_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12120__A2_N _12123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12136_ _12009_/A _18655_/A _12128_/X _12126_/X _12131_/Y vssd1 vssd1 vccd1 vccd1
+ _12138_/B sky130_fd_sc_hd__o221ai_1
XFILLER_150_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17993_ _18061_/A _18061_/B _18062_/D _18062_/C vssd1 vssd1 vccd1 vccd1 _17994_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14846__A1 _14552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19732_ _19649_/B _19643_/Y _19649_/C vssd1 vssd1 vccd1 vccd1 _19736_/C sky130_fd_sc_hd__o21ai_1
X_16944_ _15325_/X _15326_/X _12689_/A _19199_/B _19199_/C vssd1 vssd1 vccd1 vccd1
+ _16944_/Y sky130_fd_sc_hd__o2111ai_4
X_12067_ _16192_/D _18830_/A _18305_/B _17006_/D vssd1 vssd1 vccd1 vccd1 _12069_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16130__C _20745_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19663_ _19663_/A _19663_/B vssd1 vssd1 vccd1 vccd1 _19664_/C sky130_fd_sc_hd__nor2_1
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16875_ _17313_/B vssd1 vssd1 vccd1 vccd1 _17006_/A sky130_fd_sc_hd__buf_2
XFILLER_38_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18614_ _18610_/X _18611_/Y _18618_/B vssd1 vssd1 vccd1 vccd1 _18616_/A sky130_fd_sc_hd__o21ai_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17523__A _17523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15826_ _15826_/A _15849_/A _15826_/C vssd1 vssd1 vccd1 vccd1 _15826_/Y sky130_fd_sc_hd__nand3_2
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19594_ _19594_/A _19594_/B vssd1 vssd1 vccd1 vccd1 _19594_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18545_ _18156_/X _16276_/X _18091_/Y _18360_/X _18544_/X vssd1 vssd1 vccd1 vccd1
+ _18546_/C sky130_fd_sc_hd__o32a_2
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _15854_/A _15854_/B _15864_/B _15756_/X vssd1 vssd1 vccd1 vccd1 _15758_/C
+ sky130_fd_sc_hd__a31oi_4
XFILLER_18_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17548__B1 _17546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22541__A0 _14362_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ _12981_/D vssd1 vssd1 vccd1 vccd1 _13024_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17012__A2 _16732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14708_ _14815_/C _14857_/A _14951_/A _14708_/D vssd1 vssd1 vccd1 vccd1 _14711_/D
+ sky130_fd_sc_hd__nand4_1
X_18476_ _18305_/A _18459_/A _18305_/D vssd1 vssd1 vccd1 vccd1 _18478_/C sky130_fd_sc_hd__a21bo_1
X_15688_ _15682_/Y _15433_/A _15683_/Y _15687_/Y vssd1 vssd1 vccd1 vccd1 _15761_/B
+ sky130_fd_sc_hd__o22ai_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17427_ _17427_/A vssd1 vssd1 vccd1 vccd1 _17427_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ _14650_/A _14740_/B _14650_/C vssd1 vssd1 vccd1 vccd1 _14649_/B sky130_fd_sc_hd__nand3_1
XFILLER_147_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17358_ _17372_/C _17357_/X _22897_/Q vssd1 vssd1 vccd1 vccd1 _17358_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16309_ _16308_/X _15634_/Y _15632_/Y _15319_/B vssd1 vssd1 vccd1 vccd1 _16309_/Y
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ _16737_/X _16015_/A _17293_/B _17449_/A vssd1 vssd1 vccd1 vccd1 _17290_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_134_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19028_ _19012_/X _19013_/X _19029_/A _19037_/A vssd1 vssd1 vccd1 vccd1 _19028_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16826__A2 _16825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13664__C _21878_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14122__A _14122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22941_ _22943_/CLK _22941_/D vssd1 vssd1 vccd1 vccd1 _22941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22872_ _22916_/CLK _22872_/D vssd1 vssd1 vccd1 vccd1 _22872_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__19351__C _19351_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14776__B _22766_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21823_ _21834_/C _21834_/D vssd1 vssd1 vccd1 vccd1 _21823_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22532__A0 _13736_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11481__A _22790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21754_ _21486_/A _21596_/B _21591_/Y vssd1 vssd1 vccd1 vccd1 _21758_/B sky130_fd_sc_hd__o21ai_1
XFILLER_24_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20705_ _20596_/C _20596_/A _20703_/X _20704_/Y vssd1 vssd1 vccd1 vccd1 _20709_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__15888__A _15888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21685_ _21684_/X _21546_/A _21531_/X _21534_/Y vssd1 vssd1 vccd1 vccd1 _21688_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_196_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13576__A1 _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13576__B2 _13434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20636_ _20574_/X _20575_/X _20631_/Y _20737_/A vssd1 vssd1 vccd1 vccd1 _20636_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_165_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20567_ _20522_/A _20522_/B _20522_/C vssd1 vssd1 vccd1 vccd1 _20567_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_165_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22306_ _22306_/A _22306_/B _22306_/C _22263_/B vssd1 vssd1 vccd1 vccd1 _22307_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_192_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20498_ _20499_/A _20499_/B _20629_/A _20499_/D vssd1 vssd1 vccd1 vccd1 _20500_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18267__A1 _18088_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22237_ _22237_/A _22237_/B vssd1 vssd1 vccd1 vccd1 _22240_/C sky130_fd_sc_hd__nand2_1
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20074__A1 _12761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12551__A2 _12528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22168_ _13305_/A _13305_/B _22306_/B vssd1 vssd1 vccd1 vccd1 _22168_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21119_ _21119_/A _21119_/B _22943_/Q vssd1 vssd1 vccd1 vccd1 _21120_/A sky130_fd_sc_hd__or3b_1
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22099_ _22099_/A _22099_/B vssd1 vssd1 vccd1 vccd1 _22100_/B sky130_fd_sc_hd__nand2_1
X_14990_ _15186_/D vssd1 vssd1 vccd1 vccd1 _14990_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19767__A1 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19767__B2 _19176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13941_ _14110_/B vssd1 vssd1 vccd1 vccd1 _14489_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16660_ _16889_/B _16673_/A vssd1 vssd1 vccd1 vccd1 _16660_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__15789__C1 _16192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872_ _13881_/B vssd1 vssd1 vccd1 vccd1 _13986_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14686__B _14686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19519__B2 _19518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15611_ _15611_/A vssd1 vssd1 vccd1 vccd1 _16611_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12067__A1 _16192_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ _12823_/A vssd1 vssd1 vccd1 vccd1 _16320_/A sky130_fd_sc_hd__clkbuf_4
X_16591_ _16586_/A _16879_/A _16590_/X vssd1 vssd1 vccd1 vccd1 _16598_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__12067__B2 _17006_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22523__A0 _13725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__A _16515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__A _18482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18330_ _18330_/A vssd1 vssd1 vccd1 vccd1 _18330_/X sky130_fd_sc_hd__buf_4
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15542_ _15538_/X _15541_/X _12968_/B vssd1 vssd1 vccd1 vccd1 _15542_/X sky130_fd_sc_hd__a21o_2
XFILLER_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _13044_/C vssd1 vssd1 vccd1 vccd1 _12754_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _18261_/A _18261_/B _18600_/A vssd1 vssd1 vccd1 vccd1 _18261_/X sky130_fd_sc_hd__and3_1
X_11705_ _11738_/A vssd1 vssd1 vccd1 vccd1 _11705_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15556__A2 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15473_ _15309_/B _15472_/X _15574_/C _19016_/A _17246_/A vssd1 vssd1 vccd1 vccd1
+ _15474_/C sky130_fd_sc_hd__o2111ai_2
X_12685_ _16498_/A vssd1 vssd1 vccd1 vccd1 _16067_/D sky130_fd_sc_hd__clkbuf_2
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _17603_/B vssd1 vssd1 vccd1 vccd1 _17518_/C sky130_fd_sc_hd__inv_2
XFILLER_175_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11636_ _11636_/A vssd1 vssd1 vccd1 vccd1 _11636_/X sky130_fd_sc_hd__buf_2
X_14424_ _22717_/Q _14418_/X _14410_/X _22749_/Q _14423_/X vssd1 vssd1 vccd1 vccd1
+ _14424_/X sky130_fd_sc_hd__a221o_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18192_ _18192_/A vssd1 vssd1 vccd1 vccd1 _19353_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12934__B _16078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17143_ _15495_/X _16226_/B _12046_/X _16242_/X vssd1 vssd1 vccd1 vccd1 _17401_/C
+ sky130_fd_sc_hd__o31ai_4
X_11567_ _11561_/X _11563_/X _11565_/Y _11566_/X vssd1 vssd1 vccd1 vccd1 _11899_/A
+ sky130_fd_sc_hd__a211o_2
X_14355_ _14355_/A vssd1 vssd1 vccd1 vccd1 _14355_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14532__C_N _22863_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13306_ _13297_/A _21329_/A _13319_/A vssd1 vssd1 vccd1 vccd1 _13309_/B sky130_fd_sc_hd__a21oi_2
X_17074_ _22896_/Q vssd1 vssd1 vccd1 vccd1 _17220_/A sky130_fd_sc_hd__inv_2
XFILLER_171_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14286_ _14054_/A _14115_/B _14115_/C _14285_/A _14285_/B vssd1 vssd1 vccd1 vccd1
+ _14288_/B sky130_fd_sc_hd__a32o_1
XFILLER_144_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11498_ _11792_/B vssd1 vssd1 vccd1 vccd1 _18131_/C sky130_fd_sc_hd__buf_2
XFILLER_196_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20870__C _20870_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12527__C1 _16488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16025_ _15970_/A _15970_/B _15927_/Y vssd1 vssd1 vccd1 vccd1 _16026_/A sky130_fd_sc_hd__o21ai_1
X_13237_ _13423_/A _21259_/B _21259_/C vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__or3_1
XFILLER_108_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12950__A _20390_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16269__B1 _11568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20065__A1 _20064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16808__A2 _15933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13168_ _13513_/A _21448_/A _13168_/C _21595_/B vssd1 vssd1 vccd1 vccd1 _13465_/A
+ sky130_fd_sc_hd__nand4_4
XANTENNA__17237__B _17631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14819__A1 _15188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11566__A _11818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _12116_/X _16014_/A _11634_/A _16016_/A vssd1 vssd1 vccd1 vccd1 _12119_/X
+ sky130_fd_sc_hd__o22a_2
X_17976_ _19454_/C vssd1 vssd1 vccd1 vccd1 _18028_/A sky130_fd_sc_hd__buf_2
XFILLER_112_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13099_ _13095_/X _13099_/B _14380_/A vssd1 vssd1 vccd1 vccd1 _13101_/A sky130_fd_sc_hd__nand3b_1
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1080 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19758__A1 _22919_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15492__A1 _12758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17218__C1 _17373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19715_ _19793_/C _19792_/A _19615_/A _19714_/X vssd1 vssd1 vccd1 vccd1 _19715_/X
+ sky130_fd_sc_hd__a31o_1
X_16927_ _16920_/Y _16922_/X _16923_/Y _16926_/Y vssd1 vssd1 vccd1 vccd1 _17341_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11285__B _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14299__D input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19646_ _19540_/A _19540_/B _19540_/C _19543_/A vssd1 vssd1 vccd1 vccd1 _19650_/B
+ sky130_fd_sc_hd__a31o_1
X_16858_ _16858_/A vssd1 vssd1 vccd1 vccd1 _16869_/B sky130_fd_sc_hd__inv_2
XFILLER_26_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15809_ _12772_/X _12774_/X _14432_/A _15808_/X _11672_/X vssd1 vssd1 vccd1 vccd1
+ _15812_/C sky130_fd_sc_hd__o221a_2
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19577_ _19577_/A _19577_/B vssd1 vssd1 vccd1 vccd1 _19663_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16789_ _17636_/A _16179_/X _16781_/Y _16787_/Y _16788_/X vssd1 vssd1 vccd1 vccd1
+ _16789_/X sky130_fd_sc_hd__o311a_1
XFILLER_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15795__A2 _12607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16992__A1 _11504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18528_ _18495_/A _18495_/B _18326_/Y vssd1 vssd1 vccd1 vccd1 _18528_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18459_ _18459_/A _19687_/C _18459_/C vssd1 vssd1 vccd1 vccd1 _18464_/A sky130_fd_sc_hd__and3_1
XANTENNA__15547__A2 _15546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16744__A1 _16742_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20540__A2 _15890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21470_ _21578_/A _21307_/C _21580_/B vssd1 vssd1 vccd1 vccd1 _21476_/A sky130_fd_sc_hd__a21o_1
XFILLER_53_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20421_ _20286_/A _20286_/B _20286_/C _20298_/B _20319_/B vssd1 vssd1 vccd1 vccd1
+ _20423_/C sky130_fd_sc_hd__a32oi_4
XFILLER_193_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13659__C _13659_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13021__A _20697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20352_ _20457_/B _20457_/A _20083_/X _20339_/A vssd1 vssd1 vccd1 vccd1 _20353_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20780__C _20853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20283_ _20284_/B _20284_/C _20177_/A _20429_/B vssd1 vssd1 vccd1 vccd1 _20401_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__19346__C _19504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22022_ _22016_/X _22017_/X _22018_/Y _22021_/B vssd1 vssd1 vccd1 vccd1 _22290_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_114_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_48 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18259__A _18259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22924_ _22948_/CLK _22924_/D vssd1 vssd1 vccd1 vccd1 _22924_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22855_ _22937_/CLK _22867_/Q vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17313__D _17313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21806_ _22229_/B _13630_/A _21667_/Y _21805_/X vssd1 vssd1 vccd1 vccd1 _21806_/X
+ sky130_fd_sc_hd__a31o_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15114__C _15114_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22786_ _22787_/CLK _22786_/D vssd1 vssd1 vccd1 vccd1 _22786_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21737_ _21737_/A _21737_/B vssd1 vssd1 vccd1 vccd1 _21737_/Y sky130_fd_sc_hd__nor2_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16735__A1 _11821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12470_ _22690_/Q vssd1 vssd1 vccd1 vccd1 _12470_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_138_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21668_ _21651_/X _21665_/Y _21667_/Y _13630_/A _21990_/B vssd1 vssd1 vccd1 vccd1
+ _21677_/A sky130_fd_sc_hd__o2111a_2
XFILLER_184_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11421_ _11421_/A vssd1 vssd1 vccd1 vccd1 _18319_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_137_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20619_ _20620_/B _20620_/C _20620_/A vssd1 vssd1 vccd1 vccd1 _20621_/A sky130_fd_sc_hd__a21o_1
X_21599_ _21645_/A vssd1 vssd1 vccd1 vccd1 _21846_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14140_ _14238_/B _14239_/B vssd1 vssd1 vccd1 vccd1 _14141_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11352_ _11369_/A _11369_/B _11345_/X _11351_/X vssd1 vssd1 vccd1 vccd1 _11352_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14071_ _14510_/C _14686_/B _14506_/C vssd1 vssd1 vccd1 vccd1 _14071_/Y sky130_fd_sc_hd__nand3_1
XFILLER_153_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11283_ _22787_/Q vssd1 vssd1 vccd1 vccd1 _11860_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_141_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _13022_/A _13022_/B _13022_/C _13022_/D vssd1 vssd1 vccd1 vccd1 _13022_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_105_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input51_A wb_dat_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20598__A2 _17111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17830_ _17890_/B _17831_/C _17831_/A vssd1 vssd1 vccd1 vccd1 _17871_/A sky130_fd_sc_hd__a21o_1
XFILLER_121_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18660__A1 _19199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17761_ _17736_/X _17761_/B _17761_/C vssd1 vssd1 vccd1 vccd1 _17765_/A sky130_fd_sc_hd__and3b_1
XFILLER_121_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14973_ _14970_/X _14971_/Y _14914_/C _14972_/Y vssd1 vssd1 vccd1 vccd1 _14977_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_120_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19500_ _19500_/A vssd1 vssd1 vccd1 vccd1 _19500_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16712_ _20471_/A _20471_/B _16712_/C vssd1 vssd1 vccd1 vccd1 _16712_/X sky130_fd_sc_hd__and3_1
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13924_ _13924_/A vssd1 vssd1 vccd1 vccd1 _13924_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17692_ _17579_/Y _17585_/Y _17583_/Y vssd1 vssd1 vccd1 vccd1 _17693_/C sky130_fd_sc_hd__a21boi_1
XFILLER_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19431_ _19302_/Y _19147_/X _19299_/Y _19663_/A _19430_/X vssd1 vssd1 vccd1 vccd1
+ _19446_/A sky130_fd_sc_hd__o2111ai_2
X_16643_ _16613_/D _17039_/C _16879_/B _16351_/X vssd1 vssd1 vccd1 vccd1 _16644_/C
+ sky130_fd_sc_hd__a31o_2
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13855_ _13761_/B _13707_/A _13707_/B _13845_/B _13810_/C vssd1 vssd1 vccd1 vccd1
+ _13930_/A sky130_fd_sc_hd__o311ai_4
XANTENNA__15777__A2 _11505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17801__A _18044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19362_ _19357_/B _19359_/X _19360_/Y _19361_/Y vssd1 vssd1 vccd1 vccd1 _19362_/Y
+ sky130_fd_sc_hd__a22oi_2
X_12806_ _12596_/A _15637_/A _12817_/A vssd1 vssd1 vccd1 vccd1 _12810_/A sky130_fd_sc_hd__o21ai_2
XFILLER_76_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16574_ _22701_/Q _16320_/A _16320_/B _22702_/Q _15369_/B vssd1 vssd1 vccd1 vccd1
+ _20579_/B sky130_fd_sc_hd__o311ai_4
XFILLER_90_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13786_ _13786_/A _13786_/B vssd1 vssd1 vccd1 vccd1 _14165_/C sky130_fd_sc_hd__nand2_1
XFILLER_43_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18313_ _18313_/A _18313_/B _18677_/C _18677_/B vssd1 vssd1 vccd1 vccd1 _18313_/Y
+ sky130_fd_sc_hd__nand4_4
X_15525_ _12209_/A _12211_/A _16759_/A _16473_/A vssd1 vssd1 vccd1 vccd1 _15589_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_16_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17520__B _17523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19293_ _19293_/A vssd1 vssd1 vccd1 vccd1 _19293_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_163_1043 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15529__A2 _15524_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12460__A1 _16477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12737_ _12737_/A _12737_/B _12950_/B _12737_/D vssd1 vssd1 vccd1 vccd1 _12933_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12945__A _20129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15959__C _17816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14863__C _14863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18259_/B _18258_/A vssd1 vssd1 vccd1 vccd1 _18246_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15321__A _20611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15456_ _11820_/A _15546_/A _15302_/A _15302_/B vssd1 vssd1 vccd1 vccd1 _15457_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_176_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12668_ _12668_/A _12668_/B _12745_/A _12745_/B vssd1 vssd1 vccd1 vccd1 _12741_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14407_ _22711_/Q _14403_/X _14396_/X _22743_/Q _14406_/X vssd1 vssd1 vccd1 vccd1
+ _14407_/X sky130_fd_sc_hd__a221o_1
XFILLER_128_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18175_ _18113_/Y _18114_/X _18163_/Y _18404_/A vssd1 vssd1 vccd1 vccd1 _18181_/A
+ sky130_fd_sc_hd__o211ai_1
X_11619_ _11619_/A _11619_/B _18115_/A vssd1 vssd1 vccd1 vccd1 _11974_/C sky130_fd_sc_hd__nand3_2
XANTENNA__19676__B1 _22918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15387_ _17423_/A _17424_/A _15358_/X vssd1 vssd1 vccd1 vccd1 _15389_/A sky130_fd_sc_hd__a21o_2
X_12599_ _20323_/A vssd1 vssd1 vccd1 vccd1 _16261_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_156_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12383__C _20207_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17126_ _17122_/A _17122_/B _17122_/C _17125_/X vssd1 vssd1 vccd1 vccd1 _17127_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_184_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14338_ _14354_/A vssd1 vssd1 vccd1 vccd1 _14338_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13776__A _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17057_ _17603_/A _17603_/B vssd1 vssd1 vccd1 vccd1 _17058_/B sky130_fd_sc_hd__nor2_1
XFILLER_132_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14269_ _14269_/A _14279_/A _14269_/C _14269_/D vssd1 vssd1 vccd1 vccd1 _14279_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12680__A _20478_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1071 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16008_ _16000_/A _16000_/B _16000_/C _16047_/C _16047_/D vssd1 vssd1 vccd1 vccd1
+ _16008_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15991__A _16129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11296__A _11968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18651__A1 _11598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11727__C _11727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _17959_/A _17959_/B _17959_/C vssd1 vssd1 vccd1 vccd1 _17960_/D sky130_fd_sc_hd__nand3_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20970_ _17928_/A _20843_/X _20967_/Y _20969_/Y vssd1 vssd1 vccd1 vccd1 _20982_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19629_ _19709_/C _19629_/B vssd1 vssd1 vccd1 vccd1 _19630_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22640_ _22640_/A vssd1 vssd1 vccd1 vccd1 _22807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22571_ _22571_/A vssd1 vssd1 vccd1 vccd1 _22580_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_167_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21522_ _21522_/A _21522_/B _21522_/C _21522_/D vssd1 vssd1 vccd1 vccd1 _21524_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_178_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16193__A2 _15978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21453_ _21767_/A _21341_/A _21216_/B _21352_/X vssd1 vssd1 vccd1 vccd1 _21453_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22266__A2 _21594_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20404_ _20403_/A _20403_/B _20403_/C vssd1 vssd1 vccd1 vccd1 _20404_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21384_ _21383_/X _21341_/X _21216_/B _21352_/X _21460_/A vssd1 vssd1 vccd1 vccd1
+ _21385_/B sky130_fd_sc_hd__o221ai_1
XFILLER_174_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11962__B1 _11935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15153__B1 _14942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20335_ _20335_/A _20335_/B _20335_/C vssd1 vssd1 vccd1 vccd1 _20336_/B sky130_fd_sc_hd__and3_1
XFILLER_190_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16062__A _16062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20266_ _20266_/A vssd1 vssd1 vccd1 vccd1 _20397_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22005_ _22007_/A _22007_/B _21909_/A vssd1 vssd1 vccd1 vccd1 _22005_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__17445__A2 _17731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20197_ _20197_/A _20197_/B vssd1 vssd1 vccd1 vccd1 _20197_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15456__A1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11934__A _19316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _18648_/D _18167_/A _18875_/D _18875_/C vssd1 vssd1 vccd1 vccd1 _11970_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22907_ _22949_/CLK _22907_/D vssd1 vssd1 vccd1 vccd1 _22907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13640_ _13647_/A _13640_/B vssd1 vssd1 vccd1 vccd1 _13640_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22838_ _22850_/CLK _22850_/Q vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__22884__D input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12978__C1 _20697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16885__A_N _16884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13571_ _21212_/C vssd1 vssd1 vccd1 vccd1 _21938_/B sky130_fd_sc_hd__clkbuf_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20504__A2 _20123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22769_ _22801_/CLK _22769_/D vssd1 vssd1 vccd1 vccd1 _22769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_630 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12765__A _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15310_ _15302_/B _15306_/Y _15502_/A _15694_/A _15774_/C vssd1 vssd1 vccd1 vccd1
+ _15313_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14683__C _14684_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14719__B1 _13748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12522_/A _12522_/B vssd1 vssd1 vccd1 vccd1 _12523_/A sky130_fd_sc_hd__nand2_1
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16290_ _16290_/A _16596_/A _16595_/B vssd1 vssd1 vccd1 vccd1 _16290_/X sky130_fd_sc_hd__and3_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ _15241_/A _15241_/B vssd1 vssd1 vccd1 vccd1 _15242_/B sky130_fd_sc_hd__nand2_1
X_12453_ _12461_/A _12424_/Y _20323_/B _20466_/B _12449_/Y vssd1 vssd1 vccd1 vccd1
+ _12454_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_185_679 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11404_ _11404_/A _11404_/B _11404_/C _11404_/D vssd1 vssd1 vccd1 vccd1 _16481_/A
+ sky130_fd_sc_hd__nor4_2
XFILLER_138_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15172_ _15173_/A _15173_/B _15173_/C vssd1 vssd1 vccd1 vccd1 _15174_/A sky130_fd_sc_hd__o21ai_2
X_12384_ _12384_/A vssd1 vssd1 vccd1 vccd1 _12550_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11335_ _11404_/C vssd1 vssd1 vccd1 vccd1 _11423_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ _13930_/A _13930_/B _14274_/A vssd1 vssd1 vccd1 vccd1 _14123_/X sky130_fd_sc_hd__a21o_1
X_19980_ _19750_/X _19963_/A _19963_/B _19965_/B vssd1 vssd1 vccd1 vccd1 _20005_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_181_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15695__A1 _15298_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18931_ _18978_/A _18931_/B _18977_/B vssd1 vssd1 vccd1 vccd1 _18932_/C sky130_fd_sc_hd__nand3_1
XFILLER_119_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14054_ _14054_/A _14055_/B vssd1 vssd1 vccd1 vccd1 _14054_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13005_ _13004_/C _13004_/A _13004_/B vssd1 vssd1 vccd1 vccd1 _13006_/B sky130_fd_sc_hd__a21o_1
X_18862_ _18862_/A _18862_/B vssd1 vssd1 vccd1 vccd1 _18869_/D sky130_fd_sc_hd__nand2_1
XFILLER_122_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17813_ _17929_/A vssd1 vssd1 vccd1 vccd1 _19896_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18793_ _18770_/C _18779_/B _18776_/Y vssd1 vssd1 vccd1 vccd1 _18955_/A sky130_fd_sc_hd__a21oi_2
Xclkbuf_4_5_0_bq_clk_i clkbuf_4_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _22944_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_48_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11844__A _15377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17744_ _17744_/A _17826_/B vssd1 vssd1 vccd1 vccd1 _17755_/B sky130_fd_sc_hd__nand2_1
X_14956_ _14952_/Y _14954_/X _14955_/A vssd1 vssd1 vccd1 vccd1 _14956_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_130_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12659__B _20723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_796 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13907_ _13907_/A vssd1 vssd1 vccd1 vccd1 _13907_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17675_ _16585_/A _16585_/B _16016_/X _17564_/B vssd1 vssd1 vccd1 vccd1 _17678_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14887_ _14947_/A _14887_/B _14887_/C vssd1 vssd1 vccd1 vccd1 _14887_/Y sky130_fd_sc_hd__nand3_1
XFILLER_130_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19414_ _19407_/X _19408_/X _19401_/X vssd1 vssd1 vccd1 vccd1 _19414_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12378__C _12378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17531__A _19772_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16626_ _16637_/A _16637_/B vssd1 vssd1 vccd1 vccd1 _16631_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13838_ _13807_/Y _13808_/Y _13830_/Y _13837_/Y vssd1 vssd1 vccd1 vccd1 _13838_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14422__A2 _14418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13225__A3 _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19345_ _11598_/X _16758_/X _17393_/X _11474_/X vssd1 vssd1 vccd1 vccd1 _19455_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_188_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16557_ _16557_/A _16557_/B _16557_/C vssd1 vssd1 vccd1 vccd1 _16599_/C sky130_fd_sc_hd__nand3_4
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13769_ _14110_/C vssd1 vssd1 vccd1 vccd1 _14181_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_189_985 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14593__C _22764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19361__A2 _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15508_ _15502_/C _15502_/D _15507_/X vssd1 vssd1 vccd1 vccd1 _15508_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19276_ _19131_/B _19131_/A _19147_/X _19295_/A vssd1 vssd1 vccd1 vccd1 _19284_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__11787__A3 _11786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16488_ _16488_/A _17139_/A _17140_/A vssd1 vssd1 vccd1 vccd1 _16762_/A sky130_fd_sc_hd__nand3_2
XFILLER_149_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18227_ _18228_/A _18228_/B _18227_/C vssd1 vssd1 vccd1 vccd1 _18227_/X sky130_fd_sc_hd__and3_1
X_15439_ _15439_/A vssd1 vssd1 vccd1 vccd1 _15439_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_129_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17109__D1 _17386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14725__A3 _14911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19113__A2 _19941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20259__A1 _20252_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21456__B1 _13326_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13933__A1 _13948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12736__A2 _12735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18158_ _18995_/A vssd1 vssd1 vccd1 vccd1 _18158_/X sky130_fd_sc_hd__buf_2
XFILLER_7_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17109_ _12827_/X _15617_/X _11672_/A _11666_/X _17386_/B vssd1 vssd1 vccd1 vccd1
+ _17110_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17675__A2 _16585_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18089_ _12162_/Y _12172_/Y _12156_/X vssd1 vssd1 vccd1 vccd1 _18098_/A sky130_fd_sc_hd__a21boi_1
XFILLER_117_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16313__C _16313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20120_ _20120_/A _20120_/B vssd1 vssd1 vccd1 vccd1 _20121_/C sky130_fd_sc_hd__nand2_1
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22034__D _22229_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17128__D _19496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20051_ _20051_/A _20051_/B vssd1 vssd1 vccd1 vccd1 _22907_/D sky130_fd_sc_hd__nor2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16610__A _16996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15989__A2 _15450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater131 _22846_/Q vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11754__A _17280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater142 _22765_/CLK vssd1 vssd1 vccd1 vccd1 _22799_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater153 _22749_/CLK vssd1 vssd1 vccd1 vccd1 _22812_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater164 _22801_/CLK vssd1 vssd1 vccd1 vccd1 _22738_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11473__B _18093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ _20951_/X _20989_/A _20894_/B _20894_/Y vssd1 vssd1 vccd1 vccd1 _20954_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_26_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _20884_/A _20884_/B _20884_/C vssd1 vssd1 vccd1 vccd1 _20887_/B sky130_fd_sc_hd__nor3_1
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17160__B _17270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22623_ _22623_/A vssd1 vssd1 vccd1 vccd1 _22799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22554_ _22769_/Q input43/X _22558_/S vssd1 vssd1 vccd1 vccd1 _22555_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21505_ _21508_/B _21649_/B _21508_/A vssd1 vssd1 vccd1 vccd1 _21658_/B sky130_fd_sc_hd__nand3b_1
XFILLER_195_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22485_ _22485_/A vssd1 vssd1 vccd1 vccd1 _22738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21436_ _21294_/C _21434_/Y _21433_/Y _21432_/X vssd1 vssd1 vccd1 vccd1 _21437_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17115__A1 _16976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20307__A _20432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20655__D1 _20454_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21367_ _21367_/A _21367_/B _21367_/C vssd1 vssd1 vccd1 vccd1 _21449_/A sky130_fd_sc_hd__nand3_2
XFILLER_163_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14305__A _14305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17319__C _17520_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20318_ _20311_/A _20311_/B _20311_/C _20562_/A _20317_/B vssd1 vssd1 vccd1 vccd1
+ _20441_/A sky130_fd_sc_hd__a32o_2
XFILLER_162_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21298_ _21419_/A _21276_/C _21264_/Y vssd1 vssd1 vccd1 vccd1 _21415_/A sky130_fd_sc_hd__a21oi_4
XFILLER_150_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20249_ _20249_/A _20249_/B _20249_/C vssd1 vssd1 vccd1 vccd1 _20249_/Y sky130_fd_sc_hd__nand3_1
XFILLER_118_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22882__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15429__A1 _15427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20973__A2 _21083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11664__A _18459_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14810_ _13820_/X _13821_/Y _14624_/A _13823_/Y vssd1 vssd1 vccd1 vccd1 _14810_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _20359_/A vssd1 vssd1 vccd1 vccd1 _15792_/A sky130_fd_sc_hd__buf_2
XFILLER_92_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A wb_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ _14745_/B _14745_/C vssd1 vssd1 vccd1 vccd1 _14741_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16929__A1 _16930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _16447_/A vssd1 vssd1 vccd1 vccd1 _16912_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20725__A2 _17643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _17460_/A vssd1 vssd1 vccd1 vccd1 _17981_/D sky130_fd_sc_hd__buf_2
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _13814_/A _13814_/B _14670_/A vssd1 vssd1 vccd1 vccd1 _14672_/X sky130_fd_sc_hd__a21o_1
XFILLER_72_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11884_ _11895_/C _11894_/A _11894_/B _11895_/B vssd1 vssd1 vccd1 vccd1 _11886_/B
+ sky130_fd_sc_hd__nand4_1
X_16411_ _16206_/X _15879_/X _16210_/Y vssd1 vssd1 vccd1 vccd1 _16412_/B sky130_fd_sc_hd__o21a_1
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13623_ _13623_/A _21498_/B vssd1 vssd1 vccd1 vccd1 _13624_/B sky130_fd_sc_hd__nand2_1
X_17391_ _17391_/A vssd1 vssd1 vccd1 vccd1 _17822_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_73_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12495__A _12532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19130_ _19147_/A _19130_/B vssd1 vssd1 vccd1 vccd1 _19131_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16342_ _16342_/A _16342_/B _16342_/C vssd1 vssd1 vccd1 vccd1 _16369_/A sky130_fd_sc_hd__nand3_4
XFILLER_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _13554_/A vssd1 vssd1 vccd1 vccd1 _13556_/B sky130_fd_sc_hd__inv_2
XFILLER_160_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19061_ _19061_/A _19199_/B _19199_/C vssd1 vssd1 vccd1 vccd1 _19062_/B sky130_fd_sc_hd__and3_1
X_12505_ _12621_/B _12504_/Y _12455_/A vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__o21a_1
X_16273_ _16016_/A _12922_/X _15472_/X _16040_/A _15580_/X vssd1 vssd1 vccd1 vccd1
+ _16273_/X sky130_fd_sc_hd__o32a_1
X_13485_ _13485_/A _13485_/B _13485_/C vssd1 vssd1 vccd1 vccd1 _13556_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12179__B1 _12173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18012_ _18012_/A _18012_/B vssd1 vssd1 vccd1 vccd1 _18053_/B sky130_fd_sc_hd__nand2_1
XFILLER_145_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15224_ _15224_/A _15224_/B _15224_/C _15224_/D vssd1 vssd1 vccd1 vccd1 _15224_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__13915__A1 _13924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12436_ _16778_/A _16779_/A _20466_/B vssd1 vssd1 vccd1 vccd1 _12436_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_154_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21989__A1 _22167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15155_ _15188_/B _15240_/C _15212_/A _14503_/X vssd1 vssd1 vccd1 vccd1 _15155_/X
+ sky130_fd_sc_hd__o22a_1
X_12367_ _22691_/Q _22690_/Q _22688_/Q _12518_/A vssd1 vssd1 vccd1 vccd1 _16323_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14106_ _14184_/B vssd1 vssd1 vccd1 vccd1 _14231_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_114_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11318_ _18690_/B vssd1 vssd1 vccd1 vccd1 _16308_/C sky130_fd_sc_hd__clkbuf_4
X_19963_ _19963_/A _19963_/B vssd1 vssd1 vccd1 vccd1 _19965_/A sky130_fd_sc_hd__nand2_1
XFILLER_153_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15086_ _15086_/A _15086_/B vssd1 vssd1 vccd1 vccd1 _15089_/A sky130_fd_sc_hd__xor2_2
X_12298_ _12424_/C vssd1 vssd1 vccd1 vccd1 _20694_/A sky130_fd_sc_hd__buf_2
XANTENNA__14340__A1 _11430_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17526__A _17634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18914_ _18914_/A _18914_/B _18914_/C vssd1 vssd1 vccd1 vccd1 _18978_/A sky130_fd_sc_hd__nand3_2
XFILLER_141_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14037_ _14035_/A _14523_/A _14035_/B vssd1 vssd1 vccd1 vccd1 _14037_/X sky130_fd_sc_hd__a21o_1
XANTENNA__14340__B2 _13815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19894_ _19894_/A _19921_/A vssd1 vssd1 vccd1 vccd1 _19922_/A sky130_fd_sc_hd__or2_1
XFILLER_164_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14891__A2 _14722_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18845_ _19194_/D vssd1 vssd1 vccd1 vccd1 _19504_/A sky130_fd_sc_hd__buf_2
XFILLER_80_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1069 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18776_ _18768_/A _18768_/B _18768_/C vssd1 vssd1 vccd1 vccd1 _18776_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__21990__B _21990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15988_ _15988_/A _15988_/B _16781_/B vssd1 vssd1 vccd1 vccd1 _15988_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__12103__B1 _16912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14643__A2 _14057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17727_ _17628_/Y _17629_/Y _17682_/Y _17683_/X vssd1 vssd1 vccd1 vccd1 _17727_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19031__A1 _19689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14939_ _14932_/A _14934_/Y _14936_/X vssd1 vssd1 vccd1 vccd1 _14939_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_82_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18357__A _18663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17658_ _17643_/X _17536_/X _17655_/X _17657_/Y vssd1 vssd1 vccd1 vccd1 _17660_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16609_ _15918_/X _17874_/A _17875_/A _16316_/Y _16351_/X vssd1 vssd1 vccd1 vccd1
+ _16609_/X sky130_fd_sc_hd__o32a_1
XFILLER_63_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17589_ _17701_/C _17585_/B _17579_/Y _17583_/Y vssd1 vssd1 vccd1 vccd1 _17590_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12406__B2 _20358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19328_ _19168_/Y _19323_/A _18659_/D _19319_/Y _18896_/C vssd1 vssd1 vccd1 vccd1
+ _19330_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_189_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16308__C _16308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19259_ _19149_/X _19254_/X _19252_/X _19250_/Y vssd1 vssd1 vccd1 vccd1 _19259_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_148_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19619__C _19900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22270_ _22272_/C _22309_/A _22271_/A _22271_/B vssd1 vssd1 vccd1 vccd1 _22273_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_129_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20127__A _20502_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21221_ _13344_/X _13345_/X _13350_/A vssd1 vssd1 vccd1 vccd1 _21237_/A sky130_fd_sc_hd__a21o_1
XANTENNA__18820__A _19061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__A1 _11911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21152_ _22945_/Q _21165_/A _21150_/Y _21151_/X vssd1 vssd1 vccd1 vccd1 _21154_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11468__B _15415_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20103_ _20119_/C _20119_/D vssd1 vssd1 vccd1 vccd1 _20118_/B sky130_fd_sc_hd__nand2_2
XFILLER_160_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17436__A _17436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21083_ _21083_/A _21083_/B _21083_/C vssd1 vssd1 vccd1 vccd1 _21083_/X sky130_fd_sc_hd__and3_1
XFILLER_160_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20034_ _20058_/C _20034_/B vssd1 vssd1 vccd1 vccd1 _20035_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A wb_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19651__A _19651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12299__B _20323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21985_ _21857_/A _21857_/B _21857_/C _21865_/C vssd1 vssd1 vccd1 vccd1 _21986_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18801__A2_N _12171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _20925_/Y _20936_/B _20936_/C _20936_/D vssd1 vssd1 vccd1 vccd1 _20980_/A
+ sky130_fd_sc_hd__nand4b_2
XANTENNA__16387__A2 _15339_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _20864_/Y _20865_/Y _20864_/B _20866_/X _20851_/Y vssd1 vssd1 vccd1 vccd1
+ _20869_/D sky130_fd_sc_hd__o221ai_2
XANTENNA__14937__A3 _14575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19325__A2 _19315_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22606_ _11771_/X input65/X _22608_/S vssd1 vssd1 vccd1 vccd1 _22607_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20798_ _20797_/B _20797_/C _20797_/D _20797_/A vssd1 vssd1 vccd1 vccd1 _20799_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21421__A _21421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12465__D _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22537_ _22537_/A vssd1 vssd1 vccd1 vccd1 _22761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16544__C1 _16496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16515__A _16515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13270_ _22849_/Q vssd1 vssd1 vccd1 vccd1 _13271_/A sky130_fd_sc_hd__inv_2
X_22468_ _22468_/A vssd1 vssd1 vccd1 vccd1 _22730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12221_ _12221_/A _18223_/A vssd1 vssd1 vccd1 vccd1 _12230_/C sky130_fd_sc_hd__xor2_4
XANTENNA__14570__A1 _13973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21419_ _21419_/A _21419_/B _21440_/A _21440_/B vssd1 vssd1 vccd1 vccd1 _21560_/B
+ sky130_fd_sc_hd__nand4_4
X_22399_ _22399_/A vssd1 vssd1 vccd1 vccd1 _22700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12581__B1 _12583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12152_ _12146_/Y _12148_/Y _18099_/A _22794_/Q vssd1 vssd1 vccd1 vccd1 _18339_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16311__A2 _15792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16960_ _16949_/Y _16952_/X _16954_/Y _16959_/Y vssd1 vssd1 vccd1 vccd1 _16978_/B
+ sky130_fd_sc_hd__o211ai_4
X_12083_ _12083_/A _12083_/B vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__nand2_1
XANTENNA__15792__C _15792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22396__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15911_ _15911_/A vssd1 vssd1 vccd1 vccd1 _17407_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16891_ _16890_/X _16672_/X _16889_/C vssd1 vssd1 vccd1 vccd1 _16892_/C sky130_fd_sc_hd__o21bai_1
XANTENNA__15807__D1 _17436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16075__A1 _11845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18630_ _19507_/C vssd1 vssd1 vccd1 vccd1 _19504_/C sky130_fd_sc_hd__buf_2
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _15842_/A _15842_/B vssd1 vssd1 vccd1 vccd1 _15944_/C sky130_fd_sc_hd__nor2_1
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22398__S _22402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14086__B1 _14191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _18561_/A _18561_/B _18561_/C vssd1 vssd1 vccd1 vccd1 _18568_/C sky130_fd_sc_hd__nand3_2
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _16209_/A _15773_/B vssd1 vssd1 vccd1 vccd1 _16208_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12097__C1 _15559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ _15799_/B vssd1 vssd1 vccd1 vccd1 _20452_/B sky130_fd_sc_hd__buf_2
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17512_ _17344_/Y _17347_/Y _17351_/Y vssd1 vssd1 vccd1 vccd1 _17513_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__17024__B1 _17023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _14727_/A _14727_/B _14727_/C _15061_/A vssd1 vssd1 vccd1 vccd1 _14726_/C
+ sky130_fd_sc_hd__nand4_2
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ _18492_/A vssd1 vssd1 vccd1 vccd1 _18493_/A sky130_fd_sc_hd__clkbuf_2
X_11936_ _11936_/A _18093_/D _11936_/C _18093_/C vssd1 vssd1 vccd1 vccd1 _11936_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17443_ _17443_/A vssd1 vssd1 vccd1 vccd1 _17444_/A sky130_fd_sc_hd__buf_2
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14655_ _14655_/A _14655_/B vssd1 vssd1 vccd1 vccd1 _14655_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _19154_/C vssd1 vssd1 vccd1 vccd1 _16106_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_177_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ _13566_/X _13599_/Y _13602_/Y _13605_/Y vssd1 vssd1 vccd1 vccd1 _13608_/B
+ sky130_fd_sc_hd__a2bb2oi_1
X_17374_ _17350_/A _17346_/Y _17347_/Y vssd1 vssd1 vccd1 vccd1 _17375_/A sky130_fd_sc_hd__o21ai_4
X_14586_ _14786_/A vssd1 vssd1 vccd1 vccd1 _14785_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11798_ _11541_/A _11639_/A _11791_/X _11789_/X _11976_/A vssd1 vssd1 vccd1 vccd1
+ _11799_/C sky130_fd_sc_hd__o221ai_4
X_19113_ _12064_/X _19941_/A _19983_/B _19043_/X vssd1 vssd1 vccd1 vccd1 _19113_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_41_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16325_ _16325_/A _16325_/B vssd1 vssd1 vccd1 vccd1 _16344_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15338__B1 _16720_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13537_ _13537_/A _13537_/B vssd1 vssd1 vccd1 vccd1 _13538_/C sky130_fd_sc_hd__nand2_1
XFILLER_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17878__A2 _17806_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15889__A1 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19044_ _19045_/A _19065_/A _19043_/X _18814_/X vssd1 vssd1 vccd1 vccd1 _19044_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__15889__B2 _15888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16256_ _16256_/A _16256_/B _16256_/C _16256_/D vssd1 vssd1 vccd1 vccd1 _16256_/Y
+ sky130_fd_sc_hd__nand4_4
X_13468_ _13468_/A _13468_/B _13468_/C vssd1 vssd1 vccd1 vccd1 _13469_/A sky130_fd_sc_hd__nand3_1
XANTENNA__16550__A2 _15617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15207_ _15207_/A vssd1 vssd1 vccd1 vccd1 _22683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12419_ _12577_/A _12576_/A _12578_/A vssd1 vssd1 vccd1 vccd1 _15335_/A sky130_fd_sc_hd__o21ai_4
XFILLER_154_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16187_ _16145_/Y _16148_/Y _16185_/Y _16186_/Y vssd1 vssd1 vccd1 vccd1 _16187_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_127_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13399_ _13399_/A _13399_/B _13399_/C vssd1 vssd1 vccd1 vccd1 _13495_/B sky130_fd_sc_hd__nand3_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15138_ _15089_/B _15089_/A _15095_/B _15135_/B vssd1 vssd1 vccd1 vccd1 _15139_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19455__B _19945_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19946_ _19946_/A _19946_/B _19946_/C vssd1 vssd1 vccd1 vccd1 _19948_/A sky130_fd_sc_hd__nand3_1
X_15069_ _15069_/A vssd1 vssd1 vccd1 vccd1 _15152_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22387__A1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold22_A hold22/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19877_ _19881_/C _19881_/B _19881_/A vssd1 vssd1 vccd1 vccd1 _19878_/B sky130_fd_sc_hd__nand3b_1
XFILLER_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18828_ _18828_/A vssd1 vssd1 vccd1 vccd1 _18830_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15813__A1 _15631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12627__A1 _15586_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18759_ _18757_/X _18758_/Y _18754_/X _18764_/B vssd1 vssd1 vccd1 vccd1 _18762_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19621__D _19793_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15504__A _16178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_552 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21770_ _21604_/A _21604_/B _21604_/C _21769_/Y vssd1 vssd1 vccd1 vccd1 _21770_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_24_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17566__A1 _11821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20721_ _20721_/A _20721_/B _20721_/C vssd1 vssd1 vccd1 vccd1 _20812_/A sky130_fd_sc_hd__nand3_2
XFILLER_196_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20652_ _20652_/A _20652_/B _20652_/C vssd1 vssd1 vccd1 vccd1 _20652_/Y sky130_fd_sc_hd__nand3_2
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18515__B1 _18680_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20583_ _12968_/A _16611_/A _20577_/B vssd1 vssd1 vccd1 vccd1 _20695_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__20322__B1 _20608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22322_ _22323_/A _22323_/B _22685_/Q vssd1 vssd1 vccd1 vccd1 _22324_/A sky130_fd_sc_hd__a21oi_1
XFILLER_164_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16054__B _18984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11479__A _15633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22253_ _22253_/A _22253_/B vssd1 vssd1 vccd1 vccd1 _22940_/D sky130_fd_sc_hd__xor2_1
XFILLER_191_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21204_ _21201_/Y _21202_/Y _21203_/X vssd1 vssd1 vccd1 vccd1 _21204_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_191_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19491__A1 _19687_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18294__A2 _17635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15893__B _15901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22184_ _22184_/A vssd1 vssd1 vccd1 vccd1 _22265_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_160_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21135_ _21135_/A _21135_/B vssd1 vssd1 vccd1 vccd1 _21135_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22378__A1 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21066_ _21066_/A vssd1 vssd1 vccd1 vccd1 _21066_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16057__A1 _11912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20017_ _18030_/A _18029_/D _19901_/B _19901_/C _19985_/X vssd1 vssd1 vccd1 vccd1
+ _20018_/B sky130_fd_sc_hd__a41oi_4
XFILLER_150_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16462__D1 _20608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22920__CLK _22922_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11942__A _11942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15414__A _20092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _13024_/A _20390_/B _12769_/Y _12645_/A vssd1 vssd1 vccd1 vccd1 _12886_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_161_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21968_ _21972_/A vssd1 vssd1 vccd1 vccd1 _21968_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22550__A1 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _15481_/A _16226_/C _11721_/C vssd1 vssd1 vccd1 vccd1 _11750_/A sky130_fd_sc_hd__nand3b_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ _20919_/A _20919_/B vssd1 vssd1 vccd1 vccd1 _20920_/C sky130_fd_sc_hd__nand2_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21899_ _21899_/A _21899_/B _21899_/C _21899_/D vssd1 vssd1 vccd1 vccd1 _21909_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14440_/A vssd1 vssd1 vccd1 vccd1 _22952_/D sky130_fd_sc_hd__clkbuf_2
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11652_ _15476_/A vssd1 vssd1 vccd1 vccd1 _15694_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14371_ _22733_/Q vssd1 vssd1 vccd1 vccd1 _21580_/B sky130_fd_sc_hd__clkbuf_2
X_11583_ _18663_/A _11583_/B _16313_/C _18875_/C vssd1 vssd1 vccd1 vccd1 _11583_/Y
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12773__A _12773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16110_ _16160_/A _16110_/B _16166_/B vssd1 vssd1 vccd1 vccd1 _16111_/B sky130_fd_sc_hd__and3_1
XFILLER_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13322_ _13322_/A _13322_/B vssd1 vssd1 vccd1 vccd1 _13322_/Y sky130_fd_sc_hd__nand2_1
XFILLER_195_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17090_ _17081_/Y _17084_/X _16997_/C _17006_/A vssd1 vssd1 vccd1 vccd1 _17094_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16041_ _15936_/X _15932_/X _20728_/B _15935_/X _16414_/B vssd1 vssd1 vccd1 vccd1
+ _16041_/X sky130_fd_sc_hd__o41a_1
XANTENNA__11389__A _18482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13253_ _21724_/C _21250_/C _21250_/A _21629_/B _13259_/A vssd1 vssd1 vccd1 vccd1
+ _13262_/A sky130_fd_sc_hd__a32o_1
XFILLER_182_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20616__A1 _20241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12204_ _18203_/B vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18285__A2 _11308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17088__A3 _16997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13184_ _13161_/A _13234_/C _13112_/D vssd1 vssd1 vccd1 vccd1 _13185_/B sky130_fd_sc_hd__a21o_1
XANTENNA__16296__A1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19800_ _19860_/A _19798_/C _19799_/Y _19719_/X vssd1 vssd1 vccd1 vccd1 _19865_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_124_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12135_ _12135_/A _12135_/B vssd1 vssd1 vccd1 vccd1 _18655_/A sky130_fd_sc_hd__nand2_1
X_17992_ _18062_/D _18062_/C _18061_/A _18061_/B vssd1 vssd1 vccd1 vccd1 _17994_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19731_ _19731_/A _19731_/B _19726_/A vssd1 vssd1 vccd1 vccd1 _19731_/Y sky130_fd_sc_hd__nor3b_1
X_16943_ _18193_/A vssd1 vssd1 vccd1 vccd1 _19199_/C sky130_fd_sc_hd__buf_2
X_12066_ _16106_/B vssd1 vssd1 vccd1 vccd1 _17006_/D sky130_fd_sc_hd__buf_4
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11340__B1_N _11334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19662_ _19271_/Y _19268_/Y _19130_/B _19147_/A _19274_/Y vssd1 vssd1 vccd1 vccd1
+ _19664_/B sky130_fd_sc_hd__o2111a_1
X_16874_ _16874_/A _16874_/B _16874_/C vssd1 vssd1 vccd1 vccd1 _16885_/B sky130_fd_sc_hd__nand3_2
XFILLER_64_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18613_ _18613_/A _18613_/B vssd1 vssd1 vccd1 vccd1 _18618_/B sky130_fd_sc_hd__nand2_1
X_15825_ _15825_/A _15825_/B _15825_/C vssd1 vssd1 vccd1 vccd1 _15826_/C sky130_fd_sc_hd__nand3_2
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17523__B _17523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19593_ _17730_/A _19176_/X _19596_/C _19596_/B vssd1 vssd1 vccd1 vccd1 _19594_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12948__A _15991_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _15842_/A _15756_/B _15756_/C vssd1 vssd1 vccd1 vccd1 _15756_/X sky130_fd_sc_hd__and3_2
X_18544_ _11979_/Y _11980_/X _12111_/X _16276_/A _11474_/X vssd1 vssd1 vccd1 vccd1
+ _18544_/X sky130_fd_sc_hd__o32a_1
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17548__A1 _17731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12968_ _12968_/A _12968_/B _20697_/A _12968_/D vssd1 vssd1 vccd1 vccd1 _12989_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_92_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22541__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14707_ _14494_/C _14951_/A _14815_/C _14708_/D vssd1 vssd1 vccd1 vccd1 _14711_/C
+ sky130_fd_sc_hd__a22o_1
X_18475_ _18471_/X _18472_/X _18473_/Y _18474_/Y vssd1 vssd1 vccd1 vccd1 _18478_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__17012__A3 _16723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _11606_/X _11914_/Y _11918_/Y vssd1 vssd1 vccd1 vccd1 _11924_/C sky130_fd_sc_hd__o21ai_1
X_15687_ _15676_/C _15676_/D _15686_/Y vssd1 vssd1 vccd1 vccd1 _15687_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12899_ _12898_/A _12898_/B _12665_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _12900_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _17426_/A _20854_/B _20854_/A _19614_/A vssd1 vssd1 vccd1 vccd1 _17431_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ _14650_/A _14740_/B _14650_/C vssd1 vssd1 vccd1 vccd1 _14638_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17357_ _17226_/X _17227_/X _17228_/Y _17215_/Y vssd1 vssd1 vccd1 vccd1 _17357_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13779__A _22873_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16508__C1 _16496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14569_ _14468_/B _14685_/A _14568_/Y vssd1 vssd1 vccd1 vccd1 _14575_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__16155__A _16155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16308_ _20608_/B _20608_/C _16308_/C vssd1 vssd1 vccd1 vccd1 _16308_/X sky130_fd_sc_hd__and3_1
XANTENNA__20855__A1 _20514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17288_ _17288_/A _17288_/B vssd1 vssd1 vccd1 vccd1 _17290_/B sky130_fd_sc_hd__nand2_1
XFILLER_147_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19027_ _18158_/X _19023_/X _19024_/Y _19026_/Y vssd1 vssd1 vccd1 vccd1 _19037_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_174_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16239_ _16504_/A vssd1 vssd1 vccd1 vccd1 _16530_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_118_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16602__B _16602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19929_ _19293_/X _19294_/X _19878_/Y _19880_/Y _19926_/A vssd1 vssd1 vccd1 vccd1
+ _19970_/C sky130_fd_sc_hd__o221ai_4
XANTENNA__22943__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22940_ _22943_/CLK _22940_/D vssd1 vssd1 vccd1 vccd1 _22940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22871_ _22915_/CLK _22871_/D vssd1 vssd1 vccd1 vccd1 _22871_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11762__A _11762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21822_ _21700_/X _21701_/X _21815_/B _21702_/B vssd1 vssd1 vccd1 vccd1 _21822_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12076__A2 _11606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22532__A1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21753_ _21589_/Y _21753_/B _21753_/C vssd1 vssd1 vccd1 vccd1 _21760_/A sky130_fd_sc_hd__nand3b_1
XFILLER_19_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20704_ _20704_/A _20704_/B vssd1 vssd1 vccd1 vccd1 _20704_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21684_ _21399_/B _22229_/B _21399_/A _21547_/A vssd1 vssd1 vccd1 vccd1 _21684_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__14773__A1 _14362_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13576__A2 _13126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20635_ _20738_/A _20738_/B _20738_/C vssd1 vssd1 vccd1 vccd1 _20737_/A sky130_fd_sc_hd__nand3_4
XANTENNA__16065__A _18130_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20846__A1 _16585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20566_ _20566_/A _20566_/B vssd1 vssd1 vccd1 vccd1 _20566_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22305_ _22306_/C _22306_/A _22265_/B _22263_/B vssd1 vssd1 vccd1 vccd1 _22307_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20497_ _20493_/X _20581_/B _20495_/Y _20496_/Y vssd1 vssd1 vccd1 vccd1 _20629_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_164_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12536__B1 _16759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22236_ _22193_/B _22178_/B _22238_/B _22219_/Y vssd1 vssd1 vccd1 vccd1 _22237_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16278__B2 _16277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20074__A2 _20429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22167_ _22167_/A vssd1 vssd1 vccd1 vccd1 _22306_/B sky130_fd_sc_hd__buf_2
XFILLER_191_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14313__A _14351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21118_ _21118_/A _21135_/A _21118_/C vssd1 vssd1 vccd1 vccd1 _21119_/B sky130_fd_sc_hd__and3_1
X_22098_ _21330_/A _21330_/B _21269_/A vssd1 vssd1 vccd1 vccd1 _22098_/X sky130_fd_sc_hd__a21o_1
XFILLER_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19767__A2 _17822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13940_ _13975_/D vssd1 vssd1 vccd1 vccd1 _14210_/A sky130_fd_sc_hd__buf_2
XFILLER_47_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_912 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21049_ _21017_/C _17839_/B _17839_/C _21046_/B vssd1 vssd1 vccd1 vccd1 _21050_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15789__B1 _16058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ _13875_/A _13989_/A _14722_/C vssd1 vssd1 vccd1 vccd1 _13881_/B sky130_fd_sc_hd__nand3_1
XFILLER_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11672__A _11672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15610_ _20463_/A _20463_/B vssd1 vssd1 vccd1 vccd1 _15611_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12822_ _12822_/A _12822_/B _16323_/C vssd1 vssd1 vccd1 vccd1 _12823_/A sky130_fd_sc_hd__nand3_2
X_16590_ _16585_/A _16585_/B _15918_/A vssd1 vssd1 vccd1 vccd1 _16590_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12067__A2 _18830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22523__A1 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15541_ _15548_/B vssd1 vssd1 vccd1 vccd1 _15541_/X sky130_fd_sc_hd__buf_4
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12753_ _12895_/A _12895_/B _12895_/C vssd1 vssd1 vccd1 vccd1 _13044_/C sky130_fd_sc_hd__and3_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _18589_/A _18590_/A vssd1 vssd1 vccd1 vccd1 _18600_/A sky130_fd_sc_hd__or2_1
X_11704_ _11737_/A vssd1 vssd1 vccd1 vccd1 _11704_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15472_ _15472_/A vssd1 vssd1 vccd1 vccd1 _15472_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_588 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12684_ _20593_/D vssd1 vssd1 vccd1 vccd1 _20793_/B sky130_fd_sc_hd__buf_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17603_/B _17079_/Y _17213_/C vssd1 vssd1 vccd1 vccd1 _17370_/A sky130_fd_sc_hd__o21bai_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _22813_/Q _14411_/X _14412_/X _14413_/X _22781_/Q vssd1 vssd1 vccd1 vccd1
+ _14423_/X sky130_fd_sc_hd__a32o_1
X_18191_ _18191_/A vssd1 vssd1 vccd1 vccd1 _18276_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_11635_ _11614_/Y _11623_/X _19043_/A _17083_/A vssd1 vssd1 vccd1 vccd1 _11635_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__22816__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17142_ _17142_/A vssd1 vssd1 vccd1 vccd1 _17142_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12934__C _15696_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14354_ _14354_/A vssd1 vssd1 vccd1 vccd1 _14354_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11566_ _11818_/A vssd1 vssd1 vccd1 vccd1 _11566_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13305_ _13305_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _21207_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17073_ _17073_/A _17073_/B vssd1 vssd1 vccd1 vccd1 _22955_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14285_ _14285_/A _14285_/B _14285_/C vssd1 vssd1 vccd1 vccd1 _14288_/A sky130_fd_sc_hd__nand3_1
XFILLER_155_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12008__A _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11497_ _11420_/A _12148_/B _12146_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11792_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_157_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16024_ _16024_/A _16024_/B _16024_/C vssd1 vssd1 vccd1 vccd1 _16024_/Y sky130_fd_sc_hd__nor3_1
XFILLER_6_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13236_ _13633_/C vssd1 vssd1 vccd1 vccd1 _21259_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16269__B2 _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11847__A _16078_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _13340_/A _13286_/B _13166_/Y vssd1 vssd1 vccd1 vccd1 _13396_/A sky130_fd_sc_hd__a21o_1
XFILLER_124_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19207__A1 _19203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12118_ _12118_/A vssd1 vssd1 vccd1 vccd1 _16016_/A sky130_fd_sc_hd__buf_2
X_17975_ _19896_/B vssd1 vssd1 vccd1 vccd1 _19454_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13098_ _13098_/A vssd1 vssd1 vccd1 vccd1 _14380_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19714_ _17442_/A _19517_/A _16016_/X _19838_/A vssd1 vssd1 vccd1 vccd1 _19714_/X
+ sky130_fd_sc_hd__o22a_1
X_16926_ _16926_/A _16926_/B vssd1 vssd1 vccd1 vccd1 _16926_/Y sky130_fd_sc_hd__nand2_1
X_12049_ _19197_/C vssd1 vssd1 vccd1 vccd1 _19490_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19645_ _19640_/X _19641_/X _19642_/X _19540_/Y _19644_/Y vssd1 vssd1 vccd1 vccd1
+ _19740_/A sky130_fd_sc_hd__o2111ai_4
X_16857_ _16594_/B _16594_/C _16594_/A _16601_/Y vssd1 vssd1 vccd1 vccd1 _16858_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12678__A _16256_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11582__A _18690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15808_ _15808_/A vssd1 vssd1 vccd1 vccd1 _15808_/X sky130_fd_sc_hd__buf_4
X_19576_ _19427_/C _19437_/Y _19439_/A _19439_/B _19565_/Y vssd1 vssd1 vccd1 vccd1
+ _19682_/A sky130_fd_sc_hd__a221o_1
X_16788_ _15530_/A _15531_/A _12294_/A _12294_/B vssd1 vssd1 vccd1 vccd1 _16788_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14452__B1 _14448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16992__A2 _11505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15739_ _15860_/B _15766_/A vssd1 vssd1 vccd1 vccd1 _15758_/B sky130_fd_sc_hd__nand2_1
X_18527_ _18527_/A _18527_/B _18527_/C vssd1 vssd1 vccd1 vccd1 _18527_/Y sky130_fd_sc_hd__nand3_2
XFILLER_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18194__A1 _11502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18194__B2 _17381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18458_ _18458_/A _18458_/B _18458_/C vssd1 vssd1 vccd1 vccd1 _18462_/A sky130_fd_sc_hd__nand3_1
XFILLER_179_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17409_ _17402_/Y _17404_/X _17390_/Y _17408_/Y vssd1 vssd1 vccd1 vccd1 _17410_/A
+ sky130_fd_sc_hd__o211ai_1
X_18389_ _18389_/A _18389_/B _18389_/C vssd1 vssd1 vccd1 vccd1 _18389_/X sky130_fd_sc_hd__and3_1
XFILLER_159_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20420_ _20420_/A _20545_/A _20420_/C vssd1 vssd1 vccd1 vccd1 _20423_/B sky130_fd_sc_hd__nand3_2
XFILLER_174_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13659__D _21938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14117__B _14785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20351_ _20343_/A _20464_/A _20347_/B _20339_/Y vssd1 vssd1 vccd1 vccd1 _20353_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_174_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20282_ _20269_/X _20274_/Y _20280_/Y _20281_/X vssd1 vssd1 vccd1 vccd1 _20286_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_127_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19346__D _19504_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22021_ _22021_/A _22021_/B vssd1 vssd1 vccd1 vccd1 _22936_/D sky130_fd_sc_hd__xor2_1
XANTENNA__11741__A1 _18203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17444__A _17444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18259__B _18259_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22923_ _22948_/CLK _22923_/D vssd1 vssd1 vccd1 vccd1 _22923_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22854_ _22943_/CLK _22866_/Q vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15899__A _16308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21805_ _21651_/X _21805_/B _22231_/D _21805_/D vssd1 vssd1 vccd1 vccd1 _21805_/X
+ sky130_fd_sc_hd__and4b_2
XANTENNA__14994__A1 _15004_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14994__B2 _15050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22785_ _22787_/CLK _22785_/D vssd1 vssd1 vccd1 vccd1 _22785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15114__D _15114_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22839__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21736_ _21790_/A vssd1 vssd1 vccd1 vccd1 _21736_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16735__A2 _15935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21667_ _21269_/A _13343_/X _21514_/C _21666_/Y vssd1 vssd1 vccd1 vccd1 _21667_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14308__A _14370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11420_ _11420_/A _11420_/B _11420_/C _11420_/D vssd1 vssd1 vccd1 vccd1 _11428_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20618_ _17407_/A _17131_/B _20917_/A _20504_/X vssd1 vssd1 vccd1 vccd1 _20620_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21598_ _21771_/A _21771_/B _21771_/C vssd1 vssd1 vccd1 vccd1 _21645_/A sky130_fd_sc_hd__nand3_2
XFILLER_153_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ _12090_/B vssd1 vssd1 vccd1 vccd1 _11351_/X sky130_fd_sc_hd__buf_2
XANTENNA__18893__C1 _17313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20549_ _20549_/A _20549_/B _20549_/C _20549_/D vssd1 vssd1 vccd1 vccd1 _20549_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_165_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14070_ _13857_/X _13725_/Y _14184_/C _13728_/A vssd1 vssd1 vccd1 vccd1 _14085_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__17338__B _17338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11282_ _11306_/A _11421_/A vssd1 vssd1 vccd1 vccd1 _11860_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11667__A _15435_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17448__B1 _16124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ _20697_/A vssd1 vssd1 vccd1 vccd1 _13022_/B sky130_fd_sc_hd__clkbuf_4
X_22219_ _22219_/A _22219_/B vssd1 vssd1 vccd1 vccd1 _22219_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input44_A wb_dat_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18660__A2 _19320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17760_ _17760_/A _17760_/B _17760_/C vssd1 vssd1 vccd1 vccd1 _17761_/C sky130_fd_sc_hd__nand3_1
X_14972_ _14972_/A _14972_/B vssd1 vssd1 vccd1 vccd1 _14972_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19272__C _19272_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12142__D1 _15357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16711_ _17281_/B _20593_/A _16711_/C _17312_/A vssd1 vssd1 vccd1 vccd1 _16711_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13923_ _13923_/A vssd1 vssd1 vccd1 vccd1 _13923_/X sky130_fd_sc_hd__clkbuf_2
X_17691_ _17626_/B _17626_/A _17627_/X _17697_/B _17697_/C vssd1 vssd1 vccd1 vccd1
+ _17693_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19430_ _18958_/B _19132_/Y _19429_/Y vssd1 vssd1 vccd1 vccd1 _19430_/X sky130_fd_sc_hd__a21o_1
X_16642_ _17806_/D vssd1 vssd1 vccd1 vccd1 _17039_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13854_ _13854_/A vssd1 vssd1 vccd1 vccd1 _14061_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_142_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ _12329_/A _12803_/X _12804_/Y _15409_/A vssd1 vssd1 vccd1 vccd1 _12817_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_19361_ _12234_/X _12237_/X _19350_/A vssd1 vssd1 vccd1 vccd1 _19361_/Y sky130_fd_sc_hd__a21oi_1
X_16573_ _20579_/A vssd1 vssd1 vccd1 vccd1 _20584_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ _14079_/A _14489_/B _13765_/X vssd1 vssd1 vccd1 vccd1 _13786_/B sky130_fd_sc_hd__o21ai_1
XFILLER_163_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15524_ _15521_/X _15522_/X _12929_/A _15523_/X vssd1 vssd1 vccd1 vccd1 _15524_/X
+ sky130_fd_sc_hd__a211o_4
X_18312_ _22796_/Q vssd1 vssd1 vccd1 vccd1 _18678_/C sky130_fd_sc_hd__clkinv_2
X_19292_ _19292_/A _19292_/B vssd1 vssd1 vccd1 vccd1 _22896_/D sky130_fd_sc_hd__nor2_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _12734_/X _12735_/X _12950_/C vssd1 vssd1 vccd1 vccd1 _12737_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__17520__C _17520_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12460__A2 _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _18251_/B vssd1 vssd1 vccd1 vccd1 _18257_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15455_ _15455_/A vssd1 vssd1 vccd1 vccd1 _15546_/A sky130_fd_sc_hd__buf_2
XANTENNA__15321__B _16712_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12667_ _12668_/A _12668_/B _12745_/A _12745_/B vssd1 vssd1 vccd1 vccd1 _12741_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14406_ _22807_/Q _14397_/X _14398_/X _14391_/X _22775_/Q vssd1 vssd1 vccd1 vccd1
+ _14406_/X sky130_fd_sc_hd__a32o_1
X_18174_ _18174_/A vssd1 vssd1 vccd1 vccd1 _18404_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11618_ _22790_/Q _12148_/A _12148_/B _12146_/A vssd1 vssd1 vccd1 vccd1 _11619_/A
+ sky130_fd_sc_hd__nand4b_1
X_15386_ _15386_/A vssd1 vssd1 vccd1 vccd1 _15517_/A sky130_fd_sc_hd__buf_2
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12598_ _12598_/A vssd1 vssd1 vccd1 vccd1 _15450_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_129_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17125_ _16926_/B _16915_/Y _16913_/X _16911_/X vssd1 vssd1 vccd1 vccd1 _17125_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_144_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21483__A1 _13050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14337_ _14351_/A vssd1 vssd1 vccd1 vccd1 _14337_/X sky130_fd_sc_hd__clkbuf_2
X_11549_ _11401_/Y _11895_/A _11895_/B _11547_/Y _11548_/X vssd1 vssd1 vccd1 vccd1
+ _11840_/A sky130_fd_sc_hd__o2111ai_2
XFILLER_128_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11971__A1 _15904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17056_ _17076_/C _17053_/Y _17048_/Y _16659_/B vssd1 vssd1 vccd1 vccd1 _17058_/A
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_7_595 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14268_ _14269_/A _14279_/A _14269_/C _14269_/D vssd1 vssd1 vccd1 vccd1 _14280_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16007_ _16045_/A _16045_/B _16045_/C vssd1 vssd1 vccd1 vccd1 _16007_/X sky130_fd_sc_hd__and3_1
XFILLER_83_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13219_ _21362_/A vssd1 vssd1 vccd1 vccd1 _21638_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_152_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _14199_/A _14684_/B vssd1 vssd1 vccd1 vccd1 _14259_/B sky130_fd_sc_hd__nand2_2
XFILLER_112_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15991__B _15991_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18651__A2 _16275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17958_ _17958_/A _17958_/B vssd1 vssd1 vccd1 vccd1 _18002_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16909_ _16830_/Y _16831_/X _16834_/A vssd1 vssd1 vccd1 vccd1 _16909_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17889_ _17889_/A _17889_/B vssd1 vssd1 vccd1 vccd1 _17891_/A sky130_fd_sc_hd__xnor2_1
XFILLER_93_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19628_ _19709_/C _19629_/B _19636_/B vssd1 vssd1 vccd1 vccd1 _19634_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19559_ _19549_/Y _19545_/Y _19553_/X vssd1 vssd1 vccd1 vccd1 _19559_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12987__B1 _20793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22570_ _22570_/A vssd1 vssd1 vccd1 vccd1 _22776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21521_ _21519_/X _21520_/Y _21374_/A vssd1 vssd1 vccd1 vccd1 _21522_/B sky130_fd_sc_hd__o21ai_1
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21452_ _21365_/B _21633_/A _21632_/A _21805_/B _21449_/Y vssd1 vssd1 vccd1 vccd1
+ _21460_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20403_ _20403_/A _20403_/B _20403_/C vssd1 vssd1 vccd1 vccd1 _20403_/X sky130_fd_sc_hd__and3_1
XANTENNA__17439__A _17732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21383_ _21383_/A vssd1 vssd1 vccd1 vccd1 _21383_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11962__A1 _11751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20334_ _20335_/A _20335_/B _20335_/C vssd1 vssd1 vccd1 vccd1 _20336_/A sky130_fd_sc_hd__a21oi_1
XFILLER_162_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21226__A1 _22057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18627__C1 _18626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20265_ _20397_/A _20266_/A _20260_/Y _20264_/Y vssd1 vssd1 vccd1 vccd1 _20268_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_163_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22004_ _21997_/Y _22002_/Y _21999_/Y _22003_/X vssd1 vssd1 vccd1 vccd1 _22008_/D
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12911__B1 _16498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20196_ _20195_/Y _20065_/Y _20189_/B _20189_/C vssd1 vssd1 vccd1 vccd1 _20309_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_89_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15456__A2 _15546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15310__D1 _15774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14948__D _15115_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22906_ _22949_/CLK _22906_/D vssd1 vssd1 vccd1 vccd1 _22906_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_1_1_0_bq_clk_i_A clkbuf_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12111__A _12111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14416__B1 _14413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12690__A2 _20793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22837_ _22929_/CLK _22849_/Q vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11950__A _12003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12978__B1 _12968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15422__A _16477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _21739_/B vssd1 vssd1 vccd1 vccd1 _21866_/C sky130_fd_sc_hd__clkbuf_4
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22768_ _22768_/CLK _22768_/D vssd1 vssd1 vccd1 vccd1 _22768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20504__A3 _15341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14719__A1 _13851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ _12550_/C _12549_/A vssd1 vssd1 vccd1 vccd1 _12522_/B sky130_fd_sc_hd__nand2_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21719_ _21719_/A _21719_/B vssd1 vssd1 vccd1 vccd1 _21721_/A sky130_fd_sc_hd__nor2_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22699_ _22701_/CLK _22699_/D vssd1 vssd1 vccd1 vccd1 _22699_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15240_/A _15240_/B _15240_/C _15240_/D vssd1 vssd1 vccd1 vccd1 _15241_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_36_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12452_ _15314_/A vssd1 vssd1 vccd1 vccd1 _20323_/B sky130_fd_sc_hd__buf_4
XFILLER_138_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11403_ _11512_/A vssd1 vssd1 vccd1 vccd1 _18292_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_184_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15171_ _15171_/A _15171_/B vssd1 vssd1 vccd1 vccd1 _15173_/C sky130_fd_sc_hd__and2_1
X_12383_ _15352_/A _12383_/B _20207_/C vssd1 vssd1 vccd1 vccd1 _12487_/C sky130_fd_sc_hd__nand3_2
XFILLER_125_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20673__C1 _17386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14122_ _14122_/A vssd1 vssd1 vccd1 vccd1 _14274_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11334_ _11404_/B vssd1 vssd1 vccd1 vccd1 _11334_/X sky130_fd_sc_hd__buf_2
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15695__A2 _15309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11397__A _11968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18930_ _18978_/A _18931_/B _18977_/B vssd1 vssd1 vccd1 vccd1 _18932_/B sky130_fd_sc_hd__a21o_1
X_14053_ _14052_/C _14052_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14094_/C sky130_fd_sc_hd__a21o_1
XFILLER_98_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ _13004_/A _13004_/B _13004_/C vssd1 vssd1 vccd1 vccd1 _13006_/A sky130_fd_sc_hd__nand3_1
X_18861_ _18861_/A _18861_/B vssd1 vssd1 vccd1 vccd1 _18863_/A sky130_fd_sc_hd__nand2_1
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17841__B1 _19793_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17812_ _17812_/A _17895_/B vssd1 vssd1 vccd1 vccd1 _17827_/A sky130_fd_sc_hd__and2_1
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18792_ _18792_/A _18792_/B vssd1 vssd1 vccd1 vccd1 _22893_/D sky130_fd_sc_hd__xnor2_1
XFILLER_43_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17743_ _17882_/C _18305_/C _17826_/A _17743_/D vssd1 vssd1 vccd1 vccd1 _17826_/B
+ sky130_fd_sc_hd__nand4_2
X_14955_ _14955_/A _14955_/B vssd1 vssd1 vccd1 vccd1 _14955_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13117__A _22841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13906_ _13897_/Y _13745_/C _22761_/Q vssd1 vssd1 vccd1 vccd1 _14465_/A sky130_fd_sc_hd__a21o_2
X_17674_ _19619_/D _21083_/A _21083_/B _19793_/C _17431_/C vssd1 vssd1 vccd1 vccd1
+ _17678_/B sky130_fd_sc_hd__a32o_1
X_14886_ _14881_/A _14952_/B _14879_/Y _14880_/X vssd1 vssd1 vccd1 vccd1 _14886_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_63_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19413_ _19244_/Y _19400_/X _19407_/X _19408_/X vssd1 vssd1 vccd1 vccd1 _19413_/X
+ sky130_fd_sc_hd__o211a_1
X_16625_ _16625_/A _16625_/B _16625_/C vssd1 vssd1 vccd1 vccd1 _16637_/B sky130_fd_sc_hd__nand3_2
X_13837_ _13837_/A _13865_/A vssd1 vssd1 vccd1 vccd1 _13837_/Y sky130_fd_sc_hd__nand2_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19344_ _19530_/A _19530_/C _19530_/D vssd1 vssd1 vccd1 vccd1 _19344_/Y sky130_fd_sc_hd__nand3_1
X_16556_ _16098_/A _17111_/A _16295_/Y _16550_/Y _16552_/Y vssd1 vssd1 vccd1 vccd1
+ _16557_/C sky130_fd_sc_hd__o221ai_4
XFILLER_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13768_ _13707_/A _13776_/B _13745_/C _13761_/B vssd1 vssd1 vccd1 vccd1 _14110_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_31_620 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22350__C1 _22352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15507_ _15580_/A _12735_/X _15449_/X _15452_/Y vssd1 vssd1 vccd1 vccd1 _15507_/X
+ sky130_fd_sc_hd__o31a_1
X_12719_ _12719_/A vssd1 vssd1 vccd1 vccd1 _12968_/D sky130_fd_sc_hd__buf_2
X_19275_ _19268_/Y _19271_/Y _19274_/Y vssd1 vssd1 vccd1 vccd1 _19295_/A sky130_fd_sc_hd__o21ai_1
X_16487_ _16100_/D _16491_/B _16964_/A _15810_/C _16231_/X vssd1 vssd1 vccd1 vccd1
+ _16493_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13699_ _14506_/B vssd1 vssd1 vccd1 vccd1 _14808_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15438_ _16473_/A _16473_/B _16488_/A vssd1 vssd1 vccd1 vccd1 _15439_/A sky130_fd_sc_hd__nand3_2
X_18226_ _18275_/A _18275_/B _18226_/C vssd1 vssd1 vccd1 vccd1 _18226_/Y sky130_fd_sc_hd__nand3_1
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14186__A2 _14561_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17109__C1 _11666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20259__A2 _20261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18157_ _11904_/A _11905_/A _19165_/A _19168_/C vssd1 vssd1 vccd1 vccd1 _18995_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_50_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _15369_/A _15369_/B _15369_/C vssd1 vssd1 vccd1 vccd1 _17423_/A sky130_fd_sc_hd__nand3_2
XANTENNA__13933__A2 _13949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17108_ _19012_/D _17108_/B _20593_/A _17672_/A vssd1 vssd1 vccd1 vccd1 _17116_/A
+ sky130_fd_sc_hd__nand4_4
XANTENNA__11944__B2 _11774_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18088_ _22910_/Q vssd1 vssd1 vccd1 vccd1 _18088_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22405__A0 _20069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17039_ _17039_/A _17840_/A _17039_/C _17039_/D vssd1 vssd1 vccd1 vccd1 _17040_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16883__B2 _16644_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20050_ _20049_/C _20049_/B _20049_/A vssd1 vssd1 vccd1 vccd1 _20051_/B sky130_fd_sc_hd__a21oi_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22684__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater132 _22696_/CLK vssd1 vssd1 vccd1 vccd1 _22701_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater143 _22803_/CLK vssd1 vssd1 vccd1 vccd1 _22815_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater154 _22747_/CLK vssd1 vssd1 vccd1 vccd1 _22749_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater165 _22768_/CLK vssd1 vssd1 vccd1 vccd1 _22801_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16399__B1 _16398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20195__A1 _13045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20952_ _20952_/A vssd1 vssd1 vccd1 vccd1 _20989_/A sky130_fd_sc_hd__inv_2
XFILLER_54_734 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_49 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14162__A2_N _14147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__B1 _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ _20843_/X _20884_/A _15935_/X _20806_/Y _20884_/C vssd1 vssd1 vccd1 vccd1
+ _20887_/C sky130_fd_sc_hd__o311a_1
XFILLER_42_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22622_ _18258_/A input41/X _22630_/S vssd1 vssd1 vccd1 vccd1 _22623_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22553_ _22553_/A vssd1 vssd1 vccd1 vccd1 _22768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17363__A2 _17959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21504_ _21504_/A _21504_/B _21504_/C vssd1 vssd1 vccd1 vccd1 _21508_/A sky130_fd_sc_hd__nand3_1
XFILLER_166_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22484_ _22738_/Q input44/X _22486_/S vssd1 vssd1 vccd1 vccd1 _22485_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_628 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21435_ _21432_/X _21433_/Y _21434_/Y _21294_/C vssd1 vssd1 vccd1 vccd1 _21437_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_5_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21366_ _21632_/A _21177_/A _21372_/A _21372_/B vssd1 vssd1 vccd1 vccd1 _21369_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17319__D _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20317_ _20317_/A _20317_/B vssd1 vssd1 vccd1 vccd1 _22911_/D sky130_fd_sc_hd__xor2_4
XFILLER_135_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21297_ _21422_/A _21424_/C _21423_/A vssd1 vssd1 vccd1 vccd1 _21297_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_1_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20248_ _20133_/Y _20247_/Y _20244_/A _20242_/X vssd1 vssd1 vccd1 vccd1 _20249_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20323__A _20323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15429__A2 _15933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17823__B1 _17928_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15417__A _20611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20179_ _12765_/X _20843_/A _12878_/X _12781_/B vssd1 vssd1 vccd1 vccd1 _20179_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20973__A3 _21083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__B _18666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17632__A _17632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14740_ _14740_/A _14740_/B _14740_/C _14740_/D vssd1 vssd1 vccd1 vccd1 _14745_/C
+ sky130_fd_sc_hd__nand4_2
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _11846_/Y _11774_/Y _11951_/Y vssd1 vssd1 vccd1 vccd1 _11952_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16929__A2 _17341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13860__A1 _13930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11871__B1 _19000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14671_ _13930_/A _13930_/B _14516_/C _14522_/C _15213_/A vssd1 vssd1 vccd1 vccd1
+ _14750_/A sky130_fd_sc_hd__a221o_1
XFILLER_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _11883_/A _11883_/B _11883_/C vssd1 vssd1 vccd1 vccd1 _11895_/C sky130_fd_sc_hd__nand3_1
XFILLER_33_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19328__B1 _18659_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16410_ _16408_/Y _16035_/C _16421_/C _16421_/D vssd1 vssd1 vccd1 vccd1 _16657_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11680__A _15484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13622_ _13566_/X _13599_/Y _13602_/Y _13605_/Y vssd1 vssd1 vccd1 vccd1 _13672_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17390_ _17145_/B _17247_/X _17257_/B _17249_/Y vssd1 vssd1 vccd1 vccd1 _17390_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_73_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19879__A1 _19293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16341_ _16354_/A _16617_/A _16354_/C vssd1 vssd1 vccd1 vccd1 _16342_/C sky130_fd_sc_hd__nand3b_1
X_13553_ _13559_/A _13559_/B _13559_/C _13677_/B _13677_/C vssd1 vssd1 vccd1 vccd1
+ _13558_/C sky130_fd_sc_hd__a32oi_4
XFILLER_41_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19060_ _17388_/A _18371_/X _19059_/Y _19051_/X _19055_/Y vssd1 vssd1 vccd1 vccd1
+ _19063_/B sky130_fd_sc_hd__o221ai_4
X_12504_ _12454_/B _12454_/C _12454_/A vssd1 vssd1 vccd1 vccd1 _12504_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16272_ _16272_/A _16272_/B _16272_/C vssd1 vssd1 vccd1 vccd1 _16596_/A sky130_fd_sc_hd__nand3_2
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13484_ _13484_/A _13484_/B _13484_/C vssd1 vssd1 vccd1 vccd1 _13485_/C sky130_fd_sc_hd__nand3_1
XFILLER_186_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18011_ _17970_/Y _18009_/Y _18010_/Y vssd1 vssd1 vccd1 vccd1 _18012_/B sky130_fd_sc_hd__o21ai_1
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12179__B2 _12174_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15223_ _15223_/A _15223_/B vssd1 vssd1 vccd1 vccd1 _15223_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12435_ _22818_/Q vssd1 vssd1 vccd1 vccd1 _20466_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_138_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11926__A1 _11693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21989__A2 _21341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15154_ _15154_/A _15154_/B _15215_/A _15154_/D vssd1 vssd1 vccd1 vccd1 _15154_/X
+ sky130_fd_sc_hd__and4_2
X_12366_ _22689_/Q vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__buf_2
XFILLER_153_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13128__B1 _13126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14105_ _14184_/A vssd1 vssd1 vccd1 vccd1 _14231_/A sky130_fd_sc_hd__clkbuf_2
X_11317_ _11790_/C vssd1 vssd1 vccd1 vccd1 _18690_/B sky130_fd_sc_hd__buf_2
X_19962_ _19962_/A _19962_/B _19962_/C vssd1 vssd1 vccd1 vccd1 _19963_/B sky130_fd_sc_hd__nand3_1
XANTENNA__17807__A _17833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15085_ _15085_/A _15085_/B vssd1 vssd1 vccd1 vccd1 _15086_/B sky130_fd_sc_hd__xor2_2
X_12297_ _12415_/A _12411_/A vssd1 vssd1 vccd1 vccd1 _12424_/C sky130_fd_sc_hd__nor2_1
XANTENNA__16711__A _17281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18913_ _18908_/C _18908_/B _18911_/Y _18912_/X vssd1 vssd1 vccd1 vccd1 _18914_/C
+ sky130_fd_sc_hd__o2bb2ai_2
X_14036_ _14052_/A _14036_/B vssd1 vssd1 vccd1 vccd1 _14036_/Y sky130_fd_sc_hd__nand2_1
X_19893_ _19893_/A _19893_/B _22921_/Q vssd1 vssd1 vccd1 vccd1 _19976_/C sky130_fd_sc_hd__nand3_1
XFILLER_171_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11855__A _18706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18844_ _19470_/D _19161_/A _19587_/B _16062_/A _18862_/B vssd1 vssd1 vccd1 vccd1
+ _18854_/A sky130_fd_sc_hd__a41o_1
XANTENNA__14891__A3 _14722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21048__B _21048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15046__B _15046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18775_ _18772_/Y _18773_/Y _18774_/Y _18774_/D vssd1 vssd1 vccd1 vccd1 _19132_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15987_ _16261_/B vssd1 vssd1 vccd1 vccd1 _17539_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__12103__A1 _11625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20528__A2_N _20381_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17726_ _17790_/D _17790_/C _17726_/C _17726_/D vssd1 vssd1 vccd1 vccd1 _17726_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19031__A2 _19334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14938_ _14996_/D _14934_/Y _14936_/X _14937_/X vssd1 vssd1 vccd1 vccd1 _14945_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18357__B _19322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17657_ _17535_/B _17652_/Y _17648_/Y _18305_/C _17816_/A vssd1 vssd1 vccd1 vccd1
+ _17657_/Y sky130_fd_sc_hd__o2111ai_4
XANTENNA__16158__A _17085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14869_ _14869_/A _14869_/B _14869_/C vssd1 vssd1 vccd1 vccd1 _14871_/A sky130_fd_sc_hd__nand3_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12686__A _22817_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18790__A1 _18432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16608_ _16608_/A vssd1 vssd1 vccd1 vccd1 _16624_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12406__A2 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17588_ _17584_/X _17586_/Y _17590_/B vssd1 vssd1 vccd1 vccd1 _17624_/A sky130_fd_sc_hd__o21bai_1
XFILLER_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19327_ _19317_/Y _19319_/Y _12114_/X _18856_/A vssd1 vssd1 vccd1 vccd1 _19330_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__15997__A _18984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16539_ _16289_/Y _16290_/X _16288_/C vssd1 vssd1 vccd1 vccd1 _16540_/B sky130_fd_sc_hd__o21ai_1
XFILLER_188_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18542__A1 _17434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14159__A2 _14857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19258_ _19117_/A _19117_/B _19117_/C _19116_/B vssd1 vssd1 vccd1 vccd1 _19258_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_137_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19619__D _19619_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18209_ _18216_/B _18216_/A vssd1 vssd1 vccd1 vccd1 _18212_/A sky130_fd_sc_hd__xor2_1
XFILLER_117_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19189_ _19190_/A _19190_/B _19190_/C vssd1 vssd1 vccd1 vccd1 _19343_/B sky130_fd_sc_hd__a21o_1
XFILLER_191_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21220_ _21220_/A vssd1 vssd1 vccd1 vccd1 _21220_/X sky130_fd_sc_hd__buf_2
XANTENNA__16324__C _16324_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16305__B1 _15711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__A2 _11381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21151_ _21142_/A _21151_/B vssd1 vssd1 vccd1 vccd1 _21151_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11468__C _11942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20102_ _20110_/A _20110_/B _20250_/C _20096_/Y _16261_/B vssd1 vssd1 vccd1 vccd1
+ _20119_/D sky130_fd_sc_hd__o2111ai_4
XFILLER_144_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21082_ _21082_/A _21082_/B _21082_/C _21081_/C vssd1 vssd1 vccd1 vccd1 _21086_/A
+ sky130_fd_sc_hd__or4b_2
XANTENNA__17436__B _21011_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20143__A _20143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20033_ _20033_/A vssd1 vssd1 vccd1 vccd1 _20034_/B sky130_fd_sc_hd__inv_2
XANTENNA__21601__A1 _13633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19651__B _19651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12299__C _20694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21984_ _22029_/A _21994_/A vssd1 vssd1 vccd1 vccd1 _21993_/A sky130_fd_sc_hd__nand2_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ _20924_/X _20926_/X _20937_/A vssd1 vssd1 vccd1 vccd1 _20935_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_183_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16387__A3 _15339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20866_ _20866_/A _20866_/B vssd1 vssd1 vccd1 vccd1 _20866_/X sky130_fd_sc_hd__and2_1
XFILLER_168_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22605_ _22605_/A vssd1 vssd1 vccd1 vccd1 _22791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20797_ _20797_/A _20797_/B _20797_/C _20797_/D vssd1 vssd1 vccd1 vccd1 _20869_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_50_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15700__A _15707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22536_ _22761_/Q input66/X _22536_/S vssd1 vssd1 vccd1 vccd1 _22537_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20340__A1 _12450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16515__B _18192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22617__A0 _18698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22467_ _21329_/B input36/X _22475_/S vssd1 vssd1 vccd1 vccd1 _22468_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14929__D_N _14845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ _12220_/A _12220_/B vssd1 vssd1 vccd1 vccd1 _18223_/A sky130_fd_sc_hd__nand2_2
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21418_ _21553_/A _21417_/B _21299_/X _21251_/X vssd1 vssd1 vccd1 vccd1 _21440_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_136_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22398_ _22700_/Q input38/X _22402_/S vssd1 vssd1 vccd1 vccd1 _22399_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12581__A1 _20486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12151_ _18339_/A vssd1 vssd1 vccd1 vccd1 _19016_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12581__B2 _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21349_ _13101_/A _13101_/B _13350_/A vssd1 vssd1 vccd1 vccd1 _21349_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16311__A3 _15792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12082_ _12029_/Y _12039_/Y _12081_/Y vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__a21o_1
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15910_ _15978_/A _15978_/B _15792_/B _15933_/A vssd1 vssd1 vccd1 vccd1 _16011_/A
+ sky130_fd_sc_hd__o2bb2ai_4
XANTENNA__19842__A _19842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16890_ _16444_/Y _16445_/X _16644_/Y _16645_/X vssd1 vssd1 vccd1 vccd1 _16890_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15807__C1 _16106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16075__A2 _20728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _15748_/A _15748_/B _12765_/X _15840_/X vssd1 vssd1 vccd1 vccd1 _15842_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14086__B2 _14270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17362__A _17373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _18519_/Y _18523_/Y _18527_/Y _18548_/A _18548_/B vssd1 vssd1 vccd1 vccd1
+ _18561_/C sky130_fd_sc_hd__o2111ai_1
XANTENNA__12097__B1 _15557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _15350_/Y _15646_/X _15389_/C _15389_/A vssd1 vssd1 vccd1 vccd1 _16209_/C
+ sky130_fd_sc_hd__a22o_1
X_12984_ _15799_/A vssd1 vssd1 vccd1 vccd1 _20452_/A sky130_fd_sc_hd__buf_2
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _17719_/B _17511_/B vssd1 vssd1 vccd1 vccd1 _22958_/D sky130_fd_sc_hd__xor2_1
XANTENNA__17024__B2 _16742_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11935_ _18292_/A _11935_/B _11935_/C vssd1 vssd1 vccd1 vccd1 _11935_/X sky130_fd_sc_hd__or3_4
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14723_ _13950_/X _14619_/A _14722_/Y vssd1 vssd1 vccd1 vccd1 _14727_/C sky130_fd_sc_hd__o21ai_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ _18491_/A vssd1 vssd1 vccd1 vccd1 _18915_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_884 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17442_ _17442_/A vssd1 vssd1 vccd1 vccd1 _17442_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _14536_/Y _14524_/Y _14541_/D vssd1 vssd1 vccd1 vccd1 _14655_/B sky130_fd_sc_hd__o21a_1
XFILLER_178_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _18985_/C vssd1 vssd1 vccd1 vccd1 _19154_/C sky130_fd_sc_hd__buf_2
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13605_ _13627_/C _13589_/X _13627_/B _13603_/Y _13604_/X vssd1 vssd1 vccd1 vccd1
+ _13605_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_177_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17373_ _17373_/A vssd1 vssd1 vccd1 vccd1 _18044_/A sky130_fd_sc_hd__clkbuf_2
X_14585_ _14571_/A _14583_/Y _14863_/A vssd1 vssd1 vccd1 vccd1 _14786_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__14794__C1 _13873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_720 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18193__A _18193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11797_ _11797_/A _11797_/B vssd1 vssd1 vccd1 vccd1 _11799_/B sky130_fd_sc_hd__nand2_1
X_19112_ _19112_/A _19112_/B _19303_/A _19116_/A vssd1 vssd1 vccd1 vccd1 _19122_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_14_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13536_ _13533_/Y _13534_/Y _13455_/Y vssd1 vssd1 vccd1 vccd1 _13537_/A sky130_fd_sc_hd__o21ai_1
X_16324_ _22701_/Q _16324_/B _16324_/C vssd1 vssd1 vccd1 vccd1 _16325_/B sky130_fd_sc_hd__nand3b_2
XFILLER_159_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22608__A0 _12107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19043_ _19043_/A vssd1 vssd1 vccd1 vccd1 _19043_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16255_ _16540_/A _16288_/C vssd1 vssd1 vccd1 vccd1 _16282_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15889__A2 _16155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13467_ _13455_/Y _13537_/B _13470_/A vssd1 vssd1 vccd1 vccd1 _13468_/C sky130_fd_sc_hd__a21boi_1
XFILLER_127_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15206_ _15206_/A _15206_/B vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__or2_1
XFILLER_145_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12418_ _12418_/A vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__buf_4
XFILLER_161_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16186_ _16186_/A _16186_/B vssd1 vssd1 vccd1 vccd1 _16186_/Y sky130_fd_sc_hd__nor2_1
X_13398_ _13339_/Y _13353_/Y _13359_/X _13391_/B vssd1 vssd1 vccd1 vccd1 _13399_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_127_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16838__A1 _16451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ _15092_/A _15095_/B _15135_/B vssd1 vssd1 vccd1 vccd1 _15173_/A sky130_fd_sc_hd__a21oi_1
X_12349_ _22819_/Q vssd1 vssd1 vccd1 vccd1 _20338_/C sky130_fd_sc_hd__buf_2
XANTENNA__19455__C _19455_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14849__B1 _14552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19945_ _19945_/A _19945_/B _19945_/C _19945_/D vssd1 vssd1 vccd1 vccd1 _19946_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15068_ _15114_/C vssd1 vssd1 vccd1 vccd1 _15154_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16160__B _16997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14019_ _13867_/A _14169_/C _13838_/X vssd1 vssd1 vccd1 vccd1 _14022_/A sky130_fd_sc_hd__a21oi_1
XFILLER_96_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19876_ _19834_/Y _19835_/Y _19881_/C vssd1 vssd1 vccd1 vccd1 _19878_/A sky130_fd_sc_hd__o21ai_1
XFILLER_122_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18460__B1 _17817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18827_ _18827_/A _18827_/B vssd1 vssd1 vccd1 vccd1 _18827_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15274__B1 _15271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15813__A2 _12493_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18758_ _18748_/B _18748_/A _18608_/Y _18609_/Y vssd1 vssd1 vccd1 vccd1 _18758_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12627__A2 _20502_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13824__A1 _13820_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17015__A1 _17006_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17709_ _17226_/A _17227_/A _17623_/Y _17705_/Y _17708_/Y vssd1 vssd1 vccd1 vccd1
+ _17709_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_36_564 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18689_ _11394_/A _18116_/D _18677_/B _18128_/A vssd1 vssd1 vccd1 vccd1 _18890_/A
+ sky130_fd_sc_hd__o211a_2
XANTENNA__17566__A2 _17728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13305__A _13305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16319__C _16319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20720_ _20720_/A _20720_/B _20720_/C vssd1 vssd1 vccd1 vccd1 _20721_/C sky130_fd_sc_hd__nand3_1
XANTENNA__16774__B1 _15538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19199__A _19199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20651_ _20538_/B _20538_/C _20653_/A vssd1 vssd1 vccd1 vccd1 _20652_/C sky130_fd_sc_hd__a21boi_1
XFILLER_189_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18515__B2 _18510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22872__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20322__A1 _12680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20582_ _20582_/A _20792_/C _20582_/C vssd1 vssd1 vccd1 vccd1 _20697_/B sky130_fd_sc_hd__nand3_2
XFILLER_192_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22321_ _22300_/B _22300_/A _22284_/C _22341_/C vssd1 vssd1 vccd1 vccd1 _22323_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_178_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16054__C _16498_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22252_ _22208_/B _22211_/B _22208_/A vssd1 vssd1 vccd1 vccd1 _22253_/B sky130_fd_sc_hd__a21boi_1
XFILLER_191_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21203_ _13305_/A _13305_/B _13577_/A vssd1 vssd1 vccd1 vccd1 _21203_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17447__A _19012_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13975__A _14112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22183_ _22186_/A _22186_/B vssd1 vssd1 vccd1 vccd1 _22183_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__19491__A2 _17632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21134_ _21086_/C _21086_/D _21086_/B _21112_/B _21112_/A vssd1 vssd1 vccd1 vccd1
+ _21135_/B sky130_fd_sc_hd__a32oi_4
XFILLER_120_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20592__A1_N _20593_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20389__A1 _20378_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21065_ _21068_/A _21068_/B _21037_/D _21079_/A vssd1 vssd1 vccd1 vccd1 _21065_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21586__B1 _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17254__A1 _16040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16057__A2 _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20016_ _20016_/A _20016_/B vssd1 vssd1 vccd1 vccd1 _20018_/A sky130_fd_sc_hd__xnor2_1
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18278__A _18278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16462__C1 _15694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11942__B _18107_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21967_ _21767_/X _21970_/A _21740_/X _22045_/A vssd1 vssd1 vccd1 vccd1 _21967_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11720_/A vssd1 vssd1 vccd1 vccd1 _11721_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__21353__A3 _21220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20918_ _21009_/A _17733_/A _17460_/A _20917_/Y _20910_/Y vssd1 vssd1 vccd1 vccd1
+ _20920_/B sky130_fd_sc_hd__o221ai_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21898_ _21902_/B _21901_/A vssd1 vssd1 vccd1 vccd1 _21899_/D sky130_fd_sc_hd__nand2_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21432__A _22674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11651_ _11942_/A vssd1 vssd1 vccd1 vccd1 _18459_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20849_ _13022_/B _17728_/A _20697_/B _20848_/Y vssd1 vssd1 vccd1 vccd1 _20849_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14370_ _14370_/A vssd1 vssd1 vccd1 vccd1 _14370_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11582_ _18690_/B vssd1 vssd1 vccd1 vccd1 _16313_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13321_ _21606_/A _13319_/X _13126_/X _21318_/A vssd1 vssd1 vccd1 vccd1 _13321_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_168_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22519_ _13776_/A input46/X _22525_/S vssd1 vssd1 vccd1 vccd1 _22520_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15725__D1 _20870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ _16040_/A vssd1 vssd1 vccd1 vccd1 _20728_/B sky130_fd_sc_hd__buf_4
XFILLER_108_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13252_ _13504_/B _13504_/C vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__nor2_1
XANTENNA__15367__A2_N _15382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input74_A x[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12203_ _19587_/C vssd1 vssd1 vccd1 vccd1 _19772_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__12554__A1 _12771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21813__A1 _21805_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20616__A2 _15723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_439 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13183_ _13143_/A _13143_/B _13158_/A _21473_/A vssd1 vssd1 vccd1 vccd1 _13185_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__16261__A _19322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12134_ _12134_/A _12134_/B vssd1 vssd1 vccd1 vccd1 _12138_/A sky130_fd_sc_hd__nand2_1
XFILLER_150_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17991_ _17991_/A _17991_/B _17991_/C vssd1 vssd1 vccd1 vccd1 _18061_/A sky130_fd_sc_hd__and3_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17507__D _17959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19730_ _19725_/B _19725_/C _19725_/A vssd1 vssd1 vccd1 vccd1 _19731_/B sky130_fd_sc_hd__a21oi_1
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16942_ _18192_/A vssd1 vssd1 vccd1 vccd1 _19199_/B sky130_fd_sc_hd__buf_2
X_12065_ _12065_/A vssd1 vssd1 vccd1 vccd1 _16192_/D sky130_fd_sc_hd__buf_2
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15175__A_N _15101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14212__C _15004_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19661_ _19132_/A _19132_/B _19132_/C _18973_/Y vssd1 vssd1 vccd1 vccd1 _19664_/A
+ sky130_fd_sc_hd__a31o_1
X_16873_ _16873_/A _16873_/B _16873_/C _16873_/D vssd1 vssd1 vccd1 vccd1 _16874_/C
+ sky130_fd_sc_hd__nand4_1
X_18612_ _12170_/X _12171_/X _19197_/C _19197_/D vssd1 vssd1 vccd1 vccd1 _18613_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__16453__C1 _16452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ _15824_/A _15824_/B _15824_/C vssd1 vssd1 vccd1 vccd1 _15849_/A sky130_fd_sc_hd__and3_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ _19359_/X _19500_/X _19497_/B _19494_/Y vssd1 vssd1 vccd1 vccd1 _19594_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_93_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17523__C _17523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _18543_/A _18543_/B _18543_/C vssd1 vssd1 vccd1 vccd1 _18553_/B sky130_fd_sc_hd__nand3_2
XANTENNA__11817__B1 _11685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15755_ _15755_/A _15755_/B vssd1 vssd1 vccd1 vccd1 _15842_/A sky130_fd_sc_hd__nor2_2
X_12967_ _12967_/A vssd1 vssd1 vccd1 vccd1 _20697_/A sky130_fd_sc_hd__buf_2
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17548__A2 _17388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_512 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22895__CLK _22952_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _11918_/A _11918_/B vssd1 vssd1 vccd1 vccd1 _11918_/Y sky130_fd_sc_hd__nand2_1
X_14706_ _14779_/A _14706_/B _14861_/A _15115_/B vssd1 vssd1 vccd1 vccd1 _14708_/D
+ sky130_fd_sc_hd__nand4_2
X_18474_ _18474_/A _18474_/B vssd1 vssd1 vccd1 vccd1 _18474_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20552__A1 _20195_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15686_ _15766_/A _15859_/D _15738_/A vssd1 vssd1 vccd1 vccd1 _15686_/Y sky130_fd_sc_hd__a21boi_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12898_ _12898_/A _12898_/B _12898_/C vssd1 vssd1 vccd1 vccd1 _12900_/B sky130_fd_sc_hd__nand3_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17425_ _17421_/X _17422_/X _17423_/X _17424_/X vssd1 vssd1 vccd1 vccd1 _17426_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1097 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11849_ _19329_/C vssd1 vssd1 vccd1 vccd1 _17313_/D sky130_fd_sc_hd__clkbuf_4
X_14637_ _14498_/Y _14518_/Y _14522_/B vssd1 vssd1 vccd1 vccd1 _14650_/C sky130_fd_sc_hd__o21ai_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16436__A _18258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15978__C _15978_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15340__A _15797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17356_ _17226_/X _17227_/X _17228_/Y _17215_/Y _17372_/C vssd1 vssd1 vccd1 vccd1
+ _17616_/C sky130_fd_sc_hd__o221a_1
X_14568_ _14568_/A _14568_/B vssd1 vssd1 vccd1 vccd1 _14568_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19170__A1 _17421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16307_ _20605_/B vssd1 vssd1 vccd1 vccd1 _20608_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15716__D1 _17128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13519_ _13521_/A _13519_/B _13521_/C vssd1 vssd1 vccd1 vccd1 _13520_/B sky130_fd_sc_hd__nand3_2
XANTENNA__20855__A2 _17435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17287_ _17293_/A _17282_/A _17286_/X vssd1 vssd1 vccd1 vccd1 _17290_/A sky130_fd_sc_hd__a21o_1
X_14499_ _14611_/A vssd1 vssd1 vccd1 vccd1 _14499_/Y sky130_fd_sc_hd__inv_2
X_19026_ _19026_/A _19026_/B vssd1 vssd1 vccd1 vccd1 _19026_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16238_ _16532_/B _16238_/B _16532_/A vssd1 vssd1 vccd1 vccd1 _16504_/A sky130_fd_sc_hd__nand3_1
XFILLER_174_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13795__A _22868_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16169_ _16169_/A _16169_/B _16169_/C _16169_/D vssd1 vssd1 vccd1 vccd1 _16169_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_138_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16602__C _16602_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19928_ _19928_/A _19928_/B vssd1 vssd1 vccd1 vccd1 _19970_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19482__A _19482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12204__A _18203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17236__A1 _15723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18433__B1 _18432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19859_ _19859_/A vssd1 vssd1 vccd1 vccd1 _19859_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15798__A1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22870_ _22916_/CLK _22870_/D vssd1 vssd1 vccd1 vccd1 _22870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20791__A1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11762__B _11762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21821_ _21821_/A _21834_/C _21834_/D _22089_/A vssd1 vssd1 vccd1 vccd1 _21825_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_71_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17730__A _17730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21752_ _21874_/C _21748_/Y _21758_/D vssd1 vssd1 vccd1 vccd1 _21753_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__16747__B1 _16732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20703_ _12968_/A _16746_/X _20464_/B _20579_/X _20695_/A vssd1 vssd1 vccd1 vccd1
+ _20703_/X sky130_fd_sc_hd__o311a_1
XFILLER_93_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21683_ _21683_/A vssd1 vssd1 vccd1 vccd1 _22229_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20634_ _20630_/A _20634_/B _20634_/C vssd1 vssd1 vccd1 vccd1 _20738_/C sky130_fd_sc_hd__nand3b_1
XANTENNA__14773__A2 _13973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13576__A3 _13162_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20846__A2 _16585_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20565_ _22933_/Q vssd1 vssd1 vccd1 vccd1 _20565_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22304_ _22304_/A _22304_/B _22304_/C _22308_/A vssd1 vssd1 vccd1 vccd1 _22306_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_153_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15722__A1 _15649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20496_ _20347_/B _20343_/Y _20339_/Y vssd1 vssd1 vccd1 vccd1 _20496_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_180_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22235_ _22238_/B _22193_/B _22178_/B _22219_/Y _22237_/A vssd1 vssd1 vccd1 vccd1
+ _22240_/B sky130_fd_sc_hd__a311o_1
XFILLER_3_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22166_ _22084_/A _22160_/Y _22165_/X vssd1 vssd1 vccd1 vccd1 _22166_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_121_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21117_ _21135_/A _21118_/C _21118_/A vssd1 vssd1 vccd1 vccd1 _21119_/A sky130_fd_sc_hd__a21oi_1
XFILLER_132_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22097_ _21841_/A _21958_/X _22099_/A _22047_/Y _22099_/B vssd1 vssd1 vccd1 vccd1
+ _22102_/A sky130_fd_sc_hd__o221ai_2
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21048_ _21082_/B _21048_/B _21048_/C _21046_/B vssd1 vssd1 vccd1 vccd1 _21090_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11953__A _16447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15789__A1 _12413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13870_ _13799_/X _13820_/A _13826_/B _22759_/Q vssd1 vssd1 vccd1 vccd1 _14722_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13871__C _14722_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ _22696_/Q _22697_/Q vssd1 vssd1 vccd1 vccd1 _16323_/C sky130_fd_sc_hd__nor2_2
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15540_ _12046_/X _15495_/X _18258_/B _16241_/D vssd1 vssd1 vccd1 vccd1 _15548_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _12665_/A _12665_/B _12898_/A _12898_/B vssd1 vssd1 vccd1 vccd1 _12895_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__16738__B1 _16098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11703_ _11381_/X _12111_/A _11702_/X _11512_/A vssd1 vssd1 vccd1 vccd1 _11703_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15471_ _19587_/C _15586_/C _15528_/A _15901_/C vssd1 vssd1 vccd1 vccd1 _15474_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12683_/A vssd1 vssd1 vccd1 vccd1 _20593_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_188_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16256__A _16256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14213__A1 _14765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15410__B1 _15637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17603_/C _17210_/B vssd1 vssd1 vccd1 vccd1 _17213_/C sky130_fd_sc_hd__nor2_1
X_14422_ _22716_/Q _14418_/X _14410_/X _22748_/Q _14421_/X vssd1 vssd1 vccd1 vccd1
+ _14422_/X sky130_fd_sc_hd__a221o_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11634_/A vssd1 vssd1 vccd1 vccd1 _19043_/A sky130_fd_sc_hd__buf_2
XFILLER_30_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18190_ _18183_/Y _18187_/Y _18188_/Y _18189_/Y vssd1 vssd1 vccd1 vccd1 _18191_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_168_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12775__A1 _12772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17141_ _17141_/A _17532_/C _17532_/D vssd1 vssd1 vccd1 vccd1 _17142_/A sky130_fd_sc_hd__nand3_1
X_14353_ _22794_/Q vssd1 vssd1 vccd1 vccd1 _18127_/B sky130_fd_sc_hd__buf_2
XANTENNA__12934__D _20355_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11565_ _11565_/A _11565_/B vssd1 vssd1 vccd1 vccd1 _11565_/Y sky130_fd_sc_hd__nand2_2
XFILLER_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18360__C1 _11351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13304_ _13304_/A _13304_/B vssd1 vssd1 vccd1 vccd1 _13305_/B sky130_fd_sc_hd__nand2_2
X_17072_ _17071_/A _17071_/B _17071_/C vssd1 vssd1 vccd1 vccd1 _17073_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__22039__A1 _21853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14284_ _14282_/A _14282_/B _14254_/X _14283_/Y vssd1 vssd1 vccd1 vccd1 _14289_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_156_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11496_ _22790_/Q _11496_/B vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16023_ _15945_/A _15945_/B _15945_/C vssd1 vssd1 vccd1 vccd1 _16024_/B sky130_fd_sc_hd__a21oi_1
X_13235_ _13504_/C vssd1 vssd1 vccd1 vccd1 _13633_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13166_ _13286_/C _13286_/D vssd1 vssd1 vccd1 vccd1 _13166_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15319__B _15319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12117_ _12117_/A vssd1 vssd1 vccd1 vccd1 _12118_/A sky130_fd_sc_hd__buf_4
XFILLER_123_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17974_ _17974_/A vssd1 vssd1 vccd1 vccd1 _17989_/A sky130_fd_sc_hd__inv_2
XFILLER_112_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13097_ _13097_/A vssd1 vssd1 vccd1 vccd1 _13098_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19713_ _19707_/Y _19864_/A _19712_/X vssd1 vssd1 vccd1 vccd1 _19799_/B sky130_fd_sc_hd__a21o_1
XFILLER_111_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16925_ _18666_/B _17386_/B _20675_/B vssd1 vssd1 vccd1 vccd1 _16926_/B sky130_fd_sc_hd__and3_1
X_12048_ _16477_/A vssd1 vssd1 vccd1 vccd1 _19197_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_38_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_90 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20241__A _20241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19644_ _19641_/X _19643_/Y _19649_/B vssd1 vssd1 vccd1 vccd1 _19644_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15335__A _15335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16856_ _16860_/B _16860_/C _16860_/A vssd1 vssd1 vccd1 vccd1 _16856_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13781__C _14199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15807_ _15302_/A _15691_/Y _15805_/Y _16106_/A _17436_/A vssd1 vssd1 vccd1 vccd1
+ _15824_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19575_ _19575_/A _19575_/B vssd1 vssd1 vccd1 vccd1 _22898_/D sky130_fd_sc_hd__nor2_1
XFILLER_19_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16787_ _16178_/A _17634_/A _16941_/A vssd1 vssd1 vccd1 vccd1 _16787_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13999_ _14007_/B _14009_/B _14497_/A vssd1 vssd1 vccd1 vccd1 _14006_/A sky130_fd_sc_hd__nand3_1
X_18526_ _18526_/A _18526_/B _18915_/A _18526_/D vssd1 vssd1 vccd1 vccd1 _18527_/C
+ sky130_fd_sc_hd__nand4_2
X_15738_ _15738_/A _15738_/B vssd1 vssd1 vccd1 vccd1 _15860_/B sky130_fd_sc_hd__nand2_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18194__A2 _11503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18457_ _18458_/C _18458_/A _18458_/B vssd1 vssd1 vccd1 vccd1 _18457_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__12694__A _17246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15669_ _16213_/A vssd1 vssd1 vccd1 vccd1 _15673_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17408_ _17408_/A _17408_/B vssd1 vssd1 vccd1 vccd1 _17408_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12215__B1 _18445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18388_ _18388_/A vssd1 vssd1 vccd1 vccd1 _18407_/B sky130_fd_sc_hd__buf_2
XFILLER_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17339_ _17341_/A _17341_/B _17341_/C _17341_/D _17338_/X vssd1 vssd1 vccd1 vccd1
+ _17339_/X sky130_fd_sc_hd__a41o_1
XFILLER_119_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14117__C _14786_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_0_0_bq_clk_i clkbuf_2_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14507__A2 _13924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20350_ _12734_/X _16611_/A _20347_/A vssd1 vssd1 vccd1 vccd1 _20353_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__16362__D1 _16400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20416__A _20449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16613__B _17431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19009_ _19009_/A _19009_/B _19009_/C _19009_/D vssd1 vssd1 vccd1 vccd1 _19237_/A
+ sky130_fd_sc_hd__nand4_4
XANTENNA__22910__CLK _22922_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20281_ _20281_/A _20281_/B _20284_/C vssd1 vssd1 vccd1 vccd1 _20281_/X sky130_fd_sc_hd__and3_1
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22020_ _21922_/Y _21927_/X _21925_/Y vssd1 vssd1 vccd1 vccd1 _22021_/B sky130_fd_sc_hd__a21boi_1
XFILLER_161_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11757__B _12165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11741__A2 _17427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16051__D _16103_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22922_ _22922_/CLK _22922_/D vssd1 vssd1 vccd1 vccd1 _22922_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16968__B1 _15840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22853_ _22937_/CLK _22865_/Q vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17460__A _17460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21804_ _21804_/A vssd1 vssd1 vccd1 vccd1 _21913_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22784_ _22797_/CLK _22784_/D vssd1 vssd1 vccd1 vccd1 _22784_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21735_ _21737_/B _21737_/A vssd1 vssd1 vccd1 vccd1 _21790_/A sky130_fd_sc_hd__nand2_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21666_ _21666_/A _21666_/B vssd1 vssd1 vccd1 vccd1 _21666_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20617_ _20479_/Y _20614_/Y _20615_/Y _20616_/X vssd1 vssd1 vccd1 vccd1 _20620_/C
+ sky130_fd_sc_hd__o22ai_4
XFILLER_138_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21597_ _13662_/A _21594_/Y _21482_/B _21751_/A _21758_/A vssd1 vssd1 vccd1 vccd1
+ _21771_/C sky130_fd_sc_hd__o221ai_2
XFILLER_177_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16499__A2 _15435_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ _11429_/A _18099_/A _11349_/X vssd1 vssd1 vccd1 vccd1 _12090_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__18893__B1 _19771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20548_ _20754_/A _20754_/B _20445_/Y _20547_/X vssd1 vssd1 vccd1 vccd1 _20548_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11948__A _15633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ _22799_/Q vssd1 vssd1 vccd1 vccd1 _11421_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_20479_ _20482_/A _20482_/B vssd1 vssd1 vccd1 vccd1 _20479_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__17448__A1 _17426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ _16106_/A vssd1 vssd1 vccd1 vccd1 _20284_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22218_ _22195_/B _22195_/A _22217_/Y vssd1 vssd1 vccd1 vccd1 _22243_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__17448__B2 _20917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17635__A _17635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22149_ _22150_/A _22150_/B _22681_/Q vssd1 vssd1 vccd1 vccd1 _22290_/C sky130_fd_sc_hd__a21o_1
XFILLER_160_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input37_A wb_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14971_ _14971_/A _14971_/B _14971_/C vssd1 vssd1 vccd1 vccd1 _14971_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__14682__A1 _14998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12142__C1 _18510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18948__B2 _18625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11683__A _11702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16710_ _11511_/A _16708_/X _16709_/Y vssd1 vssd1 vccd1 vccd1 _16710_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__14682__B2 _14942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13922_ _13838_/X _13868_/X _13917_/Y _13921_/X vssd1 vssd1 vccd1 vccd1 _14052_/A
+ sky130_fd_sc_hd__o211ai_4
X_17690_ _17690_/A vssd1 vssd1 vccd1 vccd1 _17697_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16641_ _20972_/B vssd1 vssd1 vccd1 vccd1 _17806_/D sky130_fd_sc_hd__buf_2
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13853_ _13984_/A _13968_/C _14777_/C _14126_/A vssd1 vssd1 vccd1 vccd1 _13854_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_75_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19360_ _12202_/A _12202_/B _19176_/A vssd1 vssd1 vccd1 vccd1 _19360_/Y sky130_fd_sc_hd__a21oi_1
X_12804_ _12577_/A _12576_/A _12802_/C _12348_/A _12578_/A vssd1 vssd1 vccd1 vccd1
+ _12804_/Y sky130_fd_sc_hd__o2111ai_4
X_16572_ _16435_/B _16579_/A _16580_/A _16571_/Y vssd1 vssd1 vccd1 vccd1 _20579_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_43_640 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13784_ _13784_/A _14043_/B vssd1 vssd1 vccd1 vccd1 _13786_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18185__B _18278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18311_ _18389_/A _18389_/B _18389_/C _18310_/Y _18383_/A vssd1 vssd1 vccd1 vccd1
+ _18311_/X sky130_fd_sc_hd__a32o_1
X_15523_ _15523_/A vssd1 vssd1 vccd1 vccd1 _15523_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19291_ _19290_/A _19290_/B _19290_/C vssd1 vssd1 vccd1 vccd1 _19292_/B sky130_fd_sc_hd__a21oi_1
X_12735_ _15450_/A vssd1 vssd1 vccd1 vccd1 _12735_/X sky130_fd_sc_hd__buf_4
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17520__D _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12460__A3 _20694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _12250_/D _18236_/Y _18240_/Y _18772_/A vssd1 vssd1 vccd1 vccd1 _18251_/B
+ sky130_fd_sc_hd__a2bb2oi_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15454_ _15454_/A vssd1 vssd1 vccd1 vccd1 _15457_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12666_/A _12898_/C vssd1 vssd1 vccd1 vccd1 _12895_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11617_ _11974_/A vssd1 vssd1 vccd1 vccd1 _18328_/C sky130_fd_sc_hd__buf_2
X_14405_ _22710_/Q _14403_/X _14396_/X _22742_/Q _14404_/X vssd1 vssd1 vccd1 vccd1
+ _14405_/X sky130_fd_sc_hd__a221o_1
X_18173_ _18173_/A _18173_/B _18173_/C vssd1 vssd1 vccd1 vccd1 _18174_/A sky130_fd_sc_hd__nand3_1
X_15385_ _15385_/A vssd1 vssd1 vccd1 vccd1 _15682_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12597_ _12445_/Y _12595_/Y _12697_/A _15569_/A vssd1 vssd1 vccd1 vccd1 _12601_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_11_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17124_ _17323_/A _17122_/Y _17123_/X vssd1 vssd1 vccd1 vccd1 _17178_/A sky130_fd_sc_hd__a21o_1
X_14336_ _12387_/B _14308_/X _14313_/X _13161_/C _14335_/X vssd1 vssd1 vccd1 vccd1
+ _14336_/X sky130_fd_sc_hd__a221o_1
X_11548_ _11552_/A _11537_/A _11553_/B vssd1 vssd1 vccd1 vccd1 _11548_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11971__A2 _15905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17055_ _17603_/A _17603_/B _17048_/Y _16659_/B _17054_/Y vssd1 vssd1 vccd1 vccd1
+ _17060_/A sky130_fd_sc_hd__o221ai_4
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14267_ _14267_/A _14267_/B _14267_/C vssd1 vssd1 vccd1 vccd1 _14269_/D sky130_fd_sc_hd__nand3_1
XFILLER_143_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11479_ _15633_/A vssd1 vssd1 vccd1 vccd1 _12094_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16006_ _16006_/A _16006_/B vssd1 vssd1 vccd1 vccd1 _16045_/C sky130_fd_sc_hd__nand2_1
X_13218_ _21591_/B vssd1 vssd1 vccd1 vccd1 _21757_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_125_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18097__D1 _18810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14198_ _14198_/A _14198_/B _14198_/C _14198_/D vssd1 vssd1 vccd1 vccd1 _14255_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13149_ _22845_/Q vssd1 vssd1 vccd1 vccd1 _13502_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15991__C _16129_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13792__B _15082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17957_ _17957_/A _17957_/B vssd1 vssd1 vccd1 vccd1 _17958_/B sky130_fd_sc_hd__nor2_1
XFILLER_111_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12689__A _12689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16908_ _16908_/A _16908_/B _16908_/C vssd1 vssd1 vccd1 vccd1 _16908_/X sky130_fd_sc_hd__and3_1
XFILLER_66_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17888_ _17888_/A _17888_/B vssd1 vssd1 vccd1 vccd1 _17889_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19627_ _19621_/Y _19622_/X _19626_/X vssd1 vssd1 vccd1 vccd1 _19629_/B sky130_fd_sc_hd__a21boi_2
X_16839_ _16845_/C _16845_/D vssd1 vssd1 vccd1 vccd1 _17189_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12201__B _22662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15622__B1 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17280__A _17280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19558_ _19454_/X _19455_/X _19545_/Y _19549_/Y vssd1 vssd1 vccd1 vccd1 _19558_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13016__C _13016_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19364__A1 _11639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18509_ _18876_/A vssd1 vssd1 vccd1 vccd1 _19614_/B sky130_fd_sc_hd__buf_2
XANTENNA__12987__A1 _20452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19489_ _11639_/X _17526_/X _19215_/X _19352_/X vssd1 vssd1 vccd1 vccd1 _19489_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__21171__A1 _13434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21520_ _21369_/A _21369_/B _21369_/C _21369_/D vssd1 vssd1 vccd1 vccd1 _21520_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_167_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21451_ _21853_/A _13343_/X _21450_/Y vssd1 vssd1 vccd1 vccd1 _21460_/B sky130_fd_sc_hd__o21ai_1
XFILLER_119_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19785__A_N _19788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20402_ _20400_/Y _20272_/Y _20269_/X _20401_/Y vssd1 vssd1 vccd1 vccd1 _20427_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19000__A _19000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21382_ _21460_/A _21344_/D _21349_/X vssd1 vssd1 vccd1 vccd1 _21385_/A sky130_fd_sc_hd__a21o_1
XANTENNA__15689__B1 _12719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11962__A2 _11703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20333_ _20242_/X _20244_/X _20262_/C vssd1 vssd1 vccd1 vccd1 _20335_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__12590__C _20461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18627__B1 _18636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20264_ _20264_/A _20390_/D vssd1 vssd1 vccd1 vccd1 _20264_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22003_ _21897_/B _21842_/X _21733_/A _21841_/Y vssd1 vssd1 vccd1 vccd1 _22003_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12911__A1 _15988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16997__C _16997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13983__A _22867_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12911__B2 _20593_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16102__A1 _16103_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20195_ _13045_/A _13045_/B _20194_/Y vssd1 vssd1 vccd1 vccd1 _20195_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_163_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15310__C1 _15694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12599__A _20323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22905_ _22949_/CLK _22905_/D vssd1 vssd1 vccd1 vccd1 _22905_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22836_ _22850_/CLK _22848_/Q vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12427__B1 _12343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19355__A1 _16940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12978__A1 _12522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22956__CLK _22959_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22767_ _22805_/CLK _22767_/D vssd1 vssd1 vccd1 vccd1 _22767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_824 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ _12520_/A _12520_/B vssd1 vssd1 vccd1 vccd1 _12550_/C sky130_fd_sc_hd__nand2_2
XFILLER_72_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21718_ _21654_/A _21654_/C _21717_/Y vssd1 vssd1 vccd1 vccd1 _21719_/B sky130_fd_sc_hd__a21oi_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11650__A1 _11507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14719__A2 _13851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22698_ _22701_/CLK _22698_/D vssd1 vssd1 vccd1 vccd1 _22698_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ _12448_/Y _12449_/Y _12450_/X _12420_/X vssd1 vssd1 vccd1 vccd1 _12454_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_138_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21649_ _21649_/A _21649_/B vssd1 vssd1 vccd1 vccd1 _21650_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11402_ _11502_/A _11503_/A vssd1 vssd1 vccd1 vccd1 _11512_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17669__A1 _16124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15170_ _15169_/B _15181_/B _15169_/A vssd1 vssd1 vccd1 vccd1 _15171_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__18866__B1 _11639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ _22821_/Q vssd1 vssd1 vccd1 vccd1 _20207_/C sky130_fd_sc_hd__buf_2
XFILLER_181_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14121_ _14117_/Y _14118_/Y _14120_/Y vssd1 vssd1 vccd1 vccd1 _14237_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__11678__A _11819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20673__B1 _20853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11333_ _11333_/A vssd1 vssd1 vccd1 vccd1 _11333_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ _14052_/A _14052_/B _14052_/C vssd1 vssd1 vccd1 vccd1 _14094_/B sky130_fd_sc_hd__nand3_2
XFILLER_153_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16629__C1 _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13003_ _13003_/A _13003_/B _13003_/C vssd1 vssd1 vccd1 vccd1 _13004_/C sky130_fd_sc_hd__nand3_1
X_18860_ _15887_/X _19695_/A _19313_/A _11845_/X vssd1 vssd1 vccd1 vccd1 _19091_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_121_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20976__A1 _20917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17811_ _19844_/B _20936_/C _17895_/A _17811_/D vssd1 vssd1 vccd1 vccd1 _17895_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_122_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ _18970_/A _18970_/C vssd1 vssd1 vccd1 vccd1 _18792_/B sky130_fd_sc_hd__and2_1
XANTENNA__13458__A2 _21621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17742_ _17649_/X _17648_/Y _17652_/Y _17535_/B vssd1 vssd1 vccd1 vccd1 _17744_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14954_ _15064_/C _15070_/A _14857_/B _14952_/A _15002_/B vssd1 vssd1 vccd1 vccd1
+ _14954_/X sky130_fd_sc_hd__a32o_1
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14220__C _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ _14506_/C _13959_/A vssd1 vssd1 vccd1 vccd1 _13905_/Y sky130_fd_sc_hd__nand2_2
XFILLER_78_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17673_ _19334_/B vssd1 vssd1 vccd1 vccd1 _19793_/C sky130_fd_sc_hd__buf_2
X_14885_ _14885_/A _14885_/B vssd1 vssd1 vccd1 vccd1 _14885_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_584 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19412_ _19404_/Y _19251_/Y _19405_/X vssd1 vssd1 vccd1 vccd1 _19412_/Y sky130_fd_sc_hd__a21boi_1
X_16624_ _16624_/A _16624_/B _16624_/C _16873_/B vssd1 vssd1 vccd1 vccd1 _16625_/C
+ sky130_fd_sc_hd__nand4_1
X_13836_ _13829_/B _13877_/A _13807_/A vssd1 vssd1 vccd1 vccd1 _13865_/A sky130_fd_sc_hd__o21ai_1
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17531__C _17833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _19343_/A _19343_/B _19343_/C vssd1 vssd1 vccd1 vccd1 _19530_/D sky130_fd_sc_hd__nand3_1
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16555_ _15638_/X _16312_/X _16313_/X _16296_/Y vssd1 vssd1 vccd1 vccd1 _16557_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13767_ _14110_/A vssd1 vssd1 vccd1 vccd1 _14181_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19897__A2 _18889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15506_ _15449_/X _15505_/X _15502_/C _15502_/D vssd1 vssd1 vccd1 vccd1 _15506_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_31_632 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19274_ _19268_/Y _19272_/X _19299_/C vssd1 vssd1 vccd1 vccd1 _19274_/Y sky130_fd_sc_hd__o21bai_2
XANTENNA__11641__A1 _11636_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ _12718_/A vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__buf_4
X_16486_ _17139_/A _17140_/A _16486_/C vssd1 vssd1 vccd1 vccd1 _16491_/B sky130_fd_sc_hd__nand3_2
XFILLER_188_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13698_ _22871_/Q vssd1 vssd1 vccd1 vccd1 _14506_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_176_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18225_ _12220_/A _12220_/B _12221_/A vssd1 vssd1 vccd1 vccd1 _18275_/B sky130_fd_sc_hd__a21oi_2
X_15437_ _15482_/A _16481_/B _15486_/A _12211_/A vssd1 vssd1 vccd1 vccd1 _16473_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12972__A _16100_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17109__B1 _11672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12649_ _12510_/A _12510_/B _12644_/Y _12645_/X vssd1 vssd1 vccd1 vccd1 _12651_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_178_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18156_ _18156_/A vssd1 vssd1 vccd1 vccd1 _18156_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__14591__B1 _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15368_ _15368_/A vssd1 vssd1 vccd1 vccd1 _15389_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17107_ _16976_/B _16934_/X _16944_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _17311_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_129_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11944__A2 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14319_ _22442_/B vssd1 vssd1 vccd1 vccd1 _14355_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18087_ _18087_/A _18087_/B vssd1 vssd1 vccd1 vccd1 _22968_/D sky130_fd_sc_hd__nand2_1
XFILLER_183_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15299_ _16256_/A _16256_/B _15299_/C _15299_/D vssd1 vssd1 vccd1 vccd1 _15309_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_171_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17038_ _17038_/A _17038_/B _17038_/C vssd1 vssd1 vccd1 vccd1 _17208_/A sky130_fd_sc_hd__nand3_4
XANTENNA__22405__A1 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14343__B1 _14337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22829__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18989_ _19002_/A _19002_/B vssd1 vssd1 vccd1 vccd1 _18990_/A sky130_fd_sc_hd__nand2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19490__A _19490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater133 _22693_/CLK vssd1 vssd1 vccd1 vccd1 _22696_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12212__A _15486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater144 _22803_/CLK vssd1 vssd1 vccd1 vccd1 _22765_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater155 _22746_/CLK vssd1 vssd1 vccd1 vccd1 _22747_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater166 _22800_/CLK vssd1 vssd1 vccd1 vccd1 _22768_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20951_ _20949_/B _20949_/C _20949_/A vssd1 vssd1 vccd1 vccd1 _20951_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20195__A2 _13045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11880__A1 _11877_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20882_ _20882_/A _20882_/B vssd1 vssd1 vccd1 vccd1 _20884_/C sky130_fd_sc_hd__xnor2_1
XFILLER_35_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19337__B2 _19336_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22621_ _22643_/A vssd1 vssd1 vccd1 vccd1 _22630_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22552_ _22768_/Q input42/X _22558_/S vssd1 vssd1 vccd1 vccd1 _22553_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11632__A1 _11644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21503_ _21504_/B _21504_/C _21504_/A vssd1 vssd1 vccd1 vccd1 _21649_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22483_ _22483_/A vssd1 vssd1 vccd1 vccd1 _22737_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16354__A _16354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21434_ _21292_/A _22673_/Q _21292_/C _13689_/A vssd1 vssd1 vccd1 vccd1 _21434_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_163_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21365_ _21365_/A _21365_/B vssd1 vssd1 vccd1 vccd1 _21372_/B sky130_fd_sc_hd__nand2_1
XFILLER_174_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20316_ _22930_/Q _20191_/B _20315_/Y vssd1 vssd1 vccd1 vccd1 _20317_/B sky130_fd_sc_hd__a21oi_2
XFILLER_190_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21296_ _21296_/A vssd1 vssd1 vccd1 vccd1 _22930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20247_ _15326_/X _15325_/X _20130_/C _16932_/C vssd1 vssd1 vccd1 vccd1 _20247_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11699__A1 _11644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20323__B _20323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20178_ _20178_/A vssd1 vssd1 vccd1 vccd1 _20843_/A sky130_fd_sc_hd__buf_2
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14321__B input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13218__A _21591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11664__C _18839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21368__D1 _13630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ _11859_/X _11861_/X _15714_/A vssd1 vssd1 vccd1 vccd1 _11951_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13860__A2 _13930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11961__A _12219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11871__A1 _18984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11882_ _16564_/B _19202_/D _11333_/X _11319_/Y vssd1 vssd1 vccd1 vccd1 _11883_/C
+ sky130_fd_sc_hd__a22o_1
X_14670_ _14670_/A vssd1 vssd1 vccd1 vccd1 _15213_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11871__B2 _18288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ _13617_/B _13602_/B _13620_/Y vssd1 vssd1 vccd1 vccd1 _13672_/B sky130_fd_sc_hd__o21ai_1
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22819_ _22929_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _22819_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19879__A2 _19294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16340_ _16311_/X _16314_/Y _16309_/Y _16301_/Y vssd1 vssd1 vccd1 vccd1 _16354_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_125_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13552_ _13552_/A vssd1 vssd1 vccd1 vccd1 _13677_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__12820__B1 _12687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12503_ _12503_/A _12503_/B vssd1 vssd1 vccd1 vccd1 _12621_/B sky130_fd_sc_hd__nand2_1
XFILLER_158_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16271_ _15580_/A _15933_/A _15557_/Y _16256_/Y _16258_/Y vssd1 vssd1 vccd1 vccd1
+ _16272_/C sky130_fd_sc_hd__o221ai_4
XFILLER_13_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13483_ _13501_/A _13550_/C _13477_/X vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__a21oi_1
XFILLER_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18010_ _17967_/A _22904_/Q _17967_/C _17970_/B _22903_/Q vssd1 vssd1 vccd1 vccd1
+ _18010_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_157_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15222_ _15224_/A _15224_/C _15224_/D _15224_/B vssd1 vssd1 vccd1 vccd1 _15223_/B
+ sky130_fd_sc_hd__o22ai_1
X_12434_ _12292_/A _15608_/C _12319_/Y vssd1 vssd1 vccd1 vccd1 _16779_/A sky130_fd_sc_hd__a21oi_4
XFILLER_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11926__A2 _11565_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15153_ _14871_/A _14871_/B _14942_/A _15122_/X _15124_/Y vssd1 vssd1 vccd1 vccd1
+ _15161_/A sky130_fd_sc_hd__a2111o_1
XANTENNA__15117__A2 _15006_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12365_ _12404_/A vssd1 vssd1 vccd1 vccd1 _20089_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11316_ _11316_/A _11316_/B vssd1 vssd1 vccd1 vccd1 _11790_/C sky130_fd_sc_hd__nand2_2
X_14104_ _14104_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14553_/B sky130_fd_sc_hd__nand2_2
X_19961_ _19962_/A _19962_/B _19962_/C vssd1 vssd1 vccd1 vccd1 _19963_/A sky130_fd_sc_hd__a21o_1
XFILLER_154_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15084_ _15081_/X _15107_/B _15107_/A _15083_/Y vssd1 vssd1 vccd1 vccd1 _15085_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ _22819_/Q vssd1 vssd1 vccd1 vccd1 _12411_/A sky130_fd_sc_hd__inv_2
XFILLER_181_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16711__B _20593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18912_ _18912_/A _18912_/B _18920_/B vssd1 vssd1 vccd1 vccd1 _18912_/X sky130_fd_sc_hd__and3_1
X_14035_ _14035_/A _14035_/B vssd1 vssd1 vccd1 vccd1 _14523_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19892_ _19892_/A _19892_/B vssd1 vssd1 vccd1 vccd1 _19893_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12887__B1 _16160_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14512__A _14512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18843_ _18843_/A _18843_/B vssd1 vssd1 vccd1 vccd1 _19161_/A sky130_fd_sc_hd__nand2_2
XFILLER_45_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21048__C _21048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18774_ _18774_/A _18774_/B _18774_/C _18774_/D vssd1 vssd1 vccd1 vccd1 _18774_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12639__B1 _12742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15986_ _16005_/A _16005_/B _16006_/A _16006_/B vssd1 vssd1 vccd1 vccd1 _15986_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12103__A2 _11626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17725_ _17611_/A _17611_/B _17708_/A _17708_/B vssd1 vssd1 vccd1 vccd1 _17790_/D
+ sky130_fd_sc_hd__a22oi_1
XFILLER_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14937_ _14872_/Y _15154_/D _14575_/B _14862_/Y vssd1 vssd1 vccd1 vccd1 _14937_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_57_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12967__A _12967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18357__C _18797_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17656_ _19768_/C vssd1 vssd1 vccd1 vccd1 _18305_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_91_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14868_ _15115_/A _14868_/B _14868_/C vssd1 vssd1 vccd1 vccd1 _14998_/C sky130_fd_sc_hd__nand3_1
XANTENNA__19319__A1 _12118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16607_ _16370_/B _16377_/B _16377_/C _16606_/X vssd1 vssd1 vccd1 vccd1 _16620_/B
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__15062__B _15114_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13819_ _14126_/A _13959_/A _13828_/B _14184_/C vssd1 vssd1 vccd1 vccd1 _13819_/Y
+ sky130_fd_sc_hd__nand4_2
X_17587_ _17479_/B _17470_/B _17479_/A vssd1 vssd1 vccd1 vccd1 _17590_/B sky130_fd_sc_hd__a21bo_1
XFILLER_51_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14799_ _14805_/C _14805_/D _14885_/B vssd1 vssd1 vccd1 vccd1 _14802_/B sky130_fd_sc_hd__a21o_1
X_19326_ _19326_/A vssd1 vssd1 vccd1 vccd1 _19521_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16538_ _16534_/A _16520_/A _16536_/B vssd1 vssd1 vccd1 vccd1 _16548_/A sky130_fd_sc_hd__a21o_1
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19469__A1_N _19476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15997__B _18984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22176__A _22176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18542__A2 _11474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19257_ _19257_/A _19257_/B _19257_/C vssd1 vssd1 vccd1 vccd1 _19257_/X sky130_fd_sc_hd__and3_1
XFILLER_149_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16469_ _16842_/A _16469_/B _16842_/C vssd1 vssd1 vccd1 vccd1 _16535_/B sky130_fd_sc_hd__and3_1
XANTENNA__17750__B1 _15840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18208_ _18208_/A _18208_/B vssd1 vssd1 vccd1 vccd1 _18216_/A sky130_fd_sc_hd__and2_1
XANTENNA__13367__A1 _13423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19188_ _19017_/Y _19026_/B _19014_/X _19015_/Y vssd1 vssd1 vccd1 vccd1 _19190_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18139_ _18340_/A vssd1 vssd1 vccd1 vccd1 _18139_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_176_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21150_ _21150_/A _21150_/B _21150_/C vssd1 vssd1 vccd1 vccd1 _21150_/Y sky130_fd_sc_hd__nand3_1
XFILLER_172_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11468__D _15901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20101_ _20101_/A _20101_/B _20101_/C vssd1 vssd1 vccd1 vccd1 _20110_/B sky130_fd_sc_hd__nand3_4
XFILLER_132_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21081_ _21082_/A _21081_/B _21081_/C _21081_/D vssd1 vssd1 vccd1 vccd1 _21088_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17436__C _17462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20032_ _22926_/Q _20032_/B _20032_/C vssd1 vssd1 vccd1 vccd1 _20033_/A sky130_fd_sc_hd__nor3_1
XANTENNA__21601__A2 _21594_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16695__B_N _22889_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11550__B1 _11895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17733__A _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21255__A _21990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21983_ _21983_/A _21983_/B _21983_/C vssd1 vssd1 vccd1 vccd1 _21994_/A sky130_fd_sc_hd__nand3_1
XFILLER_66_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20934_ _20924_/X _20926_/X _20937_/A _20933_/Y vssd1 vssd1 vccd1 vccd1 _20934_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ _20860_/B _20860_/C _20793_/Y vssd1 vssd1 vccd1 vccd1 _20865_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22604_ _18115_/A input64/X _22608_/S vssd1 vssd1 vccd1 vccd1 _22605_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20796_ _20796_/A _20796_/B vssd1 vssd1 vccd1 vccd1 _20797_/D sky130_fd_sc_hd__nand2_1
XFILLER_195_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22535_ _22535_/A vssd1 vssd1 vccd1 vccd1 _22760_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16544__A1 _16155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16515__C _18193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22617__A1 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14555__B1 _14843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22466_ _22512_/S vssd1 vssd1 vccd1 vccd1 _22475_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21417_ _21553_/A _21417_/B _21417_/C vssd1 vssd1 vccd1 vccd1 _21440_/A sky130_fd_sc_hd__nand3_2
XFILLER_120_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12117__A _12117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22397_ _22397_/A vssd1 vssd1 vccd1 vccd1 _22699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12150_ _18116_/D _18128_/A vssd1 vssd1 vccd1 vccd1 _18339_/A sky130_fd_sc_hd__nand2_2
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21348_ _21348_/A vssd1 vssd1 vccd1 vccd1 _21460_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11956__A _19016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15428__A _15718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _12081_/A vssd1 vssd1 vccd1 vccd1 _12081_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21279_ _21264_/Y _21267_/X _21276_/C vssd1 vssd1 vccd1 vccd1 _21282_/A sky130_fd_sc_hd__o21ai_1
XFILLER_78_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19797__A1 _19615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _15840_/A vssd1 vssd1 vccd1 vccd1 _15840_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__17643__A _17643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17009__C1 _17008_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16480__B1 _16513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15771_ _15350_/Y _15646_/X _15389_/C _15389_/A vssd1 vssd1 vccd1 vccd1 _16402_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12983_ _12989_/A _12989_/B _12989_/C vssd1 vssd1 vccd1 vccd1 _12990_/A sky130_fd_sc_hd__a21o_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16259__A _19016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17510_ _17616_/B _17616_/C _17616_/A _17719_/A _17719_/C vssd1 vssd1 vccd1 vccd1
+ _17511_/B sky130_fd_sc_hd__o32a_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14722_ _14722_/A _14808_/D _14722_/C vssd1 vssd1 vccd1 vccd1 _14722_/Y sky130_fd_sc_hd__nand3_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _19316_/A vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__clkbuf_4
X_18490_ _18490_/A _18490_/B _18490_/C vssd1 vssd1 vccd1 vccd1 _18491_/A sky130_fd_sc_hd__nand3_1
XFILLER_40_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _17442_/A _17439_/X _17110_/B _17880_/A _16015_/X vssd1 vssd1 vccd1 vccd1
+ _17441_/X sky130_fd_sc_hd__o32a_1
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13046__B1 _13045_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14653_ _14656_/C _14656_/B vssd1 vssd1 vccd1 vccd1 _14655_/A sky130_fd_sc_hd__nand2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _16712_/C vssd1 vssd1 vccd1 vccd1 _17085_/C sky130_fd_sc_hd__buf_4
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output106_A _14428_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _13565_/Y _13524_/X _13526_/X vssd1 vssd1 vccd1 vccd1 _13604_/X sky130_fd_sc_hd__a21o_1
X_17372_ _17372_/A _17372_/B _17372_/C vssd1 vssd1 vccd1 vccd1 _17507_/A sky130_fd_sc_hd__nand3_2
XFILLER_186_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11796_ _11796_/A _18328_/B _18328_/C vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__and3_1
X_14584_ _22764_/Q vssd1 vssd1 vccd1 vccd1 _14863_/A sky130_fd_sc_hd__inv_2
XFILLER_186_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19111_ _19111_/A _19116_/B vssd1 vssd1 vccd1 vccd1 _19122_/B sky130_fd_sc_hd__nand2_1
XFILLER_158_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16323_ _16323_/A _16323_/B _16323_/C _16323_/D vssd1 vssd1 vccd1 vccd1 _16324_/B
+ sky130_fd_sc_hd__nand4_4
X_13535_ _13460_/A _13460_/B _13533_/Y _13534_/Y _13455_/Y vssd1 vssd1 vccd1 vccd1
+ _13538_/B sky130_fd_sc_hd__o221ai_1
XFILLER_185_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22674__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13349__A1 _21383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19042_ _19418_/A _19504_/B _19504_/C _19202_/D vssd1 vssd1 vccd1 vccd1 _19065_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_173_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16254_ _16530_/D _16530_/A _15542_/X _16253_/Y vssd1 vssd1 vccd1 vccd1 _16288_/C
+ sky130_fd_sc_hd__o2bb2ai_4
XANTENNA__22608__A1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13466_ _13461_/Y _13463_/Y _13464_/X _13465_/Y vssd1 vssd1 vccd1 vccd1 _13470_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_167_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21050__D _21050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14226__B _15114_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15205_ _15205_/A _15205_/B _15205_/C vssd1 vssd1 vccd1 vccd1 _15206_/B sky130_fd_sc_hd__and3_1
XFILLER_138_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12417_ _16465_/A _12967_/A _20255_/C _12701_/A _12921_/A vssd1 vssd1 vccd1 vccd1
+ _12417_/X sky130_fd_sc_hd__o32a_1
XANTENNA__19485__B1 _19340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17818__A _18814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16185_ _16186_/A _16184_/Y _16181_/X vssd1 vssd1 vccd1 vccd1 _16185_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13397_ _13484_/B _13289_/A _13396_/X vssd1 vssd1 vccd1 vccd1 _13399_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__16838__A2 _16825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15136_ _15095_/A _15095_/B _15095_/C _15135_/A _15135_/B vssd1 vssd1 vccd1 vccd1
+ _15136_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_126_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12348_ _12348_/A vssd1 vssd1 vccd1 vccd1 _20341_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_154_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11866__A _18985_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19944_ _19981_/A _19987_/D _17872_/C _19901_/C vssd1 vssd1 vccd1 vccd1 _19946_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15067_ _15060_/X _15066_/Y _14996_/B vssd1 vssd1 vccd1 vccd1 _15073_/C sky130_fd_sc_hd__o21ai_1
X_12279_ _12300_/A _12279_/B _15363_/C vssd1 vssd1 vccd1 vccd1 _12607_/A sky130_fd_sc_hd__nand3_2
XANTENNA__16160__C _16160_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14018_ _14014_/X _14026_/B _14017_/X vssd1 vssd1 vccd1 vccd1 _14169_/C sky130_fd_sc_hd__o21ai_1
X_19875_ _19875_/A _19919_/A vssd1 vssd1 vccd1 vccd1 _19881_/C sky130_fd_sc_hd__or2b_1
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18460__A1 _12204_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18826_ _18826_/A _18826_/B vssd1 vssd1 vccd1 vccd1 _18827_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18460__B2 _11566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19471__C _19476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15274__A1 _22877_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18757_ _18645_/Y _18646_/X _18725_/X _18732_/Y _18737_/X vssd1 vssd1 vccd1 vccd1
+ _18757_/X sky130_fd_sc_hd__o221a_1
X_15969_ _15824_/A _15824_/B _15824_/C vssd1 vssd1 vccd1 vccd1 _15970_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12697__A _12697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17708_ _17708_/A _17708_/B vssd1 vssd1 vccd1 vccd1 _17708_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17015__A2 _17008_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18688_ _18691_/A _18691_/B _18690_/B vssd1 vssd1 vccd1 vccd1 _18877_/A sky130_fd_sc_hd__nand3_1
XANTENNA__20555__C1 _20551_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ _17633_/Y _17637_/Y _17638_/X vssd1 vssd1 vccd1 vccd1 _17661_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__13305__B _13305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16774__A1 _12571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16774__B2 _15541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20650_ _20650_/A _20650_/B _20650_/C vssd1 vssd1 vccd1 vccd1 _20652_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19199__B _19199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13024__C _15746_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19309_ _19329_/A vssd1 vssd1 vccd1 vccd1 _19618_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20581_ _20581_/A _20581_/B vssd1 vssd1 vccd1 vccd1 _20586_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22320_ _22320_/A vssd1 vssd1 vccd1 vccd1 _22341_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22251_ _22294_/A _22251_/B vssd1 vssd1 vccd1 vccd1 _22253_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17728__A _17728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21202_ _21202_/A _21301_/A vssd1 vssd1 vccd1 vccd1 _21202_/Y sky130_fd_sc_hd__nor2_2
XFILLER_133_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22182_ _22182_/A _22182_/B _22182_/C vssd1 vssd1 vccd1 vccd1 _22186_/B sky130_fd_sc_hd__nand3_1
XFILLER_2_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13975__B _14963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11776__A _19197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21133_ _20834_/X _20835_/X _21135_/A _21118_/C vssd1 vssd1 vccd1 vccd1 _21133_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_133_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21064_ _21067_/A _21067_/B _21067_/C _21067_/D vssd1 vssd1 vccd1 vccd1 _21079_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_154_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11523__B1 _11295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20389__A2 _20381_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20574__A2_N _20637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20015_ _19949_/A _19949_/B _19988_/X _20037_/B vssd1 vssd1 vccd1 vccd1 _20016_/B
+ sky130_fd_sc_hd__o31ai_1
XFILLER_171_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17254__A2 _17391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15265__A1 _14845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16462__B1 _16452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18278__B _18278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18739__C1 _18666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11942__C _18107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21966_ _21957_/A _22037_/C _22220_/A _21965_/Y _22031_/A vssd1 vssd1 vccd1 vccd1
+ _21972_/C sky130_fd_sc_hd__o2111ai_4
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _20917_/A _20917_/B vssd1 vssd1 vccd1 vccd1 _20917_/Y sky130_fd_sc_hd__nand2_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ _21897_/A _21897_/B vssd1 vssd1 vccd1 vccd1 _21901_/A sky130_fd_sc_hd__xnor2_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15711__A _15711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11650_ _11507_/X _11501_/Y _11493_/Y vssd1 vssd1 vccd1 vccd1 _11674_/A sky130_fd_sc_hd__a21boi_2
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ _20920_/A _20848_/B vssd1 vssd1 vccd1 vccd1 _20848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_888 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11581_ _11581_/A _11789_/A vssd1 vssd1 vccd1 vccd1 _11589_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20779_ _15941_/A _20123_/X _17444_/A _20682_/C vssd1 vssd1 vccd1 vccd1 _20871_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17714__B1 _22900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13320_ _21495_/C _21495_/A vssd1 vssd1 vccd1 vccd1 _21318_/A sky130_fd_sc_hd__nand2_2
XFILLER_196_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15725__C1 _19154_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22518_ _22518_/A vssd1 vssd1 vccd1 vccd1 _22752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19467__B1 _15810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22449_ _13257_/B input57/X _22453_/S vssd1 vssd1 vccd1 vccd1 _22450_/A sky130_fd_sc_hd__mux2_1
X_13251_ _21367_/C vssd1 vssd1 vccd1 vccd1 _21629_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_171_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12202_ _12202_/A _12202_/B vssd1 vssd1 vccd1 vccd1 _19587_/C sky130_fd_sc_hd__nand2_4
XANTENNA__12554__A2 _12773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13182_ _22735_/Q vssd1 vssd1 vccd1 vccd1 _21473_/A sky130_fd_sc_hd__inv_2
XFILLER_182_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input67_A wb_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21813__A2 _21677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16261__B _16261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12133_ _18348_/A _12135_/A _12135_/B vssd1 vssd1 vccd1 vccd1 _12134_/B sky130_fd_sc_hd__and3_1
X_17990_ _17989_/A _17991_/A _17989_/C vssd1 vssd1 vccd1 vccd1 _18062_/C sky130_fd_sc_hd__a21o_1
XFILLER_151_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16941_ _16941_/A vssd1 vssd1 vccd1 vccd1 _16941_/X sky130_fd_sc_hd__clkbuf_2
X_12064_ _12064_/A vssd1 vssd1 vccd1 vccd1 _12064_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17373__A _17373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19660_ _19432_/Y _19565_/Y _19439_/B _19659_/Y vssd1 vssd1 vccd1 vccd1 _19813_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_49_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16872_ _16873_/C _16873_/D _16869_/B vssd1 vssd1 vccd1 vccd1 _16874_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20511__B _20511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18611_ _12170_/X _12171_/X _17380_/X _17381_/A _18200_/A vssd1 vssd1 vccd1 vccd1
+ _18611_/Y sky130_fd_sc_hd__o221ai_4
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ _15823_/A _16106_/D _19614_/A vssd1 vssd1 vccd1 vccd1 _15824_/C sky130_fd_sc_hd__and3_1
Xclkbuf_3_2_0_bq_clk_i clkbuf_3_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19591_ _19596_/B _19596_/C _19590_/X vssd1 vssd1 vccd1 vccd1 _19591_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_65_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _17434_/A _11474_/X _18536_/Y _18537_/X _18664_/B vssd1 vssd1 vccd1 vccd1
+ _18543_/C sky130_fd_sc_hd__o221ai_4
XFILLER_92_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15752_/X _15753_/Y _15864_/A _15709_/Y vssd1 vssd1 vccd1 vccd1 _15864_/B
+ sky130_fd_sc_hd__o211ai_4
X_12966_ _12966_/A _12966_/B _12966_/C vssd1 vssd1 vccd1 vccd1 _13011_/C sky130_fd_sc_hd__nand3_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _14868_/B vssd1 vssd1 vccd1 vccd1 _15115_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__19942__B2 _19896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ _18770_/C _18461_/B _18465_/X _18467_/Y _18462_/A vssd1 vssd1 vccd1 vccd1
+ _18473_/Y sky130_fd_sc_hd__o221ai_2
X_11917_ _18830_/A _16106_/B _18629_/A _12065_/A vssd1 vssd1 vccd1 vccd1 _11918_/B
+ sky130_fd_sc_hd__and4_1
X_15685_ _15682_/A _15433_/A _15684_/Y vssd1 vssd1 vccd1 vccd1 _15766_/A sky130_fd_sc_hd__a21oi_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1054 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16717__A _18716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20552__A2 _20065_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12897_ _12741_/C _12741_/A _12741_/B _13007_/B _12750_/B vssd1 vssd1 vccd1 vccd1
+ _12900_/A sky130_fd_sc_hd__a32oi_1
XFILLER_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ _17424_/A vssd1 vssd1 vccd1 vccd1 _17424_/X sky130_fd_sc_hd__buf_2
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _14740_/A _14636_/B _14636_/C _14636_/D vssd1 vssd1 vccd1 vccd1 _14740_/B
+ sky130_fd_sc_hd__nand4_2
X_11848_ _15714_/B vssd1 vssd1 vccd1 vccd1 _19329_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_127_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16436__B _20069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15978__D _17645_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17230_/Y _17353_/X _17354_/Y vssd1 vssd1 vccd1 vccd1 _17372_/C sky130_fd_sc_hd__o21ai_2
XFILLER_14_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16508__A1 _12716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14567_ _15058_/A _15058_/B _14693_/D vssd1 vssd1 vccd1 vccd1 _14568_/B sky130_fd_sc_hd__nand3_1
XANTENNA__17166__D1 _19772_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11779_ _18107_/A _11779_/B _11779_/C vssd1 vssd1 vccd1 vccd1 _11779_/X sky130_fd_sc_hd__and3_1
XFILLER_147_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16306_ _20605_/A vssd1 vssd1 vccd1 vccd1 _20608_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__13141__A _13141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19170__A2 _17422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13518_ _21173_/A _13521_/B _21173_/C vssd1 vssd1 vccd1 vccd1 _13520_/A sky130_fd_sc_hd__nand3_1
X_17286_ _11561_/X _11563_/X _16737_/A vssd1 vssd1 vccd1 vccd1 _17286_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14498_ _14492_/Y _14611_/B _14497_/Y vssd1 vssd1 vccd1 vccd1 _14498_/Y sky130_fd_sc_hd__a21oi_1
X_19025_ _19461_/A _19496_/B _19496_/C vssd1 vssd1 vccd1 vccd1 _19026_/B sky130_fd_sc_hd__and3_1
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ _15589_/X _16474_/A _16221_/Y _19047_/B _15991_/B vssd1 vssd1 vccd1 vccd1
+ _16532_/A sky130_fd_sc_hd__o2111ai_4
X_13449_ _13449_/A _13449_/B _21312_/B vssd1 vssd1 vccd1 vccd1 _13461_/A sky130_fd_sc_hd__nand3_2
XFILLER_173_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12980__A _15774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22173__B _22173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16168_ _16168_/A _16168_/B vssd1 vssd1 vccd1 vccd1 _16168_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15068__A _15114_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15119_ _15186_/A _15119_/B _15119_/C _15119_/D vssd1 vssd1 vccd1 vccd1 _15120_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_170_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16099_ _13022_/D _16098_/X _13022_/A _15887_/X vssd1 vssd1 vccd1 vccd1 _16099_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_134_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19927_ _19878_/Y _19880_/Y _19750_/X vssd1 vssd1 vccd1 vccd1 _19928_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__19482__B _20012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17236__A2 _17379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17283__A _19615_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19858_ _19913_/B _19860_/C _19860_/A vssd1 vssd1 vccd1 vccd1 _19859_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__14700__A _22765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18809_ _18824_/A _18824_/B _18824_/C vssd1 vssd1 vccd1 vccd1 _19079_/A sky130_fd_sc_hd__nand3_2
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22517__A0 _14220_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19789_ _19789_/A _19789_/B vssd1 vssd1 vccd1 vccd1 _19796_/C sky130_fd_sc_hd__nand2_1
XANTENNA__15798__A2 _15797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20791__A2 _17435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21820_ _21820_/A vssd1 vssd1 vccd1 vccd1 _22089_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12220__A _12220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11762__C _11932_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21751_ _21751_/A _21751_/B vssd1 vssd1 vccd1 vccd1 _21758_/D sky130_fd_sc_hd__nand2_1
XANTENNA__16747__A1 _15932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16627__A _16627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15531__A _15531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20702_ _20702_/A _20702_/B _20702_/C _20702_/D vssd1 vssd1 vccd1 vccd1 _20720_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_180_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21682_ _21809_/A _21686_/A _21687_/C vssd1 vssd1 vccd1 vccd1 _21688_/A sky130_fd_sc_hd__a21o_1
XFILLER_196_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20633_ _20602_/Y _20603_/X _20630_/A vssd1 vssd1 vccd1 vccd1 _20738_/B sky130_fd_sc_hd__o21ai_1
XFILLER_138_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14147__A _14147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13981__A1 _14122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20564_ _20564_/A _20564_/B vssd1 vssd1 vccd1 vccd1 _22913_/D sky130_fd_sc_hd__xnor2_4
XFILLER_138_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22303_ _22304_/B _22304_/C _22186_/A _22308_/B vssd1 vssd1 vccd1 vccd1 _22306_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_165_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20495_ _20495_/A _20495_/B vssd1 vssd1 vccd1 vccd1 _20495_/Y sky130_fd_sc_hd__nand2_1
XFILLER_192_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22234_ _22271_/A _22271_/B vssd1 vssd1 vccd1 vccd1 _22237_/A sky130_fd_sc_hd__xor2_1
XFILLER_145_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22165_ _22080_/B _22163_/Y _22159_/B _22164_/Y vssd1 vssd1 vccd1 vccd1 _22165_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21116_ _20834_/X _20835_/X _21115_/Y _21079_/Y vssd1 vssd1 vccd1 vccd1 _21118_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_120_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22096_ _22290_/A _22290_/B vssd1 vssd1 vccd1 vccd1 _22096_/X sky130_fd_sc_hd__and2_1
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15706__A _15706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21047_ _21011_/B _17839_/B _17839_/C _21082_/A _21082_/C vssd1 vssd1 vccd1 vccd1
+ _21053_/A sky130_fd_sc_hd__a311o_1
XFILLER_87_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15789__A2 _12576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12820_ _16778_/A _16779_/A _12687_/B vssd1 vssd1 vccd1 vccd1 _12820_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_74_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21443__A _21522_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12487__D _20486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _13007_/C _12751_/B vssd1 vssd1 vccd1 vccd1 _12895_/B sky130_fd_sc_hd__nand2_1
XFILLER_188_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21949_ _21758_/C _21882_/A _21947_/Y _21948_/X vssd1 vssd1 vccd1 vccd1 _22036_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15441__A _17234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11702_ _11702_/A vssd1 vssd1 vccd1 vccd1 _11702_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15477_/A _15470_/B vssd1 vssd1 vccd1 vccd1 _15474_/A sky130_fd_sc_hd__nand2_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12682_ _12689_/A _17401_/B _12680_/X _12681_/X vssd1 vssd1 vccd1 vccd1 _12682_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__15410__A1 _11911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15410__B2 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16256__B _16256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14421_ _22812_/Q _14411_/X _14412_/X _14413_/X _22780_/Q vssd1 vssd1 vccd1 vccd1
+ _14421_/X sky130_fd_sc_hd__a32o_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11633_ _11633_/A vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17140_ _17140_/A vssd1 vssd1 vccd1 vccd1 _17532_/D sky130_fd_sc_hd__buf_2
XFILLER_129_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14352_ _21188_/B vssd1 vssd1 vccd1 vccd1 _21329_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12775__A2 _12774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11564_ _11468_/Y _18371_/A _11452_/X vssd1 vssd1 vccd1 vccd1 _11565_/B sky130_fd_sc_hd__o21ai_1
XFILLER_11_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18360__B1 _11345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13896__A _13896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ _13301_/X _21336_/B _21584_/C _13079_/A vssd1 vssd1 vccd1 vccd1 _13305_/A
+ sky130_fd_sc_hd__o211ai_4
X_17071_ _17071_/A _17071_/B _17071_/C vssd1 vssd1 vccd1 vccd1 _17073_/A sky130_fd_sc_hd__and3_1
XFILLER_144_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11495_ _11792_/A vssd1 vssd1 vccd1 vccd1 _18131_/B sky130_fd_sc_hd__buf_2
X_14283_ _14243_/A _14250_/Y _14253_/Y _14281_/Y _14282_/Y vssd1 vssd1 vccd1 vccd1
+ _14283_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_183_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16022_ _15967_/X _15971_/Y _16020_/Y _16021_/Y vssd1 vssd1 vccd1 vccd1 _16024_/A
+ sky130_fd_sc_hd__o211ai_2
X_13234_ _13234_/A _13234_/B _13234_/C vssd1 vssd1 vccd1 vccd1 _13504_/C sky130_fd_sc_hd__and3_1
XFILLER_171_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19583__A _19689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ _13384_/A _13384_/B _13385_/A vssd1 vssd1 vccd1 vccd1 _13286_/D sky130_fd_sc_hd__nand3_1
XFILLER_151_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12116_ _12116_/A vssd1 vssd1 vccd1 vccd1 _12116_/X sky130_fd_sc_hd__buf_2
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17973_ _18020_/A _18020_/B _18020_/C vssd1 vssd1 vccd1 vccd1 _17997_/A sky130_fd_sc_hd__nor3_1
X_13096_ _13096_/A vssd1 vssd1 vccd1 vccd1 _13099_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_123_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19712_ _19602_/Y _19603_/X _19685_/X _19684_/X vssd1 vssd1 vccd1 vccd1 _19712_/X
+ sky130_fd_sc_hd__a31o_1
X_12047_ _22658_/B _12046_/X _22660_/B _11721_/C vssd1 vssd1 vccd1 vccd1 _16477_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15616__A _15616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16924_ _20675_/A vssd1 vssd1 vccd1 vccd1 _17386_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21014__A3 _21044_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19643_ _19536_/A _19637_/Y _19635_/A _19724_/B vssd1 vssd1 vccd1 vccd1 _19643_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_172_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16855_ _16605_/B _16624_/A _16624_/B vssd1 vssd1 vccd1 vccd1 _16860_/A sky130_fd_sc_hd__a21boi_2
XANTENNA__16977__A1 _15545_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13781__D _15008_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16977__B2 _16944_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15806_ _15810_/A _15810_/B _16106_/A _15804_/Y _15805_/Y vssd1 vssd1 vccd1 vccd1
+ _15824_/A sky130_fd_sc_hd__a32o_1
XFILLER_19_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19574_ _19574_/A _19574_/B _19574_/C vssd1 vssd1 vccd1 vccd1 _19575_/B sky130_fd_sc_hd__and3_1
XANTENNA__14988__B1 _15046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__A _22962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16786_ _16786_/A vssd1 vssd1 vccd1 vccd1 _17634_/A sky130_fd_sc_hd__buf_2
XFILLER_168_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13998_ _13998_/A _13998_/B _13998_/C vssd1 vssd1 vccd1 vccd1 _14497_/A sky130_fd_sc_hd__nand3_2
XANTENNA__14452__A2 _11404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18525_ _18345_/A _18345_/B _18345_/C _18520_/B _18520_/A vssd1 vssd1 vccd1 vccd1
+ _18527_/B sky130_fd_sc_hd__a32oi_4
X_15737_ _15860_/A _15859_/C _15859_/D vssd1 vssd1 vccd1 vccd1 _15758_/A sky130_fd_sc_hd__nand3_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12949_ _20579_/C vssd1 vssd1 vccd1 vccd1 _12981_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16447__A _16447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18456_ _18455_/Y _18296_/B _18289_/Y vssd1 vssd1 vccd1 vccd1 _18458_/B sky130_fd_sc_hd__o21ai_2
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15668_ _15668_/A vssd1 vssd1 vccd1 vccd1 _15668_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17407_ _17407_/A _18303_/A _18303_/B vssd1 vssd1 vccd1 vccd1 _17408_/B sky130_fd_sc_hd__and3_1
XFILLER_33_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17941__A3 _17981_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14619_ _14619_/A vssd1 vssd1 vccd1 vccd1 _14619_/X sky130_fd_sc_hd__clkbuf_2
X_18387_ _18387_/A _18387_/B _18387_/C vssd1 vssd1 vccd1 vccd1 _18388_/A sky130_fd_sc_hd__and3_1
XFILLER_53_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15599_ _15510_/B _15672_/A _15672_/B vssd1 vssd1 vccd1 vccd1 _15678_/B sky130_fd_sc_hd__nand3b_1
XFILLER_18_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17338_ _17103_/C _17338_/B vssd1 vssd1 vccd1 vccd1 _17338_/X sky130_fd_sc_hd__and2b_1
XFILLER_105_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17269_ _17269_/A _17269_/B vssd1 vssd1 vccd1 vccd1 _17272_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16362__C1 _16586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19008_ _19001_/Y _19002_/Y _19007_/Y vssd1 vssd1 vccd1 vccd1 _19009_/D sky130_fd_sc_hd__o21ai_1
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16613__C _16613_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20280_ _20281_/B _20284_/C _20281_/A vssd1 vssd1 vccd1 vccd1 _20280_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14430__A _14430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22921_ _22922_/CLK _22921_/D vssd1 vssd1 vccd1 vccd1 _22921_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16968__B2 _15934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21961__A1 _21376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17090__B1 _16997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22852_ _22944_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 _22852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15640__A1 _15891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21803_ _21803_/A _21803_/B _21803_/C vssd1 vssd1 vccd1 vccd1 _21804_/A sky130_fd_sc_hd__nand3_1
X_22783_ _22803_/CLK _22783_/D vssd1 vssd1 vccd1 vccd1 _22783_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12885__A _16157_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21734_ _21963_/A _21219_/C _21633_/Y _21733_/X vssd1 vssd1 vccd1 vccd1 _21737_/A
+ sky130_fd_sc_hd__a31o_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21665_ _21713_/C _21713_/A _21805_/D _21665_/D vssd1 vssd1 vccd1 vccd1 _21665_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_40_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20616_ _20241_/A _15723_/A _15938_/A _20611_/Y _20606_/Y vssd1 vssd1 vccd1 vccd1
+ _20616_/X sky130_fd_sc_hd__o221a_1
X_21596_ _21596_/A _21596_/B vssd1 vssd1 vccd1 vccd1 _21758_/A sky130_fd_sc_hd__nand2_2
XFILLER_32_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15156__B1 _15188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20547_ _20539_/Y _20543_/Y _20546_/Y vssd1 vssd1 vccd1 vccd1 _20547_/X sky130_fd_sc_hd__o21a_2
XFILLER_4_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11280_ _22784_/Q _11374_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11860_/A sky130_fd_sc_hd__o21ai_2
X_20478_ _20579_/A _20579_/B _20478_/C vssd1 vssd1 vccd1 vccd1 _20482_/B sky130_fd_sc_hd__nand3_2
XFILLER_118_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17916__A _22903_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22217_ _22170_/A _22170_/B _22194_/B vssd1 vssd1 vccd1 vccd1 _22217_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_193_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22885__CLK _22922_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22148_ _22212_/A _22156_/A _22156_/B _22284_/C vssd1 vssd1 vccd1 vccd1 _22150_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_161_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15436__A _22961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22079_ _22075_/X _22079_/B _22079_/C vssd1 vssd1 vccd1 vccd1 _22080_/C sky130_fd_sc_hd__nand3b_1
X_14970_ _14971_/C _14971_/A _14971_/B vssd1 vssd1 vccd1 vccd1 _14970_/X sky130_fd_sc_hd__a21o_1
XFILLER_75_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18948__A2 _19983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13921_ _14021_/C _14021_/D _13916_/Y vssd1 vssd1 vccd1 vccd1 _13921_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19070__B2 _19091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16640_ _17431_/C vssd1 vssd1 vccd1 vccd1 _20972_/B sky130_fd_sc_hd__buf_2
XANTENNA__17651__A _19689_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13852_ _22869_/Q vssd1 vssd1 vccd1 vccd1 _14777_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_90_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20008__C_N _22925_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ _12803_/A vssd1 vssd1 vccd1 vccd1 _12803_/X sky130_fd_sc_hd__buf_2
XFILLER_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16571_ _22702_/Q vssd1 vssd1 vccd1 vccd1 _16571_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13783_ _14079_/A _14489_/B _13765_/X _14043_/B _13784_/A vssd1 vssd1 vccd1 vccd1
+ _14165_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_43_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18310_ _18310_/A _18310_/B vssd1 vssd1 vccd1 vccd1 _18310_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15522_ _15522_/A vssd1 vssd1 vccd1 vccd1 _15522_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18185__C _18279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19290_ _19290_/A _19290_/B _19290_/C vssd1 vssd1 vccd1 vccd1 _19292_/A sky130_fd_sc_hd__and3_1
X_12734_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12734_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18241_ _18249_/B _18241_/B vssd1 vssd1 vccd1 vccd1 _18772_/A sky130_fd_sc_hd__nand2_2
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15453_ _11820_/A _15450_/X _15452_/Y vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__o21ai_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12665_ _12665_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _12898_/C sky130_fd_sc_hd__nor2_1
XFILLER_169_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18482__A _18482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _22806_/Q _14397_/X _14398_/X _14391_/X _22774_/Q vssd1 vssd1 vccd1 vccd1
+ _14404_/X sky130_fd_sc_hd__a32o_1
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18172_ _18172_/A _18383_/B _18310_/A _18310_/B vssd1 vssd1 vccd1 vccd1 _18173_/C
+ sky130_fd_sc_hd__nand4_4
X_11616_ _11616_/A _11616_/B _11616_/C vssd1 vssd1 vccd1 vccd1 _11974_/A sky130_fd_sc_hd__nand3_2
XANTENNA__17136__A1 _12735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15384_ _15386_/A _15384_/B _15384_/C vssd1 vssd1 vccd1 vccd1 _15385_/A sky130_fd_sc_hd__nand3b_1
XFILLER_196_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12596_ _12596_/A vssd1 vssd1 vccd1 vccd1 _12697_/A sky130_fd_sc_hd__clkbuf_4
X_17123_ _16911_/X _16913_/X _16926_/B _16915_/Y vssd1 vssd1 vccd1 vccd1 _17123_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_14335_ _11349_/X _14317_/X _14320_/X _14334_/X _13826_/C vssd1 vssd1 vccd1 vccd1
+ _14335_/X sky130_fd_sc_hd__a32o_2
XANTENNA__18884__A1 _15932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11547_ _11553_/B _11552_/B _11552_/A vssd1 vssd1 vccd1 vccd1 _11547_/Y sky130_fd_sc_hd__nand3_1
XFILLER_184_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_362 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20691__A1 _20110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17054_ _17049_/Y _17050_/X _17053_/Y vssd1 vssd1 vccd1 vccd1 _17054_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_144_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14266_ _14267_/A _14267_/B _14267_/C vssd1 vssd1 vccd1 vccd1 _14269_/C sky130_fd_sc_hd__a21o_1
X_11478_ _11893_/B vssd1 vssd1 vccd1 vccd1 _11895_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__11708__B1 _11704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16005_ _16005_/A _16005_/B vssd1 vssd1 vccd1 vccd1 _16045_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13217_ _21480_/B vssd1 vssd1 vccd1 vccd1 _21591_/B sky130_fd_sc_hd__buf_2
X_14197_ _14197_/A _14197_/B vssd1 vssd1 vccd1 vccd1 _14255_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13148_ _22844_/Q vssd1 vssd1 vccd1 vccd1 _21609_/B sky130_fd_sc_hd__clkbuf_2
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15991__D _15991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15346__A _15633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17956_ _17919_/C _17954_/X _17908_/Y _17955_/Y vssd1 vssd1 vccd1 vccd1 _17958_/A
+ sky130_fd_sc_hd__o22ai_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _13079_/A _13304_/A vssd1 vssd1 vccd1 vccd1 _21351_/A sky130_fd_sc_hd__nand2_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12689__B _17401_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16907_ _16846_/B _16846_/C _16846_/A _16866_/C _16866_/D vssd1 vssd1 vccd1 vccd1
+ _16907_/Y sky130_fd_sc_hd__a32oi_2
X_17887_ _17886_/A _17886_/B _17886_/C vssd1 vssd1 vccd1 vccd1 _17888_/B sky130_fd_sc_hd__a21o_1
XANTENNA__20746__A2 _20734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19626_ _16015_/X _19941_/D _19793_/A _19476_/C vssd1 vssd1 vccd1 vccd1 _19626_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16838_ _16451_/B _16825_/X _16828_/A _16828_/B _16452_/X vssd1 vssd1 vccd1 vccd1
+ _16845_/D sky130_fd_sc_hd__o2111ai_2
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15622__A1 _11911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15622__B2 _15378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21083__A _21083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12436__A1 _16778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19557_ _12064_/X _19306_/X _18023_/X _19211_/A _19411_/X vssd1 vssd1 vccd1 vccd1
+ _19557_/X sky130_fd_sc_hd__o311a_1
X_16769_ _16506_/X _16507_/X _16489_/X _16496_/X vssd1 vssd1 vccd1 vccd1 _16776_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_19_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16177__A _16177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19364__A2 _17526_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18508_ _18508_/A _18508_/B vssd1 vssd1 vccd1 vccd1 _18508_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12987__A2 _20452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19488_ _19488_/A _19636_/A _19636_/B vssd1 vssd1 vccd1 vccd1 _19536_/B sky130_fd_sc_hd__nand3_1
XFILLER_55_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1018 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18439_ _18427_/X _18428_/Y _18773_/A vssd1 vssd1 vccd1 vccd1 _18774_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__16583__C1 _16324_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21450_ _21365_/B _21633_/A _21449_/Y vssd1 vssd1 vccd1 vccd1 _21450_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20401_ _20401_/A _20401_/B vssd1 vssd1 vccd1 vccd1 _20401_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19000__B _19161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21381_ _21247_/A _21247_/B _21380_/Y vssd1 vssd1 vccd1 vccd1 _21535_/B sky130_fd_sc_hd__a21oi_1
XFILLER_179_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15689__A1 _12968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15689__B2 _12118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20332_ _20206_/Y _20364_/A _20447_/A _20447_/B vssd1 vssd1 vccd1 vccd1 _20335_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_190_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17736__A _17736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18627__A1 _15538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20263_ _20263_/A _20263_/B vssd1 vssd1 vccd1 vccd1 _20390_/D sky130_fd_sc_hd__nand2_2
XFILLER_89_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16640__A _17431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22002_ _21993_/A _22029_/B _21996_/A _21996_/B vssd1 vssd1 vccd1 vccd1 _22002_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__20434__A1 _20553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16638__B1 _16630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12911__A2 _16078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16102__A2 _20452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20194_ _13044_/A _13044_/B _12754_/X vssd1 vssd1 vccd1 vccd1 _20194_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14160__A _22870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22904_ _22951_/CLK _22904_/D vssd1 vssd1 vccd1 vccd1 _22904_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22835_ _22929_/CLK _22847_/Q vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__19355__A2 _18718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13504__A _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12978__A2 _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22766_ _22799_/CLK _22766_/D vssd1 vssd1 vccd1 vccd1 _22766_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21717_ _21640_/C _21640_/D _21716_/Y vssd1 vssd1 vccd1 vccd1 _21717_/Y sky130_fd_sc_hd__a21oi_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22697_ _22701_/CLK _22697_/D vssd1 vssd1 vccd1 vccd1 _22697_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13927__A1 _13814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12450_ _12596_/A vssd1 vssd1 vccd1 vccd1 _12450_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_40_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21648_ _21618_/Y _21624_/Y _21662_/B _21647_/Y vssd1 vssd1 vccd1 vccd1 _21648_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_178_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20337__A _20337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11401_ _11477_/B _11477_/C _11477_/A vssd1 vssd1 vccd1 vccd1 _11401_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_166_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18866__A1 _17421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ _12606_/A _12607_/A _12574_/A vssd1 vssd1 vccd1 vccd1 _12383_/B sky130_fd_sc_hd__a21oi_1
XFILLER_181_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21579_ _21579_/A _21580_/A vssd1 vssd1 vccd1 vccd1 _21582_/A sky130_fd_sc_hd__nand2_1
XFILLER_193_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20673__A1 _15617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ _14122_/A _14057_/A _14119_/Y vssd1 vssd1 vccd1 vccd1 _14120_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__12781__C _16160_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11332_ _11709_/B _18875_/D _11372_/A _12062_/A vssd1 vssd1 vccd1 vccd1 _11333_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14051_ _14103_/B _14051_/B vssd1 vssd1 vccd1 vccd1 _14178_/B sky130_fd_sc_hd__or2_2
XFILLER_137_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13002_ _13002_/A _13002_/B _13002_/C vssd1 vssd1 vccd1 vccd1 _13003_/C sky130_fd_sc_hd__nand3_1
XFILLER_180_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21168__A _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20976__A2 _20975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17810_ _19844_/B _20972_/A _17895_/A _17811_/D vssd1 vssd1 vccd1 vccd1 _17812_/A
+ sky130_fd_sc_hd__a22o_1
X_18790_ _18432_/A _18603_/Y _18596_/B _18604_/Y vssd1 vssd1 vccd1 vccd1 _18970_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12115__B1 _12114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17741_ _17816_/B _17929_/A _17826_/A _17743_/D vssd1 vssd1 vccd1 vccd1 _17755_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_130_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14953_ _14953_/A vssd1 vssd1 vccd1 vccd1 _15064_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13904_ _22869_/Q vssd1 vssd1 vccd1 vccd1 _13904_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14220__D _14220_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17672_ _17672_/A vssd1 vssd1 vccd1 vccd1 _19334_/B sky130_fd_sc_hd__clkbuf_2
X_14884_ _14884_/A _14884_/B _14884_/C vssd1 vssd1 vccd1 vccd1 _14884_/X sky130_fd_sc_hd__and3_1
XFILLER_130_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19411_ _19422_/A vssd1 vssd1 vccd1 vccd1 _19411_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16623_ _16624_/A _16624_/B _16603_/Y _16622_/Y vssd1 vssd1 vccd1 vccd1 _16625_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_29_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13835_ _13736_/B _13833_/X _13989_/A _14112_/A vssd1 vssd1 vccd1 vccd1 _13877_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22900__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19342_ _19342_/A _19342_/B _19342_/C vssd1 vssd1 vccd1 vccd1 _19530_/C sky130_fd_sc_hd__nand3_2
X_16554_ _16554_/A _17530_/A _16554_/C vssd1 vssd1 vccd1 vccd1 _16557_/A sky130_fd_sc_hd__nand3_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17357__A1 _17226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ _13766_/A _13766_/B vssd1 vssd1 vccd1 vccd1 _14110_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11860__C _11860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17357__B2 _17215_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19897__A3 _18890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15505_ _12930_/A _15309_/B _17427_/A _15504_/X _12111_/X vssd1 vssd1 vccd1 vccd1
+ _15505_/X sky130_fd_sc_hd__o32a_1
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19273_ _19122_/Y _19123_/Y _19269_/Y vssd1 vssd1 vccd1 vccd1 _19299_/C sky130_fd_sc_hd__a21o_1
X_12717_ _15325_/A _15326_/A _22821_/Q _12579_/C _16256_/C vssd1 vssd1 vccd1 vccd1
+ _12718_/A sky130_fd_sc_hd__o2111ai_1
X_16485_ _14429_/A _16241_/C _16484_/X _11714_/A vssd1 vssd1 vccd1 vccd1 _17140_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11641__A2 _11606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_644 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13697_ _15005_/B vssd1 vssd1 vccd1 vccd1 _15114_/C sky130_fd_sc_hd__buf_2
X_18224_ _18226_/C _18275_/A _12221_/A _18223_/Y vssd1 vssd1 vccd1 vccd1 _18224_/Y
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_15_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18643__C _18933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15436_ _22961_/Q _22962_/Q vssd1 vssd1 vccd1 vccd1 _15486_/A sky130_fd_sc_hd__nor2_1
XFILLER_15_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17109__A1 _12827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12648_ _12745_/A _12745_/C _12745_/B vssd1 vssd1 vccd1 vccd1 _12651_/A sky130_fd_sc_hd__a21boi_1
XFILLER_175_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18155_ _18125_/X _18130_/Y _18154_/X vssd1 vssd1 vccd1 vccd1 _18155_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14591__A1 _13737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16317__C1 _20471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15367_ _15368_/A _15382_/B _15358_/X _15378_/A vssd1 vssd1 vccd1 vccd1 _15367_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_102_1114 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12579_ _15306_/C _15776_/D _12579_/C vssd1 vssd1 vccd1 vccd1 _12579_/X sky130_fd_sc_hd__and3_2
X_17106_ _16982_/A _17105_/Y _17188_/B vssd1 vssd1 vccd1 vccd1 _17177_/A sky130_fd_sc_hd__o21a_1
XFILLER_156_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14318_ input23/X _22586_/B vssd1 vssd1 vccd1 vccd1 _22442_/B sky130_fd_sc_hd__and2_1
X_18086_ _18079_/A _18079_/B _18084_/X _18080_/A vssd1 vssd1 vccd1 vccd1 _18087_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_144_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15298_ _12772_/A _12774_/A _14430_/A _15808_/A _18093_/D vssd1 vssd1 vccd1 vccd1
+ _15298_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_171_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17037_ _16873_/C _16858_/A _16856_/Y vssd1 vssd1 vccd1 vccd1 _17038_/C sky130_fd_sc_hd__a21o_1
XANTENNA__14343__A1 _13799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15540__B1 _18258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14343__B2 _13055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14249_ _14153_/A _14285_/C _14248_/B _14248_/A vssd1 vssd1 vccd1 vccd1 _14250_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_172_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19771__A _19771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _18493_/A _18875_/Y _18880_/B _18881_/X vssd1 vssd1 vccd1 vccd1 _19002_/B
+ sky130_fd_sc_hd__a2bb2oi_2
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_880 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17939_ _17939_/A _17991_/C vssd1 vssd1 vccd1 vccd1 _17940_/B sky130_fd_sc_hd__xor2_1
XANTENNA__19490__B _19490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater134 _22690_/CLK vssd1 vssd1 vccd1 vccd1 _22693_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater145 _22802_/CLK vssd1 vssd1 vccd1 vccd1 _22803_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater156 _22744_/CLK vssd1 vssd1 vccd1 vccd1 _22746_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15804__A _19012_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater167 _22735_/CLK vssd1 vssd1 vccd1 vccd1 _22800_/CLK sky130_fd_sc_hd__clkbuf_1
X_20950_ _20950_/A _20992_/A _20952_/A vssd1 vssd1 vccd1 vccd1 _20990_/A sky130_fd_sc_hd__nand3_1
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19609_ _19607_/A _19607_/B _19591_/Y _19594_/Y _19598_/Y vssd1 vssd1 vccd1 vccd1
+ _19610_/C sky130_fd_sc_hd__o221ai_1
XFILLER_4_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20881_ _20813_/X _20810_/A _20810_/B vssd1 vssd1 vccd1 vccd1 _20882_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__11880__A2 _11879_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15071__A2 _15154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22620_ _22620_/A vssd1 vssd1 vccd1 vccd1 _22798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22551_ _22551_/A vssd1 vssd1 vccd1 vccd1 _22767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_666 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21502_ _21485_/X _21492_/Y _21508_/B vssd1 vssd1 vccd1 vccd1 _21658_/A sky130_fd_sc_hd__o21ai_2
XFILLER_167_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22482_ _22737_/Q input43/X _22486_/S vssd1 vssd1 vccd1 vccd1 _22483_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16354__B _16617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11779__A _18107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21433_ _21433_/A _22674_/Q vssd1 vssd1 vccd1 vccd1 _21433_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11396__A1 _18259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21364_ _21367_/A _21367_/B _21448_/B vssd1 vssd1 vccd1 vccd1 _21365_/B sky130_fd_sc_hd__nand3_2
XFILLER_135_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20315_ _20191_/A _20314_/Y _20189_/Y _20192_/A vssd1 vssd1 vccd1 vccd1 _20315_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14305__D _14305_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21295_ _21295_/A _21295_/B vssd1 vssd1 vccd1 vccd1 _21296_/A sky130_fd_sc_hd__or2_1
XFILLER_190_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20246_ _20685_/A _12735_/X _20242_/X _20244_/X _20245_/X vssd1 vssd1 vccd1 vccd1
+ _20246_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_107_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20177_ _20177_/A vssd1 vssd1 vccd1 vccd1 _20178_/A sky130_fd_sc_hd__buf_2
XFILLER_190_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22923__CLK _22948_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15714__A _15714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _12003_/C vssd1 vssd1 vccd1 vccd1 _15714_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11961__B _12220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ _18445_/C vssd1 vssd1 vccd1 vccd1 _19202_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__11871__A2 _18984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13620_ _13566_/X _13599_/Y _13605_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22818_ _22850_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 _22818_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17339__A1 _17341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18536__B1 _15559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13551_ _13551_/A _13551_/B _13551_/C vssd1 vssd1 vccd1 vccd1 _13677_/B sky130_fd_sc_hd__nand3_2
X_22749_ _22749_/CLK _22749_/D vssd1 vssd1 vccd1 vccd1 _22749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12820__A1 _16778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ _12500_/X _12501_/X _12543_/A _20486_/C _12479_/B vssd1 vssd1 vccd1 vccd1
+ _12503_/B sky130_fd_sc_hd__o2111ai_1
X_16270_ _16258_/Y _16261_/Y _16269_/X vssd1 vssd1 vccd1 vccd1 _16272_/B sky130_fd_sc_hd__a21o_1
XFILLER_40_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13482_ _13484_/A _13484_/B _13484_/C vssd1 vssd1 vccd1 vccd1 _13485_/A sky130_fd_sc_hd__a21o_1
XFILLER_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15221_ _15224_/A _15224_/B _15224_/C _15224_/D vssd1 vssd1 vccd1 vccd1 _15242_/A
+ sky130_fd_sc_hd__nor4_4
X_12433_ _12403_/A _15631_/B _12413_/X _16318_/A vssd1 vssd1 vccd1 vccd1 _16778_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15152_ _15152_/A _15152_/B _15152_/C _15186_/D vssd1 vssd1 vccd1 vccd1 _15163_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_126_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ _12335_/A _12403_/D _12363_/Y _12378_/A vssd1 vssd1 vccd1 vccd1 _12404_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15117__A3 _15006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ _14103_/A _14103_/B _14103_/C vssd1 vssd1 vccd1 vccd1 _14104_/B sky130_fd_sc_hd__nand3_1
XFILLER_154_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11315_ _11325_/B _11315_/B _11404_/A vssd1 vssd1 vccd1 vccd1 _11316_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13128__A2 _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14325__A1 _11395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19960_ _20001_/A _19960_/B vssd1 vssd1 vccd1 vccd1 _19962_/C sky130_fd_sc_hd__nand2_1
XFILLER_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14325__B2 _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15083_ _15149_/A _14948_/C _15015_/A _15015_/C _15080_/Y vssd1 vssd1 vccd1 vccd1
+ _15083_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_107_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12295_ _22820_/Q vssd1 vssd1 vccd1 vccd1 _12415_/A sky130_fd_sc_hd__inv_2
XFILLER_181_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18911_ _18920_/B _18912_/A _18912_/B vssd1 vssd1 vccd1 vccd1 _18911_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16711__C _16711_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14034_ _14034_/A _14034_/B vssd1 vssd1 vccd1 vccd1 _14035_/B sky130_fd_sc_hd__nand2_1
X_19891_ _19891_/A _19891_/B _19976_/A _19891_/D vssd1 vssd1 vccd1 vccd1 _19891_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15608__B _22700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12887__B2 _20870_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18472__C1 _18387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18842_ _18259_/A _18678_/D _22798_/Q _18698_/B vssd1 vssd1 vccd1 vccd1 _18843_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_132_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18773_ _18773_/A _18773_/B _18774_/C _18774_/D vssd1 vssd1 vccd1 vccd1 _18773_/Y
+ sky130_fd_sc_hd__nand4_1
X_15985_ _15780_/B _15901_/Y _15900_/Y vssd1 vssd1 vccd1 vccd1 _16006_/A sky130_fd_sc_hd__o21ai_1
X_17724_ _17722_/Y _17723_/Y _17716_/A vssd1 vssd1 vccd1 vccd1 _17795_/B sky130_fd_sc_hd__o21bai_2
XANTENNA__15624__A _15624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14936_ _15050_/A _14861_/C _15050_/C _15114_/B _14934_/A vssd1 vssd1 vccd1 vccd1
+ _14936_/X sky130_fd_sc_hd__a32o_1
XFILLER_94_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17655_ _17739_/A _19768_/C _17645_/Y _17648_/Y vssd1 vssd1 vccd1 vccd1 _17655_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18357__D _19318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14867_ _14576_/X _14997_/A _14862_/Y _14866_/Y vssd1 vssd1 vccd1 vccd1 _14880_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_169_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19319__A2 _18135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1096 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16606_ _16606_/A _16606_/B _16606_/C vssd1 vssd1 vccd1 vccd1 _16606_/X sky130_fd_sc_hd__and3_1
X_13818_ _22868_/Q vssd1 vssd1 vccd1 vccd1 _14184_/C sky130_fd_sc_hd__clkbuf_4
X_17586_ _17579_/Y _17583_/Y _17585_/Y vssd1 vssd1 vccd1 vccd1 _17586_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15062__C _15114_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14798_ _14885_/B _14805_/C _14805_/D vssd1 vssd1 vccd1 vccd1 _14802_/A sky130_fd_sc_hd__nand3_1
XFILLER_32_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_763 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16537_ _16521_/Y _16529_/X _16531_/Y _16536_/Y vssd1 vssd1 vccd1 vccd1 _16624_/A
+ sky130_fd_sc_hd__o211ai_4
X_19325_ _18980_/C _19315_/X _19321_/Y _19324_/X vssd1 vssd1 vccd1 vccd1 _19326_/A
+ sky130_fd_sc_hd__o22ai_4
X_13749_ _13737_/X _13746_/X _13748_/X vssd1 vssd1 vccd1 vccd1 _14489_/B sky130_fd_sc_hd__a21oi_4
XFILLER_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15997__C _15997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19256_ _19116_/B _19117_/X _19116_/A _19253_/Y _19255_/Y vssd1 vssd1 vccd1 vccd1
+ _19296_/A sky130_fd_sc_hd__o2111ai_4
X_16468_ _16842_/A _16842_/B _16842_/C vssd1 vssd1 vccd1 vccd1 _16535_/A sky130_fd_sc_hd__a21oi_2
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17750__B2 _17981_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18207_ _18207_/A _18309_/A vssd1 vssd1 vccd1 vccd1 _18216_/B sky130_fd_sc_hd__nand2_2
X_15419_ _16058_/C _17131_/B _17108_/B _19154_/C vssd1 vssd1 vccd1 vccd1 _15419_/Y
+ sky130_fd_sc_hd__nand4_1
X_19187_ _19185_/B _19187_/B _19187_/C vssd1 vssd1 vccd1 vccd1 _19240_/B sky130_fd_sc_hd__nand3b_2
X_16399_ _16431_/C _16429_/A _16398_/X vssd1 vssd1 vccd1 vccd1 _16433_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12575__B1 _12988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18138_ _18140_/A _18338_/C _18140_/C vssd1 vssd1 vccd1 vccd1 _18340_/A sky130_fd_sc_hd__nand3_1
XFILLER_145_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18069_ _18066_/X _18082_/C _18069_/C _18069_/D vssd1 vssd1 vccd1 vccd1 _18075_/B
+ sky130_fd_sc_hd__nand4b_1
XFILLER_172_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20100_ _16267_/X _16266_/X _12988_/B _16268_/X vssd1 vssd1 vccd1 vccd1 _20110_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_132_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21080_ _21021_/A _21021_/B _21054_/B _21055_/B _21055_/A vssd1 vssd1 vccd1 vccd1
+ _21092_/A sky130_fd_sc_hd__a32oi_1
XANTENNA__22946__CLK _22948_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20031_ _20032_/B _20032_/C _22926_/Q vssd1 vssd1 vccd1 vccd1 _20058_/C sky130_fd_sc_hd__o21ai_1
XFILLER_98_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13319__A _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11550__A1 _11401_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19651__D _19945_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15534__A _22961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21982_ _22036_/A _22064_/A _22036_/B _22036_/C vssd1 vssd1 vccd1 vccd1 _21983_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20933_ _20933_/A _20933_/B vssd1 vssd1 vccd1 vccd1 _20933_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_148_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20864_ _20866_/B _20864_/B vssd1 vssd1 vccd1 vccd1 _20864_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22367__A _22368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_791 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22603_ _22603_/A vssd1 vssd1 vccd1 vccd1 _22790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16365__A _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20795_ _20792_/C _17313_/B _20577_/B _20793_/Y _20791_/Y vssd1 vssd1 vccd1 vccd1
+ _20797_/C sky130_fd_sc_hd__a32o_1
XFILLER_167_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22534_ _13896_/A input65/X _22536_/S vssd1 vssd1 vccd1 vccd1 _22535_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15700__C _15700_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17741__A1 _17816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16544__A2 _17391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_bq_clk_i clkbuf_4_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _22943_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14555__A1 _14843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22465_ _22465_/A vssd1 vssd1 vccd1 vccd1 _22729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_991 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21416_ _21416_/A vssd1 vssd1 vccd1 vccd1 _21417_/C sky130_fd_sc_hd__inv_2
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22396_ _16322_/B input37/X _22402_/S vssd1 vssd1 vccd1 vccd1 _22397_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21347_ _21346_/X _21198_/Y _21204_/Y _21238_/B _21237_/Y vssd1 vssd1 vccd1 vccd1
+ _21387_/B sky130_fd_sc_hd__a32oi_4
XFILLER_151_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11956__B _18093_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _12245_/A _12245_/B _12245_/C _18238_/A _18238_/B vssd1 vssd1 vccd1 vccd1
+ _12087_/B sky130_fd_sc_hd__a32oi_1
XFILLER_1_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21278_ _21278_/A _21278_/B _21278_/C vssd1 vssd1 vccd1 vccd1 _21423_/A sky130_fd_sc_hd__nand3_4
XFILLER_104_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19797__A2 _19795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20229_ _20206_/Y _20446_/B _20211_/Y _20236_/B _20236_/A vssd1 vssd1 vccd1 vccd1
+ _20229_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_104_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17643__B _18830_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17009__B1 _17006_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16480__A1 _15504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14086__A3 _14868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15444__A _15804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15770_ _15773_/B vssd1 vssd1 vccd1 vccd1 _16403_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12982_ _12982_/A _12982_/B vssd1 vssd1 vccd1 vccd1 _12989_/C sky130_fd_sc_hd__nand2_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A wb_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14721_ _14892_/A _14721_/B _15005_/B _14808_/D vssd1 vssd1 vccd1 vccd1 _14727_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _12035_/A _12035_/B _12036_/A _11931_/X _11932_/Y vssd1 vssd1 vccd1 vccd1
+ _11933_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_40_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21991__B1_N _21990_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18755__A _18765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _17440_/A vssd1 vssd1 vccd1 vccd1 _17880_/A sky130_fd_sc_hd__buf_2
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14652_ _14638_/Y _14650_/X _14651_/Y vssd1 vssd1 vccd1 vccd1 _14656_/B sky130_fd_sc_hd__o21ai_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _18875_/D vssd1 vssd1 vccd1 vccd1 _16712_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13046__A1 _12754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13603_ _13526_/A _13526_/B _13527_/Y _13530_/X _13524_/X vssd1 vssd1 vccd1 vccd1
+ _13603_/Y sky130_fd_sc_hd__o221ai_4
X_17371_ _17371_/A _17371_/B vssd1 vssd1 vccd1 vccd1 _17372_/B sky130_fd_sc_hd__nor2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14583_ _22763_/Q _14583_/B _14583_/C _14583_/D vssd1 vssd1 vccd1 vccd1 _14583_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_14_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16275__A _16275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11795_ _11789_/X _11791_/X _11976_/A vssd1 vssd1 vccd1 vccd1 _11797_/A sky130_fd_sc_hd__o21ai_1
XFILLER_159_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19110_ _19112_/A _19112_/B vssd1 vssd1 vccd1 vccd1 _19116_/B sky130_fd_sc_hd__nand2_2
XANTENNA__22819__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16322_ _16322_/A _16322_/B _22700_/Q vssd1 vssd1 vccd1 vccd1 _16323_/D sky130_fd_sc_hd__nor3_2
X_13534_ _13461_/Y _13463_/Y _13465_/Y vssd1 vssd1 vccd1 vccd1 _13534_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19041_ _18795_/A _17400_/A _17393_/X _12116_/X vssd1 vssd1 vccd1 vccd1 _19045_/A
+ sky130_fd_sc_hd__o22ai_1
X_16253_ _16253_/A _16253_/B vssd1 vssd1 vccd1 vccd1 _16253_/Y sky130_fd_sc_hd__nand2_1
X_13465_ _13465_/A _13465_/B _21362_/B _13591_/A vssd1 vssd1 vccd1 vccd1 _13465_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_186_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12308__A _22703_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15204_ _15205_/A _15205_/B _15205_/C vssd1 vssd1 vccd1 vccd1 _15206_/A sky130_fd_sc_hd__a21oi_1
X_12416_ _20130_/A _12904_/A vssd1 vssd1 vccd1 vccd1 _12921_/A sky130_fd_sc_hd__nand2_4
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16184_ _16141_/X _16140_/Y _16173_/Y vssd1 vssd1 vccd1 vccd1 _16184_/Y sky130_fd_sc_hd__o21ai_1
X_13396_ _13396_/A _13396_/B _13396_/C vssd1 vssd1 vccd1 vccd1 _13396_/X sky130_fd_sc_hd__and3_1
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15135_ _15135_/A _15135_/B vssd1 vssd1 vccd1 vccd1 _15135_/X sky130_fd_sc_hd__or2_1
XANTENNA__15619__A _16715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ _16267_/A _16266_/A _16268_/A vssd1 vssd1 vccd1 vccd1 _15314_/A sky130_fd_sc_hd__a21oi_2
XFILLER_5_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14849__A2 _14845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19943_ _19842_/D _19461_/B _19461_/C _19945_/A _19945_/D vssd1 vssd1 vccd1 vccd1
+ _19946_/A sky130_fd_sc_hd__a32o_1
X_15066_ _15062_/Y _15059_/Y _15058_/X vssd1 vssd1 vccd1 vccd1 _15066_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ _12303_/A vssd1 vssd1 vccd1 vccd1 _15363_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_141_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14017_ _13848_/A _13854_/A _13862_/A vssd1 vssd1 vccd1 vccd1 _14017_/X sky130_fd_sc_hd__a21o_1
X_19874_ _19872_/A _19872_/B _19921_/A _19921_/B vssd1 vssd1 vccd1 vccd1 _19919_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18825_ _18825_/A _18825_/B vssd1 vssd1 vccd1 vccd1 _19080_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18460__A2 _17400_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_658 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18756_ _18763_/A _18754_/X _18764_/B vssd1 vssd1 vccd1 vccd1 _18762_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13285__A1 _13475_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15968_ _15898_/Y _15913_/Y _15915_/Y _15916_/Y vssd1 vssd1 vccd1 vccd1 _15971_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17707_ _17781_/C vssd1 vssd1 vccd1 vccd1 _17708_/B sky130_fd_sc_hd__inv_2
X_14919_ _14919_/A _14919_/B _14919_/C vssd1 vssd1 vccd1 vccd1 _14921_/A sky130_fd_sc_hd__nand3_1
XFILLER_82_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18687_ _18706_/B _18876_/B vssd1 vssd1 vccd1 vccd1 _19160_/A sky130_fd_sc_hd__nand2_4
X_15899_ _16308_/C _15899_/B _20134_/B vssd1 vssd1 vccd1 vccd1 _16006_/B sky130_fd_sc_hd__and3_1
XANTENNA__20555__B1 _20548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18665__A _18665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17638_ _12234_/X _12237_/X _17440_/A vssd1 vssd1 vccd1 vccd1 _17638_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16774__A2 _12571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17569_ _17574_/A vssd1 vssd1 vccd1 vccd1 _17626_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19199__C _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11599__A1 _15932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19308_ _18843_/A _18843_/B _11511_/X vssd1 vssd1 vccd1 vccd1 _19308_/X sky130_fd_sc_hd__a21o_2
X_20580_ _20577_/Y _20578_/X _20579_/X vssd1 vssd1 vccd1 vccd1 _20586_/A sky130_fd_sc_hd__o21ai_1
XFILLER_182_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19496__A _19496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19239_ _19035_/X _19037_/X _19010_/X vssd1 vssd1 vccd1 vccd1 _19239_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16913__A _17110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21807__B1 _21806_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22250_ _22250_/A _22683_/Q _22250_/C vssd1 vssd1 vccd1 vccd1 _22251_/B sky130_fd_sc_hd__nand3_1
XFILLER_191_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21201_ _22229_/A _21195_/C _22229_/C _13309_/B _21851_/C vssd1 vssd1 vccd1 vccd1
+ _21201_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_145_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22181_ _22182_/A _22221_/C _22182_/C vssd1 vssd1 vccd1 vccd1 _22181_/Y sky130_fd_sc_hd__nand3_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14433__A _22965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21132_ _21150_/A _21150_/B vssd1 vssd1 vccd1 vccd1 _21143_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17239__B1 _17238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13049__A _22843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21063_ _21097_/A _21061_/Y _21095_/B _21095_/A vssd1 vssd1 vccd1 vccd1 _21068_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_132_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11523__A1 _11285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20014_ _18029_/D _19901_/B _20012_/X _20013_/X vssd1 vssd1 vccd1 vccd1 _20016_/A
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__18987__B1 _18986_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__B2 _11295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20243__C1 _16257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input4_A wb_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_978 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13276__A1 _21853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21965_ _21964_/X _21958_/X _21960_/Y vssd1 vssd1 vccd1 vccd1 _21965_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _20920_/A _20916_/B _20916_/C vssd1 vssd1 vccd1 vccd1 _20923_/B sky130_fd_sc_hd__nand3b_2
XFILLER_42_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21896_ _21896_/A _21933_/B vssd1 vssd1 vccd1 vccd1 _21902_/B sky130_fd_sc_hd__nand2_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_508 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20847_ _20793_/A _20792_/A _20792_/B _20936_/B _20793_/D vssd1 vssd1 vccd1 vccd1
+ _20848_/B sky130_fd_sc_hd__a32o_1
XFILLER_168_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20849__A1 _13022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11580_ _11587_/A _18339_/C _11587_/C vssd1 vssd1 vccd1 vccd1 _11789_/A sky130_fd_sc_hd__nand3_1
X_20778_ _20778_/A _20778_/B vssd1 vssd1 vccd1 vccd1 _20812_/B sky130_fd_sc_hd__nand2_1
XFILLER_168_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22517_ _14220_/D input35/X _22525_/S vssd1 vssd1 vccd1 vccd1 _22518_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15725__B1 _15991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13250_ _22848_/Q vssd1 vssd1 vccd1 vccd1 _21367_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22448_ _22448_/A vssd1 vssd1 vccd1 vccd1 _22721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12201_ _12212_/B _22662_/B vssd1 vssd1 vccd1 vccd1 _12202_/B sky130_fd_sc_hd__nand2_4
XFILLER_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _13221_/A _13181_/B _13181_/C vssd1 vssd1 vccd1 vccd1 _13475_/C sky130_fd_sc_hd__nand3b_2
XFILLER_164_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22379_ _22379_/A vssd1 vssd1 vccd1 vccd1 _22691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16261__C _17280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12132_ _12126_/X _12128_/X _12131_/Y vssd1 vssd1 vccd1 vccd1 _12134_/A sky130_fd_sc_hd__o21ai_1
XFILLER_151_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16940_ _16940_/A vssd1 vssd1 vccd1 vccd1 _16940_/X sky130_fd_sc_hd__clkbuf_4
X_12063_ _12116_/A vssd1 vssd1 vccd1 vccd1 _12064_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16871_ _16637_/A _16706_/A _16705_/Y vssd1 vssd1 vccd1 vccd1 _16874_/A sky130_fd_sc_hd__a21oi_1
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16453__A1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18610_ _11877_/Y _11879_/Y _15530_/A _15531_/A vssd1 vssd1 vccd1 vccd1 _18610_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _19317_/D vssd1 vssd1 vccd1 vccd1 _19614_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ _15522_/X _15521_/X _15523_/X _18718_/X vssd1 vssd1 vccd1 vccd1 _19590_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_18_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18541_ _18664_/B _18533_/Y _18534_/X vssd1 vssd1 vccd1 vccd1 _18543_/B sky130_fd_sc_hd__a21o_1
X_15753_ _15733_/A _15733_/B _15733_/C _15727_/B _15727_/A vssd1 vssd1 vccd1 vccd1
+ _15753_/Y sky130_fd_sc_hd__a311oi_4
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _12749_/B _12749_/A _13007_/C _13007_/B vssd1 vssd1 vccd1 vccd1 _12966_/C
+ sky130_fd_sc_hd__o211ai_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19942__A2 _19322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11916_ _18459_/C vssd1 vssd1 vccd1 vccd1 _18830_/A sky130_fd_sc_hd__buf_2
X_14704_ _14861_/A _14868_/B _14191_/C _14706_/B vssd1 vssd1 vccd1 vccd1 _14815_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15684_ _15682_/A _15512_/Y _15514_/X vssd1 vssd1 vccd1 vccd1 _15684_/Y sky130_fd_sc_hd__a21oi_1
X_18472_ _12064_/A _18372_/X _17442_/X _18105_/Y _18387_/B vssd1 vssd1 vccd1 vccd1
+ _18472_/X sky130_fd_sc_hd__o311a_1
XANTENNA__13019__A1 _15577_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12896_ _12896_/A vssd1 vssd1 vccd1 vccd1 _13007_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16717__B _20781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _17423_/A vssd1 vssd1 vccd1 vccd1 _17423_/X sky130_fd_sc_hd__buf_2
X_14635_ _14635_/A _14635_/B _14635_/C vssd1 vssd1 vccd1 vccd1 _14636_/D sky130_fd_sc_hd__nand3_2
X_11847_ _16078_/C vssd1 vssd1 vccd1 vccd1 _15978_/C sky130_fd_sc_hd__buf_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_878 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19155__B1 _19154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _17210_/B _17230_/Y _17352_/X vssd1 vssd1 vccd1 vccd1 _17354_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14566_ _14566_/A vssd1 vssd1 vccd1 vccd1 _15058_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11778_/A _11778_/B vssd1 vssd1 vccd1 vccd1 _11779_/C sky130_fd_sc_hd__nand2_4
XFILLER_174_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16305_ _15638_/X _16552_/A _15711_/A _16296_/Y _20593_/A vssd1 vssd1 vccd1 vccd1
+ _16305_/Y sky130_fd_sc_hd__o2111ai_4
X_13517_ _13517_/A _21480_/B _13517_/C vssd1 vssd1 vccd1 vccd1 _13517_/X sky130_fd_sc_hd__and3_1
X_17285_ _17288_/A _17288_/B _17285_/C _17285_/D vssd1 vssd1 vccd1 vccd1 _17285_/Y
+ sky130_fd_sc_hd__nand4_4
XANTENNA__15716__B1 _15711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14497_ _14497_/A _14497_/B vssd1 vssd1 vccd1 vccd1 _14497_/Y sky130_fd_sc_hd__nand2_2
XFILLER_9_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16236_ _16236_/A vssd1 vssd1 vccd1 vccd1 _16474_/A sky130_fd_sc_hd__buf_2
X_19024_ _19350_/A _17434_/A _19014_/X _19015_/Y _19017_/Y vssd1 vssd1 vccd1 vccd1
+ _19024_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13448_ _13050_/X _13343_/A _13446_/X _13447_/X vssd1 vssd1 vccd1 vccd1 _13455_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_162_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20255__A _20255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16167_ _16162_/X _16165_/Y _16166_/Y vssd1 vssd1 vccd1 vccd1 _16168_/B sky130_fd_sc_hd__o21a_1
X_13379_ _13502_/D vssd1 vssd1 vccd1 vccd1 _21498_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_6_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15118_ _15118_/A _15215_/A _15118_/C vssd1 vssd1 vccd1 vccd1 _15120_/B sky130_fd_sc_hd__and3_1
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16098_ _16098_/A vssd1 vssd1 vccd1 vccd1 _16098_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_141_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19926_ _19926_/A vssd1 vssd1 vccd1 vccd1 _19928_/A sky130_fd_sc_hd__inv_2
X_15049_ _15114_/B vssd1 vssd1 vccd1 vccd1 _15215_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__19482__C _20012_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19857_ _19856_/B _19913_/A _19856_/A vssd1 vssd1 vccd1 vccd1 _19860_/C sky130_fd_sc_hd__o21a_1
XFILLER_122_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18808_ _18616_/B _18618_/B _18611_/Y _18610_/X vssd1 vssd1 vccd1 vccd1 _18824_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_110_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14455__B1 _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19788_ _19788_/A _19788_/B _19837_/B vssd1 vssd1 vccd1 vccd1 _19796_/B sky130_fd_sc_hd__nand3_2
XANTENNA__12501__A _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22517__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18739_ _18826_/A _18827_/A _18664_/X _18666_/X vssd1 vssd1 vccd1 vccd1 _18741_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_3_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21750_ _21876_/A _21877_/A _21750_/C vssd1 vssd1 vccd1 vccd1 _21751_/B sky130_fd_sc_hd__nand3_1
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16747__A2 _16746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20701_ _20796_/B _20797_/A _20796_/A vssd1 vssd1 vccd1 vccd1 _20702_/D sky130_fd_sc_hd__a21o_1
XFILLER_196_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21681_ _21539_/A _21539_/B _21524_/A vssd1 vssd1 vccd1 vccd1 _21687_/C sky130_fd_sc_hd__o21ai_2
XFILLER_196_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20632_ _20501_/X _20623_/Y _20624_/X vssd1 vssd1 vccd1 vccd1 _20738_/A sky130_fd_sc_hd__a21oi_2
XFILLER_32_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14147__B _14147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17739__A _17739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20563_ _20563_/A _20563_/B vssd1 vssd1 vccd1 vccd1 _20564_/B sky130_fd_sc_hd__nand2_2
XFILLER_149_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22302_ _22302_/A _22302_/B vssd1 vssd1 vccd1 vccd1 _22302_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20494_ _12697_/A _16331_/A _20587_/A _20462_/A vssd1 vssd1 vccd1 vccd1 _20581_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_121_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21256__A1 _21683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22233_ _22233_/A _22233_/B vssd1 vssd1 vccd1 vccd1 _22271_/B sky130_fd_sc_hd__xor2_1
XFILLER_30_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22164_ _22164_/A vssd1 vssd1 vccd1 vccd1 _22164_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21115_ _21115_/A _21115_/B vssd1 vssd1 vccd1 vccd1 _21115_/Y sky130_fd_sc_hd__nand2_1
XFILLER_161_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22095_ _22290_/A _22290_/B vssd1 vssd1 vccd1 vccd1 _22937_/D sky130_fd_sc_hd__xor2_1
X_21046_ _21046_/A _21046_/B _21021_/B vssd1 vssd1 vccd1 vccd1 _21054_/A sky130_fd_sc_hd__or3b_1
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13507__A _21724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1078 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22664__CLK _22959_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21724__A _21724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _12896_/A _12750_/B vssd1 vssd1 vccd1 vccd1 _12751_/B sky130_fd_sc_hd__nand2_1
X_21948_ _21767_/X _21594_/Y _22045_/A _22045_/B _21952_/C vssd1 vssd1 vccd1 vccd1
+ _21948_/X sky130_fd_sc_hd__o221a_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11701_ _11819_/A vssd1 vssd1 vccd1 vccd1 _12111_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12681_ _12681_/A _12681_/B _20101_/C vssd1 vssd1 vccd1 vccd1 _12681_/X sky130_fd_sc_hd__and3_1
XFILLER_187_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21879_ _21383_/X _21970_/A _21742_/B _21939_/A _21972_/A vssd1 vssd1 vccd1 vccd1
+ _21879_/Y sky130_fd_sc_hd__o221ai_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _22715_/Q _14418_/X _14410_/X _22747_/Q _14419_/X vssd1 vssd1 vccd1 vccd1
+ _14420_/X sky130_fd_sc_hd__a221o_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14213__A3 _14765_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11644_/A _11645_/A _11645_/B _11553_/B _11552_/B vssd1 vssd1 vccd1 vccd1
+ _11698_/B sky130_fd_sc_hd__a32oi_2
XANTENNA__19688__A1 _19585_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14351_ _14351_/A vssd1 vssd1 vccd1 vccd1 _14351_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17649__A _20928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11563_ _11568_/B vssd1 vssd1 vccd1 vccd1 _11563_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__18360__A1 _17421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _13302_/A vssd1 vssd1 vccd1 vccd1 _21336_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_183_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17070_ _17070_/A _17070_/B vssd1 vssd1 vccd1 vccd1 _17071_/C sky130_fd_sc_hd__nand2_1
XFILLER_155_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14282_ _14282_/A _14282_/B vssd1 vssd1 vccd1 vccd1 _14282_/Y sky130_fd_sc_hd__nand2_1
XFILLER_183_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11494_ _11980_/A _11619_/B _18115_/D vssd1 vssd1 vccd1 vccd1 _11792_/A sky130_fd_sc_hd__a21o_1
XFILLER_171_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16021_ _15971_/A _15927_/Y _15970_/B _15970_/A vssd1 vssd1 vccd1 vccd1 _16021_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13233_ _13633_/B vssd1 vssd1 vccd1 vccd1 _21259_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164_ _13164_/A vssd1 vssd1 vccd1 vccd1 _13384_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__19583__B _19687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16674__A1 _17226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ _12116_/A _12111_/X _11935_/C _12114_/X _18203_/B vssd1 vssd1 vccd1 vccd1
+ _12115_/X sky130_fd_sc_hd__o32a_1
XANTENNA__17384__A _19496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17972_ _18007_/D _17972_/B vssd1 vssd1 vccd1 vccd1 _22964_/D sky130_fd_sc_hd__xor2_1
X_13095_ _13095_/A vssd1 vssd1 vccd1 vccd1 _13095_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19711_ _19720_/C vssd1 vssd1 vccd1 vccd1 _19864_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16923_ _16782_/X _16781_/Y _16792_/B _16787_/Y vssd1 vssd1 vccd1 vccd1 _16923_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
X_12046_ _12046_/A vssd1 vssd1 vccd1 vccd1 _12046_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21469__A_N _13112_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19642_ _19528_/A _19528_/B _19528_/C _19543_/Y vssd1 vssd1 vccd1 vccd1 _19642_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_38_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16854_ _16866_/A _16866_/B _16852_/Y _16853_/X vssd1 vssd1 vccd1 vccd1 _16860_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_133_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16977__A2 _15723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15805_ _12988_/A _17427_/A _15298_/Y vssd1 vssd1 vccd1 vccd1 _15805_/Y sky130_fd_sc_hd__o21ai_2
X_19573_ _19574_/A _19574_/B _19574_/C vssd1 vssd1 vccd1 vccd1 _19575_/A sky130_fd_sc_hd__a21oi_1
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16785_ _18282_/A vssd1 vssd1 vccd1 vccd1 _17636_/A sky130_fd_sc_hd__clkbuf_4
X_13997_ _13877_/B _14468_/A _13873_/A _13986_/Y _14889_/A vssd1 vssd1 vccd1 vccd1
+ _13998_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_81_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18524_ _18526_/A _18526_/B _18491_/A _18526_/D vssd1 vssd1 vccd1 vccd1 _18527_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15736_ _15859_/A _15859_/B vssd1 vssd1 vccd1 vccd1 _15860_/A sky130_fd_sc_hd__nand2_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12948_ _15991_/B vssd1 vssd1 vccd1 vccd1 _20390_/C sky130_fd_sc_hd__buf_2
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16447__B _20323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18455_ _12202_/A _12202_/B _18281_/Y vssd1 vssd1 vccd1 vccd1 _18455_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__15937__B1 _15935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15667_ _15667_/A _15673_/A vssd1 vssd1 vccd1 vccd1 _15678_/C sky130_fd_sc_hd__nand2_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _12876_/X _20870_/C _12878_/X _12776_/X vssd1 vssd1 vccd1 vccd1 _12879_/Y
+ sky130_fd_sc_hd__a211oi_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13152__A _22844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17406_ _17406_/A vssd1 vssd1 vccd1 vccd1 _18303_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17941__A4 _21081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14618_ _14618_/A vssd1 vssd1 vccd1 vccd1 _14942_/A sky130_fd_sc_hd__buf_2
XFILLER_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15598_ _15672_/A _15672_/B _15596_/Y _15597_/Y vssd1 vssd1 vccd1 vccd1 _15678_/A
+ sky130_fd_sc_hd__o2bb2ai_2
X_18386_ _18387_/A _18387_/B _18387_/C vssd1 vssd1 vccd1 vccd1 _18407_/A sky130_fd_sc_hd__a21oi_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17337_ _17337_/A vssd1 vssd1 vccd1 vccd1 _17337_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14549_ _14661_/C _14549_/B vssd1 vssd1 vccd1 vccd1 _14554_/B sky130_fd_sc_hd__xor2_4
XFILLER_159_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17268_ _17298_/B _17268_/B vssd1 vssd1 vccd1 vccd1 _17269_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16362__B1 _20793_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16901__A2 _16685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17338__A_N _17103_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19007_ _19179_/C _19007_/B vssd1 vssd1 vccd1 vccd1 _19007_/Y sky130_fd_sc_hd__nor2_1
X_16219_ _12500_/A _12501_/A _18192_/A _18193_/A vssd1 vssd1 vccd1 vccd1 _16236_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17199_ _17186_/X _17193_/Y _17197_/Y _17198_/X vssd1 vssd1 vccd1 vccd1 _17205_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16613__D _16613_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22687__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20432__B _20432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19909_ _19909_/A _19909_/B _19909_/C vssd1 vssd1 vccd1 vccd1 _19909_/X sky130_fd_sc_hd__or3_1
XANTENNA__19603__A1 _18131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__21247__C _21247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22920_ _22922_/CLK _22920_/D vssd1 vssd1 vccd1 vccd1 _22920_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14428__B1 _14351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22851_ _22929_/CLK _22863_/Q vssd1 vssd1 vccd1 vccd1 _22851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15640__A2 _15938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21802_ _21802_/A _21899_/A _21802_/C vssd1 vssd1 vccd1 vccd1 _21803_/C sky130_fd_sc_hd__nand3_1
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19014__A _19014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22782_ _22815_/CLK _22782_/D vssd1 vssd1 vccd1 vccd1 _22782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21733_ _21733_/A _22034_/A _22108_/C _22106_/A vssd1 vssd1 vccd1 vccd1 _21733_/X
+ sky130_fd_sc_hd__and4_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13062__A _22735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21664_ _21664_/A vssd1 vssd1 vccd1 vccd1 _21664_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18572__B _18572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20615_ _20606_/Y _20608_/Y _20609_/X vssd1 vssd1 vccd1 vccd1 _20615_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_178_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18342__A1 _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21595_ _21936_/A _21595_/B _21937_/A vssd1 vssd1 vccd1 vccd1 _21751_/A sky130_fd_sc_hd__nand3_1
XFILLER_193_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16353__B1 _16310_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20546_ _20658_/A _20658_/B _20544_/X _20545_/Y vssd1 vssd1 vccd1 vccd1 _20546_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_137_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18893__A2 _18856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13167__B1 _13166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14605__B _14953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14364__C1 _14363_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20477_ _20477_/A _20481_/C vssd1 vssd1 vccd1 vccd1 _20482_/A sky130_fd_sc_hd__nand2_2
XFILLER_193_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11310__A _22956_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22216_ _22216_/A _22216_/B vssd1 vssd1 vccd1 vccd1 _22216_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17448__A3 _19619_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22147_ _22156_/A _22156_/B _22212_/A _22089_/A vssd1 vssd1 vccd1 vccd1 _22150_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14667__B1 _14845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15436__B _22962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22078_ _22073_/Y _22074_/Y _22075_/X vssd1 vssd1 vccd1 vccd1 _22080_/A sky130_fd_sc_hd__o21ai_1
XFILLER_86_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13237__A _13423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18948__A3 _18626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13920_ _13920_/A _13920_/B _13920_/C vssd1 vssd1 vccd1 vccd1 _14021_/D sky130_fd_sc_hd__nand3_1
X_21029_ _21030_/B _21030_/C _21030_/A vssd1 vssd1 vccd1 vccd1 _21095_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__14419__B1 _14413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13851_ _13851_/A _13851_/B vssd1 vssd1 vccd1 vccd1 _13984_/A sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_3_4_0_bq_clk_i_A clkbuf_3_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15452__A _19322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ _12802_/A _12813_/A _12802_/C vssd1 vssd1 vccd1 vccd1 _12803_/A sky130_fd_sc_hd__nand3_1
XFILLER_142_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16570_ _16570_/A vssd1 vssd1 vccd1 vccd1 _16879_/A sky130_fd_sc_hd__buf_2
X_13782_ _14199_/A _15008_/C _13781_/A _14043_/A vssd1 vssd1 vccd1 vccd1 _13784_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15521_ _15521_/A vssd1 vssd1 vccd1 vccd1 _15521_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _12702_/A _12716_/A _12592_/B vssd1 vssd1 vccd1 vccd1 _12950_/B sky130_fd_sc_hd__o21ai_2
XFILLER_188_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15452_ _19322_/A _17280_/A _16772_/A _15997_/C vssd1 vssd1 vccd1 vccd1 _15452_/Y
+ sky130_fd_sc_hd__nand4_2
X_18240_ _18240_/A _18240_/B vssd1 vssd1 vccd1 vccd1 _18240_/Y sky130_fd_sc_hd__nor2_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _16160_/C _20723_/A _12757_/B vssd1 vssd1 vccd1 vccd1 _12665_/B sky130_fd_sc_hd__a21oi_1
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18482__B _18482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14403_ _22369_/D vssd1 vssd1 vccd1 vccd1 _14403_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11615_ _11615_/A _11995_/B vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__nand2_1
XFILLER_168_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17379__A _17379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15383_ _15664_/A _15665_/A _15665_/B _15665_/C vssd1 vssd1 vccd1 vccd1 _15384_/C
+ sky130_fd_sc_hd__nand4_1
X_18171_ _18365_/A _18995_/A _19504_/D _18125_/X _18980_/A vssd1 vssd1 vccd1 vccd1
+ _18310_/B sky130_fd_sc_hd__o2111ai_4
X_12595_ _12701_/A _12598_/A _12594_/Y vssd1 vssd1 vccd1 vccd1 _12595_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17122_ _17122_/A _17122_/B _17122_/C vssd1 vssd1 vccd1 vccd1 _17122_/Y sky130_fd_sc_hd__nand3_1
X_14334_ _14361_/A vssd1 vssd1 vccd1 vccd1 _14334_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11546_ _11644_/A _11645_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _11552_/A sky130_fd_sc_hd__nand3_1
XFILLER_184_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18884__A2 _19313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _17053_/A _17053_/B vssd1 vssd1 vccd1 vccd1 _17053_/Y sky130_fd_sc_hd__nand2_1
XFILLER_183_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14265_ _14265_/A _14265_/B vssd1 vssd1 vccd1 vccd1 _14267_/C sky130_fd_sc_hd__nand2_1
XFILLER_156_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11477_ _11477_/A _11477_/B _11477_/C vssd1 vssd1 vccd1 vccd1 _11893_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11708__A1 _11502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11708__B2 _11705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16004_ _16133_/B vssd1 vssd1 vccd1 vccd1 _16093_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18097__B1 _18849_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13216_ _13216_/A _13216_/B vssd1 vssd1 vccd1 vccd1 _13221_/B sky130_fd_sc_hd__nand2_1
XANTENNA__21629__A _21724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14196_ _14198_/C _14198_/D vssd1 vssd1 vccd1 vccd1 _14197_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13147_ _13147_/A _13147_/B vssd1 vssd1 vccd1 vccd1 _13513_/B sky130_fd_sc_hd__nand2_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _17785_/X _17954_/B _17857_/B _17857_/A vssd1 vssd1 vccd1 vccd1 _17955_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _13301_/A _13302_/A _21307_/C vssd1 vssd1 vccd1 vccd1 _13304_/A sky130_fd_sc_hd__o21ai_1
XFILLER_140_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16906_ _16906_/A _16906_/B _16906_/C vssd1 vssd1 vccd1 vccd1 _16906_/X sky130_fd_sc_hd__and3_1
X_12029_ _11930_/X _11933_/Y _12027_/Y _12028_/X vssd1 vssd1 vccd1 vccd1 _12029_/Y
+ sky130_fd_sc_hd__o211ai_2
X_17886_ _17886_/A _17886_/B _17886_/C vssd1 vssd1 vccd1 vccd1 _17888_/A sky130_fd_sc_hd__nand3_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20746__A3 _20734_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19625_ _19625_/A vssd1 vssd1 vccd1 vccd1 _19793_/A sky130_fd_sc_hd__buf_2
X_16837_ _16828_/A _16831_/B _16836_/X vssd1 vssd1 vccd1 vccd1 _16845_/C sky130_fd_sc_hd__a21o_1
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12986__A _20593_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11890__A _16157_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15622__A2 _16300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19556_ _19556_/A vssd1 vssd1 vccd1 vccd1 _19556_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21083__B _21083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16768_ _16768_/A _16768_/B _16768_/C vssd1 vssd1 vccd1 vccd1 _16972_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12436__A2 _16779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18507_ _18706_/B _18999_/A _18507_/C vssd1 vssd1 vccd1 vccd1 _18508_/B sky130_fd_sc_hd__nand3_1
XFILLER_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15719_ _11912_/A _15723_/A _15341_/X _12009_/X vssd1 vssd1 vccd1 vccd1 _15959_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_62_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19487_ _19342_/A _19342_/B _19342_/C _19340_/A vssd1 vssd1 vccd1 vccd1 _19488_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_80_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16699_ _16685_/A _16682_/Y _16698_/Y vssd1 vssd1 vccd1 vccd1 _16700_/B sky130_fd_sc_hd__o21a_1
XANTENNA__18673__A _19351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18438_ _12249_/A _18241_/B _18428_/Y _18427_/X vssd1 vssd1 vccd1 vccd1 _18438_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_178_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19488__B _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18369_ _18365_/Y _18366_/Y _18367_/Y _18368_/Y vssd1 vssd1 vccd1 vccd1 _18387_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_187_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20400_ _20397_/Y _20398_/Y _20399_/Y _20154_/B vssd1 vssd1 vccd1 vccd1 _20400_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_193_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_330 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16335__B1 _16354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21380_ _21230_/A _21230_/B _21230_/C vssd1 vssd1 vccd1 vccd1 _21380_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20331_ _20247_/Y _20326_/Y _20508_/A _20324_/Y _20129_/A vssd1 vssd1 vccd1 vccd1
+ _20447_/B sky130_fd_sc_hd__o2111a_1
XANTENNA__14346__C1 _14345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19824__A1 _19293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18627__A2 _15541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20262_ _20262_/A _20262_/B _20262_/C vssd1 vssd1 vccd1 vccd1 _20263_/A sky130_fd_sc_hd__nand3_4
XFILLER_143_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22001_ _21996_/Y _21999_/Y _22000_/X _21842_/X vssd1 vssd1 vccd1 vccd1 _22008_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20193_ _22931_/Q vssd1 vssd1 vccd1 vccd1 _20311_/A sky130_fd_sc_hd__inv_2
XANTENNA__12911__A3 _12680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16102__A3 _20452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18848__A _19194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13321__B1 _13126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17063__A1 _17226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22903_ _22951_/CLK _22903_/D vssd1 vssd1 vccd1 vccd1 _22903_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22834_ _22929_/CLK _22846_/Q vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12427__A2 _15363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11635__B1 _19043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22765_ _22765_/CLK _22765_/D vssd1 vssd1 vccd1 vccd1 _22765_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12832__C1 _20092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21716_ _21716_/A _21716_/B vssd1 vssd1 vccd1 vccd1 _21716_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22696_ _22696_/CLK _22696_/D vssd1 vssd1 vccd1 vccd1 _22696_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16574__B1 _22702_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21647_ _21485_/X _21649_/A _21645_/Y _21646_/Y vssd1 vssd1 vccd1 vccd1 _21647_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13927__A2 _13814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11400_ _11371_/X _11393_/Y _11399_/Y vssd1 vssd1 vccd1 vccd1 _11477_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__22852__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12380_ _22817_/Q vssd1 vssd1 vccd1 vccd1 _12574_/A sky130_fd_sc_hd__inv_2
XANTENNA__12060__B1 _11693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18866__A2 _17422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21578_ _21578_/A vssd1 vssd1 vccd1 vccd1 _21579_/A sky130_fd_sc_hd__buf_2
XFILLER_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11331_ _11331_/A vssd1 vssd1 vccd1 vccd1 _12062_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__20673__A2 _12827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20529_ _20529_/A vssd1 vssd1 vccd1 vccd1 _20568_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_153_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16831__A _16831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ _14054_/A _14055_/B _14049_/A _14165_/A vssd1 vssd1 vccd1 vccd1 _14051_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13001_ _13002_/A _13002_/B _13002_/C vssd1 vssd1 vccd1 vccd1 _13003_/A sky130_fd_sc_hd__a21o_1
XFILLER_106_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21622__A1 _13326_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15447__A _19047_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14351__A _14351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21168__B _22852_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20976__A3 _17806_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input42_A wb_dat_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12115__A1 _12116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12115__B2 _18203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17740_ _15941_/X _17817_/A _17652_/Y vssd1 vssd1 vccd1 vccd1 _17743_/D sky130_fd_sc_hd__o21ai_2
XFILLER_43_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14952_ _14952_/A _14952_/B _15002_/B vssd1 vssd1 vccd1 vccd1 _14952_/Y sky130_fd_sc_hd__nand3_2
XFILLER_75_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13903_ _13996_/A _13968_/C _14777_/C _13978_/A vssd1 vssd1 vccd1 vccd1 _13903_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_101_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17671_ _20792_/B vssd1 vssd1 vccd1 vccd1 _21083_/B sky130_fd_sc_hd__buf_2
XFILLER_36_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14883_ _14883_/A _14883_/B _14883_/C vssd1 vssd1 vccd1 vccd1 _14901_/A sky130_fd_sc_hd__nand3_1
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19410_ _19410_/A _19410_/B _19410_/C vssd1 vssd1 vccd1 vccd1 _19422_/A sky130_fd_sc_hd__nand3_2
XANTENNA__15182__A _15182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16622_ _16873_/B vssd1 vssd1 vccd1 vccd1 _16622_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13834_ _13834_/A vssd1 vssd1 vccd1 vccd1 _14112_/A sky130_fd_sc_hd__buf_2
X_19341_ _19336_/X _19334_/X _19512_/A _19521_/A vssd1 vssd1 vccd1 vccd1 _19342_/C
+ sky130_fd_sc_hd__o211ai_4
X_16553_ _16295_/Y _16550_/Y _16552_/Y vssd1 vssd1 vccd1 vccd1 _16554_/A sky130_fd_sc_hd__o21ai_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ _14892_/A _14079_/A _14191_/C _14230_/A _14157_/A vssd1 vssd1 vccd1 vccd1
+ _13765_/X sky130_fd_sc_hd__a32o_1
XANTENNA__11626__B1 _11306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17357__A2 _17227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22350__A2 _22338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_770 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ _16178_/A vssd1 vssd1 vccd1 vccd1 _15504_/X sky130_fd_sc_hd__buf_2
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19272_ _19296_/A _19272_/B _19272_/C vssd1 vssd1 vccd1 vccd1 _19272_/X sky130_fd_sc_hd__and3_1
X_12716_ _12716_/A vssd1 vssd1 vccd1 vccd1 _12716_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_189_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16484_ _11434_/A _16481_/C _22967_/Q vssd1 vssd1 vccd1 vccd1 _16484_/X sky130_fd_sc_hd__o21ba_2
X_13696_ _14107_/A vssd1 vssd1 vccd1 vccd1 _15005_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__11641__A3 _11639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_656 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18223_ _18223_/A vssd1 vssd1 vccd1 vccd1 _18223_/Y sky130_fd_sc_hd__inv_2
X_15435_ _22957_/Q _15435_/B _15435_/C _15435_/D vssd1 vssd1 vccd1 vccd1 _16481_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12647_ _12755_/A _12755_/B _12755_/C vssd1 vssd1 vccd1 vccd1 _12898_/A sky130_fd_sc_hd__nand3_1
XANTENNA__18717__B1_N _18862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17109__A2 _15617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18154_ _12157_/X _12158_/X _15981_/X vssd1 vssd1 vccd1 vccd1 _18154_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16317__B1 _20471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15366_ _15366_/A vssd1 vssd1 vccd1 vccd1 _15378_/A sky130_fd_sc_hd__buf_2
XFILLER_102_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14591__A2 _13746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12578_ _12578_/A vssd1 vssd1 vccd1 vccd1 _17532_/A sky130_fd_sc_hd__buf_4
XFILLER_102_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ _16980_/C _16980_/B _16980_/A vssd1 vssd1 vccd1 vccd1 _17105_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14328__C1 _14327_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14317_ _14354_/A vssd1 vssd1 vccd1 vccd1 _14317_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17837__A _21011_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11529_ _11331_/A _15797_/A _11528_/Y vssd1 vssd1 vccd1 vccd1 _11529_/Y sky130_fd_sc_hd__o21ai_4
X_18085_ _18080_/Y _18081_/Y _18084_/X vssd1 vssd1 vccd1 vccd1 _18087_/A sky130_fd_sc_hd__o21bai_1
X_15297_ _15297_/A vssd1 vssd1 vccd1 vccd1 _15808_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17036_ _17036_/A _17036_/B _17036_/C vssd1 vssd1 vccd1 vccd1 _17038_/B sky130_fd_sc_hd__nand3_1
X_14248_ _14248_/A _14248_/B _14248_/C vssd1 vssd1 vccd1 vccd1 _14250_/B sky130_fd_sc_hd__nand3_1
XANTENNA__20263__A _20263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15357__A _15357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14179_ _14178_/A _14178_/C _14178_/B vssd1 vssd1 vccd1 vccd1 _14180_/C sky130_fd_sc_hd__a21o_1
XFILLER_152_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19019__C1 _18512_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _19156_/D _18984_/Y _18986_/Y vssd1 vssd1 vccd1 vccd1 _19002_/A sky130_fd_sc_hd__o21ai_2
XFILLER_112_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13303__B1 _21584_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _17889_/A _17889_/B _17888_/B vssd1 vssd1 vccd1 vccd1 _17991_/C sky130_fd_sc_hd__o21ai_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19490__C _19490_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater135 _22797_/CLK vssd1 vssd1 vccd1 vccd1 _22795_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__17045__A1 _16880_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18387__B _18387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater146 _22805_/CLK vssd1 vssd1 vccd1 vccd1 _22762_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater157 _22743_/CLK vssd1 vssd1 vccd1 vccd1 _22744_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17869_ _17869_/A vssd1 vssd1 vccd1 vccd1 _17954_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__15804__B _17672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater168 _22733_/CLK vssd1 vssd1 vccd1 vccd1 _22735_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18793__A1 _18770_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19608_ _19608_/A _19608_/B vssd1 vssd1 vccd1 vccd1 _19610_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20880_ _20880_/A _20941_/B vssd1 vssd1 vccd1 vccd1 _20882_/A sky130_fd_sc_hd__nand2_1
X_19539_ _19536_/A _19536_/B _19537_/Y _19538_/X vssd1 vssd1 vccd1 vccd1 _19540_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_35_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18545__A1 _18156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22875__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22550_ _14863_/C input41/X _22558_/S vssd1 vssd1 vccd1 vccd1 _22551_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11632__A3 _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21501_ _21501_/A _21501_/B vssd1 vssd1 vccd1 vccd1 _21508_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22481_ _22481_/A vssd1 vssd1 vccd1 vccd1 _22736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13340__A _13340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21432_ _22674_/Q _21433_/A vssd1 vssd1 vccd1 vccd1 _21432_/X sky130_fd_sc_hd__or2_1
XFILLER_194_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20104__A1 _12697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21852__A1 _21964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17747__A _19774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21363_ _21713_/A _21629_/B _21713_/C vssd1 vssd1 vccd1 vccd1 _21365_/A sky130_fd_sc_hd__nand3_1
XFILLER_107_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20314_ _20314_/A _20314_/B _20314_/C _20442_/A vssd1 vssd1 vccd1 vccd1 _20314_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__21269__A _21269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17466__B _17466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21294_ _22672_/Q _21294_/B _21294_/C _21294_/D vssd1 vssd1 vccd1 vccd1 _21295_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20245_ _20130_/C _16932_/C _16257_/D _16477_/C _20323_/D vssd1 vssd1 vccd1 vccd1
+ _20245_/X sky130_fd_sc_hd__a32o_1
XFILLER_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11699__A3 _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17284__A1 _19336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20176_ _20165_/Y _20181_/B _20175_/Y vssd1 vssd1 vccd1 vccd1 _20184_/A sky130_fd_sc_hd__a21o_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15714__B _15714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16098__A _16098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11880_ _11877_/Y _11879_/Y _12065_/A _11333_/X _11319_/Y vssd1 vssd1 vccd1 vccd1
+ _11883_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22817_ _22850_/CLK hold13/X vssd1 vssd1 vccd1 vccd1 _22817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1112 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18536__A1 _14430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15152__D _15186_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19202__A _19346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ _13550_/A _13550_/B _13550_/C vssd1 vssd1 vccd1 vccd1 _13551_/C sky130_fd_sc_hd__nand3_1
XFILLER_73_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22748_ _22749_/CLK _22748_/D vssd1 vssd1 vccd1 vccd1 _22748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12820__A2 _16779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12501_ _12501_/A vssd1 vssd1 vccd1 vccd1 _12501_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13481_ _13481_/A _13481_/B vssd1 vssd1 vccd1 vccd1 _13484_/C sky130_fd_sc_hd__xnor2_1
X_22679_ _22944_/CLK _22679_/D vssd1 vssd1 vccd1 vccd1 _22679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15220_ _14865_/A _14865_/B _15214_/X _15240_/A _15217_/X vssd1 vssd1 vccd1 vccd1
+ _15224_/D sky130_fd_sc_hd__a2111oi_4
XANTENNA__13250__A _22848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12432_ _12432_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _12432_/Y sky130_fd_sc_hd__nand2_1
X_15151_ _15152_/B _15152_/C _15182_/A _14854_/X vssd1 vssd1 vccd1 vccd1 _15163_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_5_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12363_ _12378_/C vssd1 vssd1 vccd1 vccd1 _12363_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14102_ _14049_/B _14049_/A _14103_/C _14103_/A vssd1 vssd1 vccd1 vccd1 _14104_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ _11411_/A _22955_/Q vssd1 vssd1 vccd1 vccd1 _11315_/B sky130_fd_sc_hd__nand2_1
X_15082_ _15082_/A vssd1 vssd1 vccd1 vccd1 _15149_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12294_ _12294_/A _12294_/B vssd1 vssd1 vccd1 vccd1 _20323_/A sky130_fd_sc_hd__nand2_2
XFILLER_153_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18910_ _19602_/C _19334_/B _18865_/A _18839_/X vssd1 vssd1 vccd1 vccd1 _18912_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_107_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14033_ _14033_/A _14033_/B _14033_/C vssd1 vssd1 vccd1 vccd1 _14033_/X sky130_fd_sc_hd__and3_1
XFILLER_153_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16711__D _17312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19890_ _19890_/A _19890_/B _19893_/A vssd1 vssd1 vccd1 vccd1 _19891_/B sky130_fd_sc_hd__and3_1
XFILLER_107_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18841_ _18841_/A _18841_/B _18841_/C vssd1 vssd1 vccd1 vccd1 _18843_/A sky130_fd_sc_hd__nand3_2
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15905__A _15905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14231__D _15050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18772_ _18772_/A _18772_/B _18772_/C _18772_/D vssd1 vssd1 vccd1 vccd1 _18772_/Y
+ sky130_fd_sc_hd__nand4_2
X_15984_ _15427_/X _12716_/X _15900_/B _15983_/Y vssd1 vssd1 vccd1 vccd1 _16005_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17723_ _17608_/X _17610_/Y _17617_/Y _17508_/Y vssd1 vssd1 vccd1 vccd1 _17723_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__18224__B1 _12221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14935_ _14935_/A vssd1 vssd1 vccd1 vccd1 _15114_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20031__B1 _22926_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22898__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17654_ _17654_/A _17654_/B _17654_/C vssd1 vssd1 vccd1 vccd1 _17660_/A sky130_fd_sc_hd__nand3_1
XFILLER_91_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14866_ _15062_/A _14934_/A _14861_/C _14935_/A vssd1 vssd1 vccd1 vccd1 _14866_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_35_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16605_ _16605_/A _16605_/B vssd1 vssd1 vccd1 vccd1 _16620_/A sky130_fd_sc_hd__nand2_1
X_13817_ _13793_/Y _13826_/B _13815_/X _14122_/A vssd1 vssd1 vccd1 vccd1 _13828_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_189_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17585_ _17585_/A _17585_/B vssd1 vssd1 vccd1 vccd1 _17585_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15994__D1 _17539_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14797_ _14884_/A _14884_/B _14884_/C vssd1 vssd1 vccd1 vccd1 _14805_/D sky130_fd_sc_hd__nand3_2
XFILLER_91_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19324_ _12111_/X _19464_/A _19323_/X _19319_/Y _19320_/X vssd1 vssd1 vccd1 vccd1
+ _19324_/X sky130_fd_sc_hd__o311a_1
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16536_ _16536_/A _16536_/B vssd1 vssd1 vccd1 vccd1 _16536_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13748_ _13748_/A vssd1 vssd1 vccd1 vccd1 _13748_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_189_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19255_ _19250_/Y _19252_/X _19254_/X _19149_/X vssd1 vssd1 vccd1 vccd1 _19255_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_32_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16467_ _16269_/X _16261_/Y _16466_/X vssd1 vssd1 vccd1 vccd1 _16842_/C sky130_fd_sc_hd__a21oi_4
XFILLER_176_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13679_ _13617_/X _13674_/Y _13678_/Y vssd1 vssd1 vccd1 vccd1 _13679_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18206_ _18204_/A _18571_/B _18571_/C vssd1 vssd1 vccd1 vccd1 _18309_/A sky130_fd_sc_hd__nand3b_1
XFILLER_176_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15418_ _20355_/A vssd1 vssd1 vccd1 vccd1 _17108_/B sky130_fd_sc_hd__buf_2
XFILLER_157_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19186_ _18980_/X _18982_/X _19185_/A vssd1 vssd1 vccd1 vccd1 _19187_/B sky130_fd_sc_hd__o21ai_1
XFILLER_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16398_ _16400_/A _21050_/D _16400_/C _16397_/X vssd1 vssd1 vccd1 vccd1 _16398_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_106_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17567__A _17574_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18137_ _19197_/A _18325_/A _18876_/C vssd1 vssd1 vccd1 vccd1 _18137_/Y sky130_fd_sc_hd__nand3_2
XFILLER_157_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15349_ _15342_/Y _15343_/X _15345_/Y _15348_/Y vssd1 vssd1 vccd1 vccd1 _15665_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__16471__A _16471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18068_ _18067_/Y _18049_/B _18063_/X vssd1 vssd1 vccd1 vccd1 _18069_/D sky130_fd_sc_hd__o21bai_1
XFILLER_145_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21047__C1 _21082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17019_ _17019_/A _17019_/B vssd1 vssd1 vccd1 vccd1 _17027_/C sky130_fd_sc_hd__nand2_1
XFILLER_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20030_ _20030_/A vssd1 vssd1 vccd1 vccd1 _20032_/C sky130_fd_sc_hd__inv_2
XFILLER_99_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11550__A2 _11895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15534__B _22962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21981_ _22036_/A _22064_/A _22036_/B _22036_/C vssd1 vssd1 vccd1 vccd1 _21983_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20932_ _17928_/A _20930_/Y _20931_/X vssd1 vssd1 vccd1 vccd1 _20933_/B sky130_fd_sc_hd__o21ai_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20573__A1 _20449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_718 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20863_ _20851_/Y _20863_/B _20863_/C vssd1 vssd1 vccd1 vccd1 _20869_/C sky130_fd_sc_hd__nand3b_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20435__A1_N _20554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15550__A _19507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22602_ _11980_/C input63/X _22608_/S vssd1 vssd1 vccd1 vccd1 _22603_/A sky130_fd_sc_hd__mux2_1
X_20794_ _13022_/B _16746_/X _20791_/Y _20792_/X _20793_/Y vssd1 vssd1 vccd1 vccd1
+ _20797_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16365__B _16627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22533_ _22533_/A vssd1 vssd1 vccd1 vccd1 _22759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22464_ _13304_/B input66/X _22464_/S vssd1 vssd1 vccd1 vccd1 _22465_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14555__A2 _14552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21415_ _21415_/A _21415_/B _21415_/C vssd1 vssd1 vccd1 vccd1 _21421_/A sky130_fd_sc_hd__nand3_2
XFILLER_182_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22395_ _22395_/A vssd1 vssd1 vccd1 vccd1 _22698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19494__A2 _18856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21346_ _13324_/B _13300_/Y _13317_/X _13316_/X vssd1 vssd1 vccd1 vccd1 _21346_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_135_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_984 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_494 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21277_ _13493_/B _13493_/A _13497_/X vssd1 vssd1 vccd1 vccd1 _21278_/C sky130_fd_sc_hd__a21oi_1
XFILLER_78_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20228_ _20228_/A _20228_/B _20228_/C vssd1 vssd1 vccd1 vccd1 _20236_/A sky130_fd_sc_hd__nand3_2
XFILLER_78_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15807__A2 _15691_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20159_ _20293_/B _20161_/B _20167_/B _20167_/A vssd1 vssd1 vccd1 vccd1 _20165_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16480__A2 _17379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12981_ _15577_/D _12981_/B _12981_/C _12981_/D vssd1 vssd1 vccd1 vccd1 _12982_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20013__B1 _18778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _14719_/X _14942_/C _14591_/X vssd1 vssd1 vccd1 vccd1 _14729_/B sky130_fd_sc_hd__o21ai_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ _11932_/A _11932_/B _11932_/C vssd1 vssd1 vccd1 vccd1 _11932_/Y sky130_fd_sc_hd__nand3_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _11859_/X _11861_/X _12065_/A _11399_/Y _11393_/Y vssd1 vssd1 vccd1 vccd1
+ _12074_/B sky130_fd_sc_hd__o2111ai_4
X_14651_ _14750_/B _14651_/B vssd1 vssd1 vccd1 vccd1 _14651_/Y sky130_fd_sc_hd__nand2_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13046__A2 _12894_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19167__D1 _19461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15460__A _15810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _13617_/B _13602_/B vssd1 vssd1 vccd1 vccd1 _13602_/Y sky130_fd_sc_hd__nor2_1
X_17370_ _17370_/A _17370_/B vssd1 vssd1 vccd1 vccd1 _17372_/A sky130_fd_sc_hd__and2_1
XANTENNA__12254__B1 _12251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _11794_/A vssd1 vssd1 vccd1 vccd1 _11976_/A sky130_fd_sc_hd__clkbuf_2
X_14582_ _14863_/B _14593_/B _22764_/Q _13748_/A vssd1 vssd1 vccd1 vccd1 _14590_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16321_ _16435_/B _16579_/A _14369_/X vssd1 vssd1 vccd1 vccd1 _16325_/A sky130_fd_sc_hd__o21ai_2
XFILLER_159_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13533_ _21757_/A _21805_/B _13446_/X _13447_/X vssd1 vssd1 vccd1 vccd1 _13533_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_159_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19040_ _18912_/A _18912_/B _18853_/A vssd1 vssd1 vccd1 vccd1 _19149_/A sky130_fd_sc_hd__a21boi_1
XFILLER_158_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16252_ _15545_/X _15546_/X _16215_/A vssd1 vssd1 vccd1 vccd1 _16253_/A sky130_fd_sc_hd__o21ai_1
X_13464_ _13447_/X _13446_/X _13169_/X vssd1 vssd1 vccd1 vccd1 _13464_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__15743__A1 _15298_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15203_ _15203_/A _15209_/B vssd1 vssd1 vccd1 vccd1 _15205_/C sky130_fd_sc_hd__or2_2
X_12415_ _12415_/A vssd1 vssd1 vccd1 vccd1 _12701_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_166_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16183_ _16183_/A _16183_/B vssd1 vssd1 vccd1 vccd1 _16183_/Y sky130_fd_sc_hd__nand2_1
X_13395_ _13394_/Y _13359_/X _13391_/B vssd1 vssd1 vccd1 vccd1 _13399_/A sky130_fd_sc_hd__a21o_1
XFILLER_182_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15134_ _15134_/A _15134_/B vssd1 vssd1 vccd1 vccd1 _15135_/B sky130_fd_sc_hd__xor2_2
X_12346_ _12314_/Y _12329_/X _20346_/C _12334_/X _20086_/A vssd1 vssd1 vccd1 vccd1
+ _12346_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_126_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15619__B _20098_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19942_ _19454_/C _19322_/B _19322_/C _19901_/B _19896_/A vssd1 vssd1 vccd1 vccd1
+ _19945_/D sky130_fd_sc_hd__a32o_1
XFILLER_141_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15065_ _15060_/X _15065_/B _15065_/C vssd1 vssd1 vccd1 vccd1 _15108_/A sky130_fd_sc_hd__nand3b_2
X_12277_ _12396_/C _12385_/A _12421_/A _12384_/A vssd1 vssd1 vccd1 vccd1 _12279_/B
+ sky130_fd_sc_hd__nand4b_2
XANTENNA__12324__A _22703_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17248__A1 _16778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14016_ _14618_/A _14057_/A _13854_/A vssd1 vssd1 vccd1 vccd1 _14026_/B sky130_fd_sc_hd__o21ai_1
X_19873_ _19921_/A _19921_/B _19872_/Y vssd1 vssd1 vccd1 vccd1 _19875_/A sky130_fd_sc_hd__o21ba_1
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18824_ _18824_/A _18824_/B _18824_/C vssd1 vssd1 vccd1 vccd1 _18824_/X sky130_fd_sc_hd__and3_1
XANTENNA__15635__A _20355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18755_ _18765_/A _18765_/B vssd1 vssd1 vccd1 vccd1 _18764_/B sky130_fd_sc_hd__nand2_1
XANTENNA__15354__B _16322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15967_ _15967_/A _15967_/B _15967_/C vssd1 vssd1 vccd1 vccd1 _15967_/X sky130_fd_sc_hd__and3_1
XFILLER_110_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17706_ _17605_/B _17605_/A _17781_/B vssd1 vssd1 vccd1 vccd1 _17708_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__13155__A _22845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14918_ _14768_/A _14768_/B _14917_/X vssd1 vssd1 vccd1 vccd1 _14919_/C sky130_fd_sc_hd__a21oi_1
X_18686_ _18980_/A _19687_/A _18869_/A _18862_/A vssd1 vssd1 vccd1 vccd1 _18905_/B
+ sky130_fd_sc_hd__nand4_2
X_15898_ _15889_/X _15894_/X _15924_/C _15924_/A vssd1 vssd1 vccd1 vccd1 _15898_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16223__A2 _15450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17637_ _17730_/A _17444_/A _17732_/A _17876_/A vssd1 vssd1 vccd1 vccd1 _17637_/Y
+ sky130_fd_sc_hd__o22ai_1
X_14849_ _14845_/C _14845_/A _14552_/X vssd1 vssd1 vccd1 vccd1 _14928_/A sky130_fd_sc_hd__a21oi_1
XFILLER_36_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17568_ _17385_/Y _17412_/X _17383_/Y vssd1 vssd1 vccd1 vccd1 _17574_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__15982__A1 _12968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21522__D _21522_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19307_ _19396_/A _19396_/B _19396_/C _19192_/Y vssd1 vssd1 vccd1 vccd1 _19394_/A
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__11599__A2 _11598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16519_ _16519_/A _16519_/B _16519_/C vssd1 vssd1 vccd1 vccd1 _16520_/A sky130_fd_sc_hd__nand3_1
XFILLER_143_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20858__A2 _17444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17499_ _17726_/D _17726_/C vssd1 vssd1 vccd1 vccd1 _17853_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18681__A _18681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19238_ _19238_/A _19396_/C vssd1 vssd1 vccd1 vccd1 _19238_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19496__B _19496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22913__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19169_ _12118_/A _12167_/X _19168_/Y vssd1 vssd1 vccd1 vccd1 _19334_/A sky130_fd_sc_hd__o21ai_4
XFILLER_117_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21200_ _13295_/X _21329_/B _13073_/A _13098_/A _14359_/X vssd1 vssd1 vccd1 vccd1
+ _22229_/C sky130_fd_sc_hd__o311ai_4
XFILLER_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22180_ _22105_/X _22186_/A _22113_/B vssd1 vssd1 vccd1 vccd1 _22231_/C sky130_fd_sc_hd__o21ai_1
XFILLER_144_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21131_ _22942_/Q _21122_/X _21127_/B _21130_/Y vssd1 vssd1 vccd1 vccd1 _21150_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__12234__A _15530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1111 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21062_ _21062_/A _21062_/B vssd1 vssd1 vccd1 vccd1 _21095_/B sky130_fd_sc_hd__nand2_1
XFILLER_160_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11523__A2 _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20013_ _18023_/X _19987_/B _18778_/D _19987_/C vssd1 vssd1 vccd1 vccd1 _20013_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15545__A _18203_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20794__A1 _13022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18856__A _18856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21964_ _21964_/A vssd1 vssd1 vccd1 vccd1 _21964_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20915_ _20123_/X _17880_/A _17460_/A _20919_/B _20910_/Y vssd1 vssd1 vccd1 vccd1
+ _20916_/C sky130_fd_sc_hd__o311ai_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21895_ _21933_/A _21996_/A _21933_/B vssd1 vssd1 vccd1 vccd1 _21899_/C sky130_fd_sc_hd__nand3_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ _16585_/A _16585_/B _20790_/Y _12928_/X vssd1 vssd1 vccd1 vccd1 _20920_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15973__A1 _15972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19164__A1 _19162_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19687__A _19687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20849__A2 _17728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20777_ _20772_/B _20775_/Y _20776_/X vssd1 vssd1 vccd1 vccd1 _20839_/A sky130_fd_sc_hd__a21oi_1
XFILLER_196_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22516_ _22584_/S vssd1 vssd1 vccd1 vccd1 _22525_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__15725__A1 _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16922__B1 _15939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20626__A _20626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22447_ _13230_/X input46/X _22453_/S vssd1 vssd1 vccd1 vccd1 _22448_/A sky130_fd_sc_hd__mux2_1
X_12200_ _22963_/Q vssd1 vssd1 vccd1 vccd1 _22662_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_182_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17478__A1 _17466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13180_ _13216_/B _13180_/B vssd1 vssd1 vccd1 vccd1 _13181_/C sky130_fd_sc_hd__nand2_1
XANTENNA__22471__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22378_ _12493_/A input60/X _22380_/S vssd1 vssd1 vccd1 vccd1 _22379_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12131_ _18512_/B _12130_/Y _11974_/Y vssd1 vssd1 vccd1 vccd1 _12131_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__16261__D _17246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21329_ _21329_/A _21329_/B vssd1 vssd1 vccd1 vccd1 _21330_/B sky130_fd_sc_hd__nand2_1
XFILLER_135_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12062_ _12062_/A vssd1 vssd1 vccd1 vccd1 _12116_/A sky130_fd_sc_hd__buf_2
XFILLER_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15455__A _15455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16870_ _16705_/Y _16707_/Y _16856_/Y _16859_/X _16869_/Y vssd1 vssd1 vccd1 vccd1
+ _17042_/A sky130_fd_sc_hd__o221ai_4
XFILLER_104_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20785__A1 _20685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16453__A2 _15341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15821_ _18648_/B vssd1 vssd1 vccd1 vccd1 _19317_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18540_ _18529_/A _18529_/B _18327_/Y vssd1 vssd1 vccd1 vccd1 _18543_/A sky130_fd_sc_hd__a21oi_2
XFILLER_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _15752_/A _15752_/B _15752_/C vssd1 vssd1 vccd1 vccd1 _15752_/X sky130_fd_sc_hd__and3_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _13004_/B _12962_/Y _13004_/A vssd1 vssd1 vccd1 vccd1 _12966_/B sky130_fd_sc_hd__o21ai_1
XFILLER_161_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17402__A1 _15934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _14770_/A _14771_/A _14777_/C vssd1 vssd1 vccd1 vccd1 _14706_/B sky130_fd_sc_hd__and3_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _18471_/A _18471_/B _18471_/C vssd1 vssd1 vccd1 vccd1 _18471_/X sky130_fd_sc_hd__and3_1
X_11915_ _16157_/D _11371_/A _11371_/B _11914_/A _11914_/B vssd1 vssd1 vccd1 vccd1
+ _11918_/A sky130_fd_sc_hd__a311o_1
XANTENNA__19942__A3 _19322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _15680_/A _15680_/B _15680_/C vssd1 vssd1 vccd1 vccd1 _15683_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12895_/A _12895_/B _12895_/C vssd1 vssd1 vccd1 vccd1 _13011_/A sky130_fd_sc_hd__nand3_4
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _17422_/A vssd1 vssd1 vccd1 vccd1 _17422_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__16717__C _20781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _14635_/A _14635_/B _14635_/C vssd1 vssd1 vccd1 vccd1 _14636_/C sky130_fd_sc_hd__a21o_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _12003_/A _11846_/B _15776_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _11846_/Y
+ sky130_fd_sc_hd__nand4_4
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19155__B2 _18984_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22936__CLK _22937_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _17208_/A _17208_/B _17208_/C _17352_/X vssd1 vssd1 vccd1 vccd1 _17353_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_158_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13422__B _22041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _18445_/C _15714_/B _19496_/C _11949_/D vssd1 vssd1 vccd1 vccd1 _11777_/Y
+ sky130_fd_sc_hd__nand4_2
X_14565_ _14565_/A vssd1 vssd1 vccd1 vccd1 _15058_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _16304_/A vssd1 vssd1 vccd1 vccd1 _20593_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13516_ _13563_/A _21591_/B _13581_/A _13516_/D vssd1 vssd1 vccd1 vccd1 _13523_/B
+ sky130_fd_sc_hd__nand4_1
X_17284_ _19336_/A _17833_/B _17833_/C _17449_/A _17293_/B vssd1 vssd1 vccd1 vccd1
+ _17285_/D sky130_fd_sc_hd__a32o_1
XFILLER_186_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14496_ _14001_/Y _14002_/X _14009_/B vssd1 vssd1 vccd1 vccd1 _14497_/B sky130_fd_sc_hd__o21ai_1
X_19023_ _11459_/A _11459_/B _11778_/A _11778_/B _18856_/A vssd1 vssd1 vccd1 vccd1
+ _19023_/X sky130_fd_sc_hd__a221o_4
XFILLER_16_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16235_ _15587_/A _16231_/X _16234_/X vssd1 vssd1 vccd1 vccd1 _16238_/B sky130_fd_sc_hd__a21oi_1
XFILLER_139_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13447_ _13465_/A vssd1 vssd1 vccd1 vccd1 _13447_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20255__B _20255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22462__A1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16166_ _16166_/A _16166_/B _16166_/C vssd1 vssd1 vccd1 vccd1 _16166_/Y sky130_fd_sc_hd__nand3_1
X_13378_ _13650_/A _21632_/A _13367_/Y _13377_/Y vssd1 vssd1 vccd1 vccd1 _13385_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15117_ _15119_/D _15006_/C _15006_/A _15119_/B _15119_/C vssd1 vssd1 vccd1 vccd1
+ _15120_/A sky130_fd_sc_hd__a32o_1
XFILLER_126_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12329_ _12329_/A vssd1 vssd1 vccd1 vccd1 _12329_/X sky130_fd_sc_hd__buf_2
X_16097_ _16041_/X _16044_/Y _16096_/Y vssd1 vssd1 vccd1 vccd1 _16418_/A sky130_fd_sc_hd__o21ai_2
XFILLER_181_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19925_ _19919_/Y _19920_/Y _19962_/B vssd1 vssd1 vccd1 vccd1 _19926_/A sky130_fd_sc_hd__o21ai_4
X_15048_ _15018_/A _15018_/C _15018_/B vssd1 vssd1 vccd1 vccd1 _15076_/A sky130_fd_sc_hd__a21bo_1
XFILLER_123_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19856_ _19856_/A _19856_/B _19913_/A vssd1 vssd1 vccd1 vccd1 _19913_/B sky130_fd_sc_hd__nor3_4
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18807_ _18613_/B _18797_/Y _19455_/C _17525_/D _18798_/Y vssd1 vssd1 vccd1 vccd1
+ _18824_/B sky130_fd_sc_hd__o2111ai_2
X_19787_ _19787_/A _19787_/B _19837_/A vssd1 vssd1 vccd1 vccd1 _19837_/B sky130_fd_sc_hd__nand3_1
X_16999_ _16098_/A _17091_/A _16709_/Y _17081_/A _16994_/Y vssd1 vssd1 vccd1 vccd1
+ _17001_/B sky130_fd_sc_hd__o221ai_4
XFILLER_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18738_ _18645_/Y _18646_/X _18725_/X _18732_/Y _18737_/X vssd1 vssd1 vccd1 vccd1
+ _18738_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18669_ _17427_/X _18371_/X _18536_/Y _18537_/X vssd1 vssd1 vccd1 vccd1 _18669_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_110_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15404__B1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16747__A3 _16727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20700_ _20796_/A _20796_/B _20797_/A vssd1 vssd1 vccd1 vccd1 _20702_/C sky130_fd_sc_hd__nand3_1
XANTENNA__15955__A1 _16400_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21680_ _21680_/A _21680_/B _21680_/C vssd1 vssd1 vccd1 vccd1 _21686_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19146__A1 _22914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20631_ _20631_/A _20631_/B _20631_/C vssd1 vssd1 vccd1 vccd1 _20631_/Y sky130_fd_sc_hd__nand3_2
XFILLER_177_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20562_ _20562_/A _20562_/B _20562_/C vssd1 vssd1 vccd1 vccd1 _20563_/B sky130_fd_sc_hd__nand3_2
XANTENNA__17739__B _19769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22301_ _22301_/A _22301_/B vssd1 vssd1 vccd1 vccd1 _22314_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20493_ _12702_/A _15366_/A _15611_/A _12967_/A vssd1 vssd1 vccd1 vccd1 _20493_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14444__A _16130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22232_ _22232_/A _22232_/B vssd1 vssd1 vccd1 vccd1 _22233_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22453__A1 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22661__A _22661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22163_ _22163_/A _22163_/B vssd1 vssd1 vccd1 vccd1 _22163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21114_ _21138_/A _21138_/B _21138_/C vssd1 vssd1 vccd1 vccd1 _21118_/C sky130_fd_sc_hd__nand3_1
X_22094_ _22094_/A _22094_/B vssd1 vssd1 vccd1 vccd1 _22290_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21045_ _21020_/A _21020_/B _21044_/X vssd1 vssd1 vccd1 vccd1 _21055_/A sky130_fd_sc_hd__a21bo_1
XFILLER_113_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17093__C1 _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11308__A _11308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21724__B _21724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22959__CLK _22959_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16199__A1 _15966_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21947_ _21952_/C _21952_/A _21946_/Y vssd1 vssd1 vccd1 vccd1 _21947_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11699_/X _11689_/A _11648_/Y _11687_/Y vssd1 vssd1 vccd1 vccd1 _11700_/Y
+ sky130_fd_sc_hd__a31oi_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _20478_/C vssd1 vssd1 vccd1 vccd1 _12680_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21878_ _22221_/A _22221_/B _21878_/C vssd1 vssd1 vccd1 vccd1 _21878_/X sky130_fd_sc_hd__and3_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11647_/A _11647_/B _11630_/Y vssd1 vssd1 vccd1 vccd1 _11698_/A sky130_fd_sc_hd__a21o_1
XANTENNA__16256__D _16256_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ _20840_/A _20840_/B _20994_/A _20907_/A vssd1 vssd1 vccd1 vccd1 _20902_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19688__A2 _19689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11562_ _11668_/A _11720_/A _11560_/C vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__a21o_2
XFILLER_11_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14350_ _22761_/Q _14330_/X _14337_/X _13304_/B _14349_/X vssd1 vssd1 vccd1 vccd1
+ _14350_/X sky130_fd_sc_hd__a221o_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17649__B _20928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18360__A2 _17422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13301_ _13301_/A vssd1 vssd1 vccd1 vccd1 _13301_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14281_ _14281_/A _14281_/B _14281_/C vssd1 vssd1 vccd1 vccd1 _14281_/Y sky130_fd_sc_hd__nand3_1
XFILLER_196_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11493_ _18130_/C _18797_/C _18453_/C _16078_/C vssd1 vssd1 vccd1 vccd1 _11493_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_109_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16020_ _16093_/B _16020_/B vssd1 vssd1 vccd1 vccd1 _16020_/Y sky130_fd_sc_hd__nand2_1
X_13232_ _13504_/B vssd1 vssd1 vccd1 vccd1 _13633_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input72_A x[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ _13164_/A _13385_/A _13384_/A vssd1 vssd1 vccd1 vccd1 _13286_/C sky130_fd_sc_hd__a21o_1
XFILLER_152_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19583__C _19687_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12114_ _16921_/A vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__16674__A2 _17227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17971_ _17918_/B _17969_/Y _17970_/Y vssd1 vssd1 vccd1 vccd1 _17972_/B sky130_fd_sc_hd__a21oi_1
XFILLER_112_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13094_ _13319_/A _13125_/A _13316_/A vssd1 vssd1 vccd1 vccd1 _13322_/A sky130_fd_sc_hd__o21ai_2
XFILLER_111_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19710_ _19608_/B _19684_/X _19685_/X _19707_/Y _19864_/A vssd1 vssd1 vccd1 vccd1
+ _19720_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12045_ _19197_/D vssd1 vssd1 vccd1 vccd1 _19490_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16922_ _15792_/C _15792_/A _16921_/X _15939_/A _16016_/A vssd1 vssd1 vccd1 vccd1
+ _16922_/X sky130_fd_sc_hd__o32a_2
XANTENNA__15185__A _15213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19073__B1 _19585_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21955__B1 _21724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19641_ _19488_/A _19636_/X _19637_/Y _19635_/A _19724_/B vssd1 vssd1 vccd1 vccd1
+ _19641_/X sky130_fd_sc_hd__o2111a_1
XFILLER_78_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16853_ _16853_/A _16853_/B _16853_/C vssd1 vssd1 vccd1 vccd1 _16853_/X sky130_fd_sc_hd__and3_1
XANTENNA__18281__D1 _19358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22510__S _22512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15804_ _19012_/D _17672_/A _15804_/C _16067_/B vssd1 vssd1 vccd1 vccd1 _15804_/Y
+ sky130_fd_sc_hd__nand4_1
X_19572_ _22917_/Q _19449_/A _19449_/B _19452_/B _19452_/A vssd1 vssd1 vccd1 vccd1
+ _19574_/C sky130_fd_sc_hd__a32o_1
X_16784_ _16778_/X _16779_/X _16792_/A _19694_/A vssd1 vssd1 vccd1 vccd1 _16784_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13996_ _13996_/A vssd1 vssd1 vccd1 vccd1 _14889_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18523_ _18726_/A _18726_/B _18916_/B _18522_/Y vssd1 vssd1 vccd1 vccd1 _18523_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_92_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735_ _15740_/B _15740_/C _15740_/A _15709_/Y _15734_/X vssd1 vssd1 vccd1 vccd1
+ _15862_/A sky130_fd_sc_hd__a32o_1
XFILLER_19_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12947_ _17144_/A vssd1 vssd1 vccd1 vccd1 _15991_/B sky130_fd_sc_hd__buf_4
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22380__A0 _12387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12975__C _16106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18454_ _18451_/Y _18452_/X _18453_/X vssd1 vssd1 vccd1 vccd1 _18458_/A sky130_fd_sc_hd__o21ai_1
XFILLER_179_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15666_ _15666_/A _15668_/A vssd1 vssd1 vccd1 vccd1 _15673_/A sky130_fd_sc_hd__nor2_1
XANTENNA__15937__A1 _15932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19128__A1 _19113_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15937__B2 _15936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20391__C1 _20263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ _12886_/B vssd1 vssd1 vccd1 vccd1 _12878_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17405_ _17405_/A vssd1 vssd1 vccd1 vccd1 _18303_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _15058_/C _14765_/C _14765_/A _14616_/Y _14614_/Y vssd1 vssd1 vccd1 vccd1
+ _14621_/C sky130_fd_sc_hd__a32o_1
X_18385_ _18384_/Y _18173_/C _18163_/Y _18187_/B vssd1 vssd1 vccd1 vccd1 _18385_/Y
+ sky130_fd_sc_hd__a22oi_2
X_11829_ _11829_/A _11829_/B _11829_/C vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__nand3_1
XFILLER_92_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12049__A _19197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15597_ _15597_/A _15597_/B vssd1 vssd1 vccd1 vccd1 _15597_/Y sky130_fd_sc_hd__nand2_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17336_ _17331_/Y _17332_/Y _17333_/Y _17335_/Y vssd1 vssd1 vccd1 vccd1 _17337_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14548_ _14548_/A _14661_/B vssd1 vssd1 vccd1 vccd1 _14549_/B sky130_fd_sc_hd__nor2b_2
XANTENNA__20266__A _20266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11888__A _15912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17267_ _17239_/Y _17236_/X _17242_/Y _17298_/B _17268_/B vssd1 vssd1 vccd1 vccd1
+ _17272_/A sky130_fd_sc_hd__o2111ai_1
XANTENNA__16362__A1 _15646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14479_ _14721_/B vssd1 vssd1 vccd1 vccd1 _14494_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_174_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19006_ _19179_/C _19007_/B _19185_/A _19187_/C vssd1 vssd1 vccd1 vccd1 _19009_/C
+ sky130_fd_sc_hd__o211ai_2
X_16218_ _16218_/A vssd1 vssd1 vccd1 vccd1 _18193_/A sky130_fd_sc_hd__buf_2
XANTENNA__16587__A1_N _16599_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17198_ _17025_/B _17025_/C _17009_/X vssd1 vssd1 vccd1 vccd1 _17198_/X sky130_fd_sc_hd__a21o_1
XFILLER_162_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12923__A1 _13022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16149_ _16186_/A _16186_/B _16145_/Y _16148_/Y vssd1 vssd1 vccd1 vccd1 _16183_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_6_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21809__B _21809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19908_ _19909_/C _19909_/A _19909_/B _19907_/Y _19851_/B vssd1 vssd1 vccd1 vccd1
+ _19908_/X sky130_fd_sc_hd__o311a_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19603__A2 _19769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18811__B1 _18626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19839_ _19899_/A _19839_/B _19839_/C _19839_/D vssd1 vssd1 vccd1 vccd1 _19842_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_110_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22850_ _22850_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 _22850_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19140__B1_N _22915_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21801_ _21801_/A _21801_/B vssd1 vssd1 vccd1 vccd1 _21802_/A sky130_fd_sc_hd__xor2_2
X_22781_ _22813_/CLK _22781_/D vssd1 vssd1 vccd1 vccd1 _22781_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21174__A1 _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13651__A2 _21757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_695 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21732_ _21732_/A _21777_/B vssd1 vssd1 vccd1 vccd1 _21737_/B sky130_fd_sc_hd__nand2_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21663_ _21658_/X _21660_/Y _21661_/Y _21662_/Y vssd1 vssd1 vccd1 vccd1 _21664_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19030__A _19504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20614_ _20482_/A _20482_/B _20486_/X vssd1 vssd1 vccd1 vccd1 _20614_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_196_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21594_ _21739_/C _21738_/A vssd1 vssd1 vccd1 vccd1 _21594_/Y sky130_fd_sc_hd__nand2_2
XFILLER_177_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18342__A2 _19464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__A2 _11774_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20545_ _20545_/A vssd1 vssd1 vccd1 vccd1 _20545_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13167__A1 _13340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20476_ _20579_/A _20579_/B _12680_/X _20481_/C _16304_/A vssd1 vssd1 vccd1 vccd1
+ _20476_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22215_ _22215_/A _22215_/B vssd1 vssd1 vccd1 vccd1 _22216_/B sky130_fd_sc_hd__and2_1
XFILLER_193_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17100__A2_N _17341_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22146_ _22146_/A vssd1 vssd1 vccd1 vccd1 _22212_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14667__A1 _14843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22077_ _22080_/B _22163_/A _22163_/B vssd1 vssd1 vccd1 vccd1 _22081_/A sky130_fd_sc_hd__nand3b_1
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17066__C1 _17373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21028_ _20987_/A _20986_/A _20985_/Y vssd1 vssd1 vccd1 vccd1 _21030_/A sky130_fd_sc_hd__o21a_1
XFILLER_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11350__B1 _11349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ _13821_/B _13892_/A _13896_/A _13869_/B vssd1 vssd1 vccd1 vccd1 _13851_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12801_ _20089_/A _20605_/B vssd1 vssd1 vccd1 vccd1 _15637_/A sky130_fd_sc_hd__nand2_2
XANTENNA__15452__B _17280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13781_ _13781_/A _14043_/A _14199_/A _15008_/C vssd1 vssd1 vccd1 vccd1 _14043_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_90_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22362__B1 _22368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15520_ _15859_/A _15859_/B _15859_/D vssd1 vssd1 vccd1 vccd1 _15679_/B sky130_fd_sc_hd__nand3_1
XFILLER_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12710_/Y _12724_/Y _12739_/C _12739_/A vssd1 vssd1 vccd1 vccd1 _12732_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_163_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _15893_/C vssd1 vssd1 vccd1 vccd1 _15997_/C sky130_fd_sc_hd__buf_2
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_996 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16592__A1 _15936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12663_ _15746_/B vssd1 vssd1 vccd1 vccd1 _16160_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_31_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _22709_/Q _14370_/X _14396_/X _22741_/Q _14401_/X vssd1 vssd1 vccd1 vccd1
+ _14402_/X sky130_fd_sc_hd__a221o_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18170_ _19329_/D vssd1 vssd1 vccd1 vccd1 _18980_/A sky130_fd_sc_hd__buf_2
X_11614_ _11606_/X _18665_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _11614_/Y sky130_fd_sc_hd__nand3b_2
X_15382_ _15389_/B _15382_/B _16062_/A _17530_/A vssd1 vssd1 vccd1 vccd1 _15665_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_169_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20086__A _20086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12594_ _15558_/C _20130_/B _12610_/A vssd1 vssd1 vccd1 vccd1 _12594_/Y sky130_fd_sc_hd__nand3_1
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ _17732_/A _16015_/A _17116_/B _17116_/A vssd1 vssd1 vccd1 vccd1 _17122_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_184_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21873__C1 _22173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14333_ _13725_/A _14330_/X _14313_/X _13202_/A _14332_/X vssd1 vssd1 vccd1 vccd1
+ _14333_/X sky130_fd_sc_hd__a221o_2
X_11545_ _11578_/A _11581_/A _11529_/Y _19061_/A _16106_/C vssd1 vssd1 vccd1 vccd1
+ _11645_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17052_ _16896_/Y _16644_/Y _17050_/X _17049_/Y vssd1 vssd1 vccd1 vccd1 _17053_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_13_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14264_ _14203_/X _14185_/X _14214_/Y _14206_/Y vssd1 vssd1 vccd1 vccd1 _14267_/B
+ sky130_fd_sc_hd__o211ai_1
X_11476_ _11894_/A _11894_/B vssd1 vssd1 vccd1 vccd1 _11895_/A sky130_fd_sc_hd__nand2_2
XFILLER_171_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11708__A2 _11503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16003_ _16003_/A _16003_/B _16003_/C vssd1 vssd1 vccd1 vccd1 _16133_/B sky130_fd_sc_hd__nand3_1
XFILLER_109_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13215_ _13215_/A _13215_/B vssd1 vssd1 vccd1 vccd1 _13475_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21629__B _21629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14195_ _14195_/A _14953_/A _14212_/D _14195_/D vssd1 vssd1 vccd1 vccd1 _14198_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_98_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13146_ _13158_/A _13161_/A _13157_/A _13112_/C vssd1 vssd1 vccd1 vccd1 _13147_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17954_ _17954_/A _17954_/B vssd1 vssd1 vccd1 vccd1 _17954_/X sky130_fd_sc_hd__or2_1
XFILLER_151_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _21188_/C vssd1 vssd1 vccd1 vccd1 _13302_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_183_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16905_ _16905_/A _16905_/B vssd1 vssd1 vccd1 vccd1 _22954_/D sky130_fd_sc_hd__nor2_2
X_12028_ _12054_/A _12054_/B _12089_/A _12088_/A vssd1 vssd1 vccd1 vccd1 _12028_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17885_ _17885_/A _17885_/B vssd1 vssd1 vccd1 vccd1 _17886_/C sky130_fd_sc_hd__nand2_1
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16836_ _19615_/C _20806_/C _16452_/X _16825_/X vssd1 vssd1 vccd1 vccd1 _16836_/X
+ sky130_fd_sc_hd__a31o_1
X_19624_ _19624_/A vssd1 vssd1 vccd1 vccd1 _19941_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19555_ _19555_/A _19555_/B _19555_/C _19555_/D vssd1 vssd1 vccd1 vccd1 _19577_/A
+ sky130_fd_sc_hd__nand4_1
X_16767_ _16494_/X _16760_/X _16954_/A _15577_/D _19687_/B vssd1 vssd1 vccd1 vccd1
+ _16768_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_111_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13979_ _14002_/B _14230_/A _14191_/A _14002_/C vssd1 vssd1 vccd1 vccd1 _14009_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_62_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18506_ _18876_/B vssd1 vssd1 vccd1 vccd1 _18999_/A sky130_fd_sc_hd__clkbuf_2
X_15718_ _15718_/A vssd1 vssd1 vccd1 vccd1 _15723_/A sky130_fd_sc_hd__buf_2
XFILLER_0_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19486_ _19486_/A _19486_/B vssd1 vssd1 vccd1 vccd1 _19536_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19769__B _19769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16698_ _16698_/A _16698_/B _16698_/C vssd1 vssd1 vccd1 vccd1 _16698_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__12841__B1 _12718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18437_ _18774_/A vssd1 vssd1 vccd1 vccd1 _18437_/Y sky130_fd_sc_hd__inv_2
X_15649_ _16078_/C vssd1 vssd1 vccd1 vccd1 _15649_/X sky130_fd_sc_hd__buf_2
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16583__A1 _14369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19506__D1 _19651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18368_ _18367_/A _18367_/B _12018_/X _16921_/X vssd1 vssd1 vccd1 vccd1 _18368_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__22656__A1 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17319_ _17520_/A _17523_/A _17520_/C _17520_/D vssd1 vssd1 vccd1 vccd1 _17466_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__16335__A1 _16310_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18299_ _15538_/X _15541_/X _18778_/A vssd1 vssd1 vccd1 vccd1 _18299_/X sky130_fd_sc_hd__a21o_1
XANTENNA__20131__A2 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19000__D _19614_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14346__B1 _14337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20330_ _20508_/A _15909_/A _20323_/Y _20324_/Y vssd1 vssd1 vccd1 vccd1 _20447_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_174_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19826__A_N _22921_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20261_ _20261_/A vssd1 vssd1 vccd1 vccd1 _20264_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19824__A2 _19294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14722__A _14722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16099__B1 _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22000_ _21841_/A _21341_/X _21841_/B _21841_/C _21897_/B vssd1 vssd1 vccd1 vccd1
+ _22000_/X sky130_fd_sc_hd__o41a_1
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20192_ _20192_/A _20192_/B vssd1 vssd1 vccd1 vccd1 _22910_/D sky130_fd_sc_hd__xor2_4
XFILLER_170_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18848__B _19351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11332__B1 _11372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22902_ _22951_/CLK _22902_/D vssd1 vssd1 vccd1 vccd1 _22902_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__17063__A2 _17227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15553__A _19358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19025__A _19461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22833_ _22850_/CLK _22845_/Q vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__18864__A _19507_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22764_ _22765_/CLK _22764_/D vssd1 vssd1 vccd1 vccd1 _22764_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21715_ _13344_/X _13345_/X _21269_/A vssd1 vssd1 vccd1 vccd1 _21719_/A sky130_fd_sc_hd__a21o_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22695_ _22696_/CLK _22695_/D vssd1 vssd1 vccd1 vccd1 _22695_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13388__A1 _13339_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21646_ _21645_/A _21763_/A _21620_/X _21622_/X vssd1 vssd1 vccd1 vccd1 _21646_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_36_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14616__B _14721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19695__A _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21577_ _21530_/A _21539_/Y _21537_/Y _21538_/Y vssd1 vssd1 vccd1 vccd1 _21680_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__12060__B2 _11565_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11330_ _11371_/A _11371_/B vssd1 vssd1 vccd1 vccd1 _11331_/A sky130_fd_sc_hd__nand2_1
X_20528_ _20378_/Y _20381_/Y _20396_/B _20388_/Y vssd1 vssd1 vccd1 vccd1 _20531_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_181_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15728__A _15988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20459_ _20371_/A _20371_/B _20458_/Y _20353_/A vssd1 vssd1 vccd1 vccd1 _20459_/Y
+ sky130_fd_sc_hd__a22oi_4
X_13000_ _13037_/B _12996_/X _13037_/A vssd1 vssd1 vccd1 vccd1 _13000_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22129_ _22129_/A _22129_/B _22129_/C _22170_/A vssd1 vssd1 vccd1 vccd1 _22170_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12115__A2 _12111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input35_A wb_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14951_ _14951_/A _15002_/A _14951_/C _15061_/A vssd1 vssd1 vccd1 vccd1 _15002_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13902_ _13902_/A _13902_/B vssd1 vssd1 vccd1 vccd1 _13978_/A sky130_fd_sc_hd__nand2_2
X_17670_ _20792_/A vssd1 vssd1 vccd1 vccd1 _21083_/A sky130_fd_sc_hd__buf_2
X_14882_ _14879_/Y _14880_/X _14887_/C vssd1 vssd1 vccd1 vccd1 _14883_/C sky130_fd_sc_hd__o21ai_1
XFILLER_36_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16262__B1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16621_ _16370_/B _16377_/B _16377_/C _16606_/X vssd1 vssd1 vccd1 vccd1 _16625_/A
+ sky130_fd_sc_hd__a31o_1
X_13833_ _13897_/A _13833_/B _13833_/C vssd1 vssd1 vccd1 vccd1 _13833_/X sky130_fd_sc_hd__and3_2
XFILLER_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_610 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14079__A _14079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19340_ _19340_/A _19340_/B vssd1 vssd1 vccd1 vccd1 _19342_/B sky130_fd_sc_hd__nor2_2
X_16552_ _16552_/A _16714_/A vssd1 vssd1 vccd1 vccd1 _16552_/Y sky130_fd_sc_hd__nand2_2
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_654 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13764_ _14203_/A vssd1 vssd1 vccd1 vccd1 _14157_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15503_ _15597_/B _15596_/A _15597_/A vssd1 vssd1 vccd1 vccd1 _15510_/B sky130_fd_sc_hd__nand3_2
XFILLER_44_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19271_ _19269_/Y _19121_/A _19299_/B vssd1 vssd1 vccd1 vccd1 _19271_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12715_ _12689_/X _12712_/Y _12714_/Y vssd1 vssd1 vccd1 vccd1 _12933_/C sky130_fd_sc_hd__o21ai_2
X_16483_ _16483_/A _16483_/B vssd1 vssd1 vccd1 vccd1 _17139_/A sky130_fd_sc_hd__nand2_2
XANTENNA__16565__A1 _15617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20361__A2 _20511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13695_ _22872_/Q vssd1 vssd1 vccd1 vccd1 _14107_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__22677__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18222_ _18214_/X _18215_/Y _18220_/Y _18221_/X vssd1 vssd1 vccd1 vccd1 _18275_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_176_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15434_ _15445_/A _15445_/B _12758_/A vssd1 vssd1 vccd1 vccd1 _15755_/A sky130_fd_sc_hd__a21o_4
XFILLER_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12646_ _12644_/Y _12645_/X _12510_/A _12510_/B vssd1 vssd1 vccd1 vccd1 _12755_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_157_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12051__A1 _11932_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18153_ _18132_/Y _18136_/X _18383_/A _18383_/B vssd1 vssd1 vccd1 vccd1 _18163_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_15_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16317__A1 _15904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15365_ _20101_/A _20101_/B vssd1 vssd1 vccd1 vccd1 _15366_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12577_ _12577_/A vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__buf_4
XFILLER_129_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17104_ _17196_/A _17196_/B vssd1 vssd1 vccd1 vccd1 _17200_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _14411_/A vssd1 vssd1 vccd1 vccd1 _14354_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14328__B1 _14313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18084_ _18084_/A _18084_/B vssd1 vssd1 vccd1 vccd1 _18084_/X sky130_fd_sc_hd__and2_1
XFILLER_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11528_ _12003_/B _18691_/C _12003_/A vssd1 vssd1 vccd1 vccd1 _11528_/Y sky130_fd_sc_hd__nand3_4
XFILLER_184_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15296_ _22887_/Q _15296_/B vssd1 vssd1 vccd1 vccd1 _22875_/D sky130_fd_sc_hd__xor2_1
XFILLER_171_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17035_ _17036_/A _17036_/B _17036_/C vssd1 vssd1 vccd1 vccd1 _17038_/A sky130_fd_sc_hd__a21o_1
X_14247_ _14253_/A _14253_/B vssd1 vssd1 vccd1 vccd1 _14250_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11459_ _11459_/A _11459_/B vssd1 vssd1 vccd1 vccd1 _11506_/A sky130_fd_sc_hd__nand2_4
XANTENNA__20263__B _20263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15357__B _20355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ _14178_/A _14178_/B _14178_/C vssd1 vssd1 vccd1 vccd1 _14180_/B sky130_fd_sc_hd__nand3_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19019__B1 _18512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _13112_/Y _13097_/A _13055_/A vssd1 vssd1 vccd1 vccd1 _13449_/A sky130_fd_sc_hd__a21o_1
XFILLER_112_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18986_ _15797_/A _19160_/A _18985_/Y vssd1 vssd1 vccd1 vccd1 _18986_/Y sky130_fd_sc_hd__o21ai_4
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _17991_/A _17991_/B vssd1 vssd1 vccd1 vccd1 _17939_/A sky130_fd_sc_hd__nand2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21377__A1 _21376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19490__D _19490_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater136 _22789_/CLK vssd1 vssd1 vccd1 vccd1 _22797_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__17045__A2 _16879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18387__C _18387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater147 _22772_/CLK vssd1 vssd1 vccd1 vccd1 _22805_/CLK sky130_fd_sc_hd__clkbuf_1
X_17868_ _17868_/A _17868_/B vssd1 vssd1 vccd1 vccd1 _22962_/D sky130_fd_sc_hd__nor2_1
Xrepeater158 _22742_/CLK vssd1 vssd1 vccd1 vccd1 _22743_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_27_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15804__C _15804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater169 _22731_/CLK vssd1 vssd1 vccd1 vccd1 _22733_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19607_ _19607_/A _19607_/B vssd1 vssd1 vccd1 vccd1 _19608_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16819_ _18848_/C _20928_/A _20928_/B vssd1 vssd1 vccd1 vccd1 _16819_/X sky130_fd_sc_hd__and3_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17799_ _17799_/A _17799_/B vssd1 vssd1 vccd1 vccd1 _17910_/A sky130_fd_sc_hd__nand2_2
XFILLER_35_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11406__A _22957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19538_ _19538_/A _19538_/B _19538_/C vssd1 vssd1 vccd1 vccd1 _19538_/X sky130_fd_sc_hd__and3_1
XFILLER_62_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18545__A2 _16276_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11908__A1_N _11909_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19469_ _19476_/C _19476_/A _18514_/Y _19308_/X vssd1 vssd1 vccd1 vccd1 _19479_/B
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_62_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16556__A1 _16098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21500_ _21716_/A _21640_/A _21499_/X vssd1 vssd1 vccd1 vccd1 _21501_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22480_ _22736_/Q input42/X _22486_/S vssd1 vssd1 vccd1 vccd1 _22481_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21431_ _21431_/A _21431_/B vssd1 vssd1 vccd1 vccd1 _21433_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20104__A2 _16300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16932__A _18445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12237__A _15531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11779__C _11779_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14582__A3 _22764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12593__A2 _20471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21362_ _21362_/A _21362_/B _21724_/C _21724_/B vssd1 vssd1 vccd1 vccd1 _21372_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_135_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20313_ _20313_/A _20562_/A vssd1 vssd1 vccd1 vccd1 _20317_/A sky130_fd_sc_hd__nand2_2
XFILLER_163_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput80 x[9] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_1
X_21293_ _22672_/Q _21294_/B _21294_/C _21294_/D vssd1 vssd1 vccd1 vccd1 _21295_/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17466__C _17467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16370__C _16377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20244_ _20244_/A vssd1 vssd1 vccd1 vccd1 _20244_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18859__A _19480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17284__A2 _17833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20175_ _12886_/A _12878_/X _12781_/B vssd1 vssd1 vccd1 vccd1 _20175_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12502__C1 _20486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12700__A _15774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15714__C _16515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22816_ _22943_/CLK _22816_/D vssd1 vssd1 vccd1 vccd1 _22816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_719 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17339__A3 _17341_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18536__A2 _15297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19202__B _19507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22747_ _22747_/CLK _22747_/D vssd1 vssd1 vccd1 vccd1 _22747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12500_ _12500_/A vssd1 vssd1 vccd1 vccd1 _12500_/X sky130_fd_sc_hd__buf_4
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13480_ _13396_/X _13290_/B _13478_/X _13479_/X vssd1 vssd1 vccd1 vccd1 _13556_/C
+ sky130_fd_sc_hd__o211ai_2
X_22678_ _22944_/CLK _22678_/D vssd1 vssd1 vccd1 vccd1 _22678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12569__C1 _16319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12033__A1 _11693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ _12417_/X _12425_/X _12429_/X _12430_/Y vssd1 vssd1 vccd1 vccd1 _12432_/B
+ sky130_fd_sc_hd__o22ai_4
X_21629_ _21724_/A _21629_/B _21724_/D vssd1 vssd1 vccd1 vccd1 _21629_/Y sky130_fd_sc_hd__nand3_1
XFILLER_32_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12147__A _22792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15150_ _15146_/Y _15122_/X _15217_/A _15006_/C _15006_/A vssd1 vssd1 vccd1 vccd1
+ _15152_/C sky130_fd_sc_hd__o2111ai_2
XANTENNA__21843__A2 _21733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ _22697_/Q vssd1 vssd1 vccd1 vccd1 _12378_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_165_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14101_ _14093_/Y _14178_/B _14178_/C _14099_/Y _14100_/X vssd1 vssd1 vccd1 vccd1
+ _14103_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_181_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11313_ _11404_/B _11404_/C _11404_/D _11311_/Y _11713_/B vssd1 vssd1 vccd1 vccd1
+ _11316_/A sky130_fd_sc_hd__o311ai_2
XFILLER_180_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15081_ _15080_/Y _15017_/A _15082_/A vssd1 vssd1 vccd1 vccd1 _15081_/X sky130_fd_sc_hd__o21a_1
X_12293_ _16267_/A _12413_/A vssd1 vssd1 vccd1 vccd1 _12294_/B sky130_fd_sc_hd__nand2_4
XFILLER_181_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13533__A1 _21757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14032_ _14032_/A vssd1 vssd1 vccd1 vccd1 _14099_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17673__A _19334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18840_ _19504_/D _19013_/C _18865_/A _18839_/X vssd1 vssd1 vccd1 vccd1 _19091_/B
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__18472__A1 _12064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14512__D _15058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18771_ _18769_/Y _18770_/X _18774_/D _18587_/B vssd1 vssd1 vccd1 vccd1 _18783_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15983_ _11904_/X _11905_/X _15810_/C vssd1 vssd1 vccd1 vccd1 _15983_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_95_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17722_ _17722_/A _17722_/B vssd1 vssd1 vccd1 vccd1 _17722_/Y sky130_fd_sc_hd__nand2_1
X_14934_ _14934_/A _15154_/D vssd1 vssd1 vccd1 vccd1 _14934_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15624__C _20678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17653_ _15941_/X _17822_/A _17535_/B _17652_/Y _17648_/Y vssd1 vssd1 vccd1 vccd1
+ _17654_/C sky130_fd_sc_hd__o221ai_1
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14865_ _14865_/A _14865_/B vssd1 vssd1 vccd1 vccd1 _15062_/A sky130_fd_sc_hd__nand2_1
XFILLER_63_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17983__B1 _17039_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16604_ _16873_/A _16601_/Y _16603_/Y vssd1 vssd1 vccd1 vccd1 _16605_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13816_ _22867_/Q vssd1 vssd1 vccd1 vccd1 _14122_/A sky130_fd_sc_hd__clkinv_2
X_17584_ _17701_/C _17585_/B _17579_/Y _17583_/Y vssd1 vssd1 vccd1 vccd1 _17584_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14796_ _14884_/B _14884_/C _14884_/A vssd1 vssd1 vccd1 vccd1 _14805_/C sky130_fd_sc_hd__a21o_1
XFILLER_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19323_ _19323_/A vssd1 vssd1 vccd1 vccd1 _19323_/X sky130_fd_sc_hd__buf_2
XFILLER_189_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16535_ _16535_/A _16535_/B vssd1 vssd1 vccd1 vccd1 _16536_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13747_ _22865_/Q vssd1 vssd1 vccd1 vccd1 _13748_/A sky130_fd_sc_hd__inv_2
XFILLER_188_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19254_ _19254_/A _19254_/B _19254_/C vssd1 vssd1 vccd1 vccd1 _19254_/X sky130_fd_sc_hd__and3_1
X_16466_ _12118_/A _15903_/X _20255_/A _16921_/A _12696_/X vssd1 vssd1 vccd1 vccd1
+ _16466_/X sky130_fd_sc_hd__o32a_1
X_13678_ _13678_/A _13678_/B _13678_/C vssd1 vssd1 vccd1 vccd1 _13678_/Y sky130_fd_sc_hd__nand3_1
X_18205_ _18402_/B _18402_/A vssd1 vssd1 vccd1 vccd1 _18207_/A sky130_fd_sc_hd__nand2_1
X_15417_ _20611_/A vssd1 vssd1 vccd1 vccd1 _17131_/B sky130_fd_sc_hd__clkbuf_4
X_19185_ _19185_/A _19185_/B _19185_/C vssd1 vssd1 vccd1 vccd1 _19240_/A sky130_fd_sc_hd__nand3_2
X_12629_ _12630_/A _12630_/B _12630_/C vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__a21o_1
XFILLER_192_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16397_ _16397_/A vssd1 vssd1 vccd1 vccd1 _16397_/X sky130_fd_sc_hd__buf_2
XFILLER_157_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18136_ _15887_/A _18365_/A _19464_/A _18131_/X _18125_/X vssd1 vssd1 vccd1 vccd1
+ _18136_/X sky130_fd_sc_hd__o311a_1
X_15348_ _15315_/Y _15343_/X _15347_/X vssd1 vssd1 vccd1 vccd1 _15348_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17567__B _17574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18067_ _18067_/A vssd1 vssd1 vccd1 vccd1 _18067_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16710__A1 _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15279_ _15279_/A _22878_/Q _22879_/Q _22880_/Q vssd1 vssd1 vccd1 vccd1 _15287_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_176_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17018_ _17027_/A _17027_/B vssd1 vssd1 vccd1 vccd1 _17020_/A sky130_fd_sc_hd__nand2_1
XFILLER_160_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11535__B1 _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20270__A1 _20115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _18969_/A _18969_/B vssd1 vssd1 vccd1 vccd1 _18969_/X sky130_fd_sc_hd__or2_1
XANTENNA__22547__A0 _22766_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22842__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15534__C _22662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21980_ _21892_/A _21892_/C _21934_/Y vssd1 vssd1 vccd1 vccd1 _21983_/A sky130_fd_sc_hd__a21oi_1
XFILLER_54_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20931_ _20806_/B _17816_/B _20930_/A vssd1 vssd1 vccd1 vccd1 _20931_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20573__A2 _20728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15831__A _16809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20862_ _20866_/A _20866_/B _20864_/B vssd1 vssd1 vccd1 vccd1 _20863_/C sky130_fd_sc_hd__a21bo_1
XFILLER_148_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_760 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20449__A _20449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19715__A1 _19793_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22601_ _22601_/A vssd1 vssd1 vccd1 vccd1 _22789_/D sky130_fd_sc_hd__clkbuf_1
X_20793_ _20793_/A _20793_/B _20793_/C _20793_/D vssd1 vssd1 vccd1 vccd1 _20793_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16365__C _16369_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22532_ _13736_/C input64/X _22536_/S vssd1 vssd1 vccd1 vccd1 _22533_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_908 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22463_ _22463_/A vssd1 vssd1 vccd1 vccd1 _22728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21414_ _21411_/A _21417_/B _21416_/A vssd1 vssd1 vccd1 vccd1 _21415_/C sky130_fd_sc_hd__a21o_1
XFILLER_182_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22394_ _16322_/A input36/X _22402_/S vssd1 vssd1 vccd1 vccd1 _22395_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21345_ _21386_/A _21386_/B _21342_/X _21344_/X vssd1 vssd1 vccd1 vccd1 _21387_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_108_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_996 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21276_ _21281_/A _21419_/A _21276_/C vssd1 vssd1 vccd1 vccd1 _21278_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11956__D _18093_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20227_ _12697_/A _15378_/A _20218_/A vssd1 vssd1 vccd1 vccd1 _20228_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__17924__C _17981_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20158_ _20158_/A _20158_/B _20158_/C vssd1 vssd1 vccd1 vccd1 _20167_/A sky130_fd_sc_hd__nand3_2
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17643__D _20745_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18101__B _18127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ _15774_/D vssd1 vssd1 vccd1 vccd1 _15577_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20089_ _20089_/A _20089_/B _20341_/C vssd1 vssd1 vccd1 vccd1 _20214_/A sky130_fd_sc_hd__nand3_2
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21746__D1 _22176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20013__A1 _18023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17414__C1 _17412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _11693_/X _11736_/Y _11762_/A _11932_/B vssd1 vssd1 vccd1 vccd1 _11931_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14650_/A _14740_/B _14650_/C vssd1 vssd1 vccd1 vccd1 _14650_/X sky130_fd_sc_hd__and3_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _16106_/C vssd1 vssd1 vccd1 vccd1 _12065_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19167__C1 _19461_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20359__A _20359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13601_ _13601_/A _13618_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _13602_/B sky130_fd_sc_hd__and3_1
XFILLER_14_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15460__B _15810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _13970_/X _14581_/B _14775_/C _14581_/D vssd1 vssd1 vccd1 vccd1 _14863_/B
+ sky130_fd_sc_hd__nand4b_4
XFILLER_72_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _11793_/A _11793_/B vssd1 vssd1 vccd1 vccd1 _11794_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16320_ _16320_/A _16320_/B vssd1 vssd1 vccd1 vccd1 _16579_/A sky130_fd_sc_hd__nor2_4
XFILLER_158_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13532_ _21362_/B vssd1 vssd1 vccd1 vccd1 _21805_/B sky130_fd_sc_hd__buf_2
XFILLER_9_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16251_ _16530_/C _16530_/B _16530_/D _16530_/A vssd1 vssd1 vccd1 vccd1 _16540_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_158_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13463_ _13461_/A _13461_/B _13563_/C vssd1 vssd1 vccd1 vccd1 _13463_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_256 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15743__A2 _15309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15202_ _15171_/A _15174_/A _15200_/X vssd1 vssd1 vccd1 vccd1 _15209_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__20806__B _20806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12414_ _12292_/A _15369_/B _12413_/X vssd1 vssd1 vccd1 vccd1 _20255_/C sky130_fd_sc_hd__a21oi_4
X_16182_ _16168_/Y _16171_/Y _16176_/Y _16181_/X vssd1 vssd1 vccd1 vccd1 _16183_/B
+ sky130_fd_sc_hd__a22oi_1
X_13394_ _13340_/Y _13341_/X _13352_/Y _13393_/Y vssd1 vssd1 vccd1 vccd1 _13394_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_138_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15133_ _15133_/A _15132_/Y vssd1 vssd1 vccd1 vccd1 _15134_/B sky130_fd_sc_hd__or2b_1
XANTENNA__15188__A _15188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12345_ _15320_/A vssd1 vssd1 vccd1 vccd1 _20086_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15619__C _18876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19941_ _19941_/A _19941_/B _19981_/A _19941_/D vssd1 vssd1 vccd1 vccd1 _19945_/A
+ sky130_fd_sc_hd__or4_1
X_15064_ _15114_/A _15114_/B _15064_/C _15118_/A vssd1 vssd1 vccd1 vccd1 _15065_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_107_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12276_ _12276_/A vssd1 vssd1 vccd1 vccd1 _12421_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14015_ _13857_/X _13725_/Y _13728_/A vssd1 vssd1 vccd1 vccd1 _14057_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__17248__A2 _16779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19872_ _19872_/A _19872_/B vssd1 vssd1 vccd1 vccd1 _19872_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__22865__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18823_ _18823_/A _18823_/B _18823_/C vssd1 vssd1 vccd1 vccd1 _18835_/C sky130_fd_sc_hd__nand3_1
XFILLER_1_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18754_ _18763_/B vssd1 vssd1 vccd1 vccd1 _18754_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15966_ _17643_/A _16192_/B _17039_/A _17401_/A vssd1 vssd1 vccd1 vccd1 _15966_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_49_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17705_ _17605_/B _17605_/A _17781_/C vssd1 vssd1 vccd1 vccd1 _17705_/Y sky130_fd_sc_hd__o21ai_1
X_14917_ _15107_/C _14917_/B _14917_/C vssd1 vssd1 vccd1 vccd1 _14917_/X sky130_fd_sc_hd__and3_1
XFILLER_64_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18685_ _18980_/A _19687_/A _18869_/A _18862_/A vssd1 vssd1 vccd1 vccd1 _18905_/A
+ sky130_fd_sc_hd__a22o_1
X_15897_ _15891_/A _15504_/X _15975_/A vssd1 vssd1 vccd1 vccd1 _15924_/A sky130_fd_sc_hd__o21ai_4
XFILLER_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17636_ _17636_/A vssd1 vssd1 vccd1 vccd1 _17876_/A sky130_fd_sc_hd__clkbuf_2
X_14848_ _14848_/A vssd1 vssd1 vccd1 vccd1 _22676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17567_ _17574_/C _17574_/B vssd1 vssd1 vccd1 vccd1 _17626_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14779_ _14779_/A _14857_/B _14858_/A _14859_/A vssd1 vssd1 vccd1 vccd1 _14895_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15982__A2 _15981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13171__A _22841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19306_ _11345_/X _11351_/X _19983_/B _19983_/A _18371_/X vssd1 vssd1 vccd1 vccd1
+ _19306_/X sky130_fd_sc_hd__o32a_1
X_16518_ _16508_/X _16510_/Y _16512_/Y _16517_/Y vssd1 vssd1 vccd1 vccd1 _16519_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_108_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ _17353_/X _17230_/Y _17375_/A _17513_/B vssd1 vssd1 vccd1 vccd1 _17726_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_182_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19237_ _19237_/A _19237_/B _19237_/C _19237_/D vssd1 vssd1 vccd1 vccd1 _19396_/C
+ sky130_fd_sc_hd__nand4_4
X_16449_ _16257_/Y _16816_/A _16452_/A vssd1 vssd1 vccd1 vccd1 _16451_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__16482__A _16482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19496__C _19496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19168_ _19318_/A _19461_/B _19168_/C vssd1 vssd1 vccd1 vccd1 _19168_/Y sky130_fd_sc_hd__nand3_4
X_18119_ _22795_/Q vssd1 vssd1 vccd1 vccd1 _18500_/C sky130_fd_sc_hd__inv_2
XANTENNA__19793__A _19793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19099_ _19106_/A _19106_/B _19097_/X _19098_/X vssd1 vssd1 vccd1 vccd1 _19117_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_172_451 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21130_ _21130_/A _21130_/B vssd1 vssd1 vccd1 vccd1 _21130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21061_ _21061_/A _21061_/B vssd1 vssd1 vccd1 vccd1 _21061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18202__A _18571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20012_ _20012_/A _20012_/B _20012_/C vssd1 vssd1 vccd1 vccd1 _20012_/X sky130_fd_sc_hd__and3_1
XFILLER_86_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20243__A1 _15326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18987__A2 _18984_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20794__A2 _16746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22659__A _22659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_980 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12484__A1 _20250_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21963_ _21963_/A vssd1 vssd1 vccd1 vccd1 _22220_/A sky130_fd_sc_hd__buf_2
XFILLER_39_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ _21019_/A _21019_/B _21083_/C vssd1 vssd1 vccd1 vccd1 _20919_/B sky130_fd_sc_hd__and3_1
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21894_ _21847_/A _21847_/B _21892_/Y _21893_/X vssd1 vssd1 vccd1 vccd1 _21933_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20845_ _21082_/B _15919_/X _20717_/B _20717_/A _20683_/B vssd1 vssd1 vccd1 vccd1
+ _20884_/A sky130_fd_sc_hd__o221a_1
XANTENNA__15973__A2 _16100_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19687__B _19687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20776_ _20776_/A _22935_/Q _20776_/C vssd1 vssd1 vccd1 vccd1 _20776_/X sky130_fd_sc_hd__and3_1
XFILLER_168_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18372__B1 _11821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_936 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22515_ _22571_/A vssd1 vssd1 vccd1 vccd1 _22584_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_50_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16922__A1 _15792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15725__A2 _15631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16922__B2 _16016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22446_ _22446_/A vssd1 vssd1 vccd1 vccd1 _22720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18640__B1_N _18933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22377_ _22377_/A vssd1 vssd1 vccd1 vccd1 _22690_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__22888__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ _12130_/A _18339_/C vssd1 vssd1 vccd1 vccd1 _12130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21328_ _21336_/B _13295_/X _13297_/A _14380_/A vssd1 vssd1 vccd1 vccd1 _21330_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_190_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17935__B _21082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1086 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21259_ _21689_/A _21259_/B _21259_/C vssd1 vssd1 vccd1 vccd1 _21260_/A sky130_fd_sc_hd__or3_1
X_12061_ _12061_/A _12061_/B _12061_/C vssd1 vssd1 vccd1 vccd1 _18238_/A sky130_fd_sc_hd__nand3_1
XFILLER_150_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18112__A _18278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12172__B1 _18716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20785__A2 _15940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15820_ _15727_/A _15727_/B _15817_/A vssd1 vssd1 vccd1 vccd1 _15826_/A sky130_fd_sc_hd__o21ai_2
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _15747_/Y _15756_/B _15750_/Y vssd1 vssd1 vccd1 vccd1 _15854_/B sky130_fd_sc_hd__a21oi_2
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21473__A _21473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12963_ _12963_/A _12963_/B _12997_/A _12963_/D vssd1 vssd1 vccd1 vccd1 _13004_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21734__A1 _21963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1032 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15471__A _19587_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14702_ _14366_/X _14863_/B _14869_/B _22765_/Q vssd1 vssd1 vccd1 vccd1 _14868_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18060__C1 _21081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17402__A2 _17400_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _18457_/Y _18462_/Y _18463_/X _18407_/B _18469_/Y vssd1 vssd1 vccd1 vccd1
+ _18765_/A sky130_fd_sc_hd__o221ai_4
X_11914_ _11914_/A _11914_/B vssd1 vssd1 vccd1 vccd1 _11914_/Y sky130_fd_sc_hd__nor2_1
X_15682_ _15682_/A vssd1 vssd1 vccd1 vccd1 _15682_/Y sky130_fd_sc_hd__inv_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12894_ _12894_/A _12894_/B vssd1 vssd1 vccd1 vccd1 _12894_/Y sky130_fd_sc_hd__nor2_4
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17421_/A vssd1 vssd1 vccd1 vccd1 _17421_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _14740_/A _14636_/B _14631_/Y _14632_/X vssd1 vssd1 vccd1 vccd1 _14650_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_11845_ _15792_/B vssd1 vssd1 vccd1 vccd1 _11845_/X sky130_fd_sc_hd__buf_4
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17352_ _17344_/Y _17347_/Y _17351_/Y vssd1 vssd1 vccd1 vccd1 _17352_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14564_ _14565_/A _14566_/A _14564_/C vssd1 vssd1 vccd1 vccd1 _14685_/A sky130_fd_sc_hd__nand3_2
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _19197_/A vssd1 vssd1 vccd1 vccd1 _19496_/C sky130_fd_sc_hd__clkbuf_4
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16293_/X _16294_/X _11627_/A _20605_/A vssd1 vssd1 vccd1 vccd1 _16552_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_186_543 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13515_ _13515_/A vssd1 vssd1 vccd1 vccd1 _13563_/A sky130_fd_sc_hd__clkbuf_2
X_17283_ _19615_/C _17449_/A _17293_/B _20917_/B vssd1 vssd1 vccd1 vccd1 _17285_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__15177__B1 _15180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14495_ _14500_/A _14611_/A _14500_/B _14500_/C vssd1 vssd1 vccd1 vccd1 _14611_/B
+ sky130_fd_sc_hd__nand4_1
X_19022_ _19022_/A _19022_/B _19022_/C vssd1 vssd1 vccd1 vccd1 _19029_/A sky130_fd_sc_hd__nand3_1
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ _12719_/A _17137_/A _16506_/A vssd1 vssd1 vccd1 vccd1 _16234_/X sky130_fd_sc_hd__o21a_1
X_13446_ _13465_/B vssd1 vssd1 vccd1 vccd1 _13446_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16165_ _16166_/A _16166_/B _16166_/C vssd1 vssd1 vccd1 vccd1 _16165_/Y sky130_fd_sc_hd__a21oi_1
X_13377_ _13579_/A _21522_/A _21522_/C _21177_/D vssd1 vssd1 vccd1 vccd1 _13377_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_138_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15116_ _15188_/B _15185_/B _15115_/Y vssd1 vssd1 vccd1 vccd1 _15119_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__20473__A1 _12734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12328_ _12577_/A _12576_/A _12348_/A _12418_/A vssd1 vssd1 vccd1 vccd1 _12329_/A
+ sky130_fd_sc_hd__o211ai_1
X_16096_ _16044_/Y _16041_/X _16201_/B vssd1 vssd1 vccd1 vccd1 _16096_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14152__A1 _14165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19924_ _19921_/Y _19872_/Y _19922_/X _19923_/Y vssd1 vssd1 vccd1 vccd1 _19962_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_170_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15047_ _15039_/A _15047_/B _15047_/C vssd1 vssd1 vccd1 vccd1 _15098_/B sky130_fd_sc_hd__nand3b_1
X_12259_ _18266_/A _12259_/B vssd1 vssd1 vccd1 vccd1 _12260_/A sky130_fd_sc_hd__or2_1
XANTENNA__14550__A _14863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19855_ _19852_/Y _19853_/Y _19793_/A _19795_/X vssd1 vssd1 vccd1 vccd1 _19913_/A
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__15365__B _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17283__D _20917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18806_ _18795_/X _16799_/X _18804_/A vssd1 vssd1 vccd1 vccd1 _18824_/A sky130_fd_sc_hd__o21ai_1
X_19786_ _19782_/A _19782_/B _19784_/C _19784_/A vssd1 vssd1 vccd1 vccd1 _19788_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__14455__A2 _15435_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16998_ _16998_/A vssd1 vssd1 vccd1 vccd1 _17081_/A sky130_fd_sc_hd__buf_2
XFILLER_3_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21383__A _21383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18737_ _18743_/B vssd1 vssd1 vccd1 vccd1 _18737_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15949_ _15949_/A _15949_/B vssd1 vssd1 vccd1 vccd1 _16035_/C sky130_fd_sc_hd__nand2_2
XFILLER_97_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15812__C _15812_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18668_ _11979_/Y _11980_/X _16276_/X _15580_/X _11639_/X vssd1 vssd1 vccd1 vccd1
+ _18668_/X sky130_fd_sc_hd__o32a_1
XANTENNA__15404__A1 _12606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16601__B1 _16600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17619_ _17720_/A _17619_/B vssd1 vssd1 vccd1 vccd1 _22959_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__12218__A1 _18830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15955__A2 _17816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18599_ _12258_/A _18251_/Y _18598_/Y _18601_/A _18601_/B vssd1 vssd1 vccd1 vccd1
+ _18599_/X sky130_fd_sc_hd__a32o_1
XFILLER_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14612__C1 _13823_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20630_ _20630_/A _20634_/B _20634_/C vssd1 vssd1 vccd1 vccd1 _20631_/C sky130_fd_sc_hd__nand3_1
XFILLER_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20561_ _20560_/Y _20315_/Y _20313_/A vssd1 vssd1 vccd1 vccd1 _20562_/B sky130_fd_sc_hd__o21ai_1
XFILLER_192_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22300_ _22300_/A _22300_/B vssd1 vssd1 vccd1 vccd1 _22341_/A sky130_fd_sc_hd__nor2_1
X_20492_ _20458_/Y _20353_/A _20366_/A _20366_/B vssd1 vssd1 vccd1 vccd1 _20500_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22231_ _22265_/C _22231_/B _22231_/C _22231_/D vssd1 vssd1 vccd1 vccd1 _22232_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_117_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15259__C _15259_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22162_ _22158_/Y _21836_/A _22161_/X vssd1 vssd1 vccd1 vccd1 _22162_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_117_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21113_ _21107_/Y _21108_/Y _21138_/C vssd1 vssd1 vccd1 vccd1 _21135_/A sky130_fd_sc_hd__o21bai_2
X_22093_ _22092_/A _22092_/B _22680_/Q vssd1 vssd1 vccd1 vccd1 _22094_/B sky130_fd_sc_hd__a21oi_1
XFILLER_182_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13351__C1 _21767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21044_ _21082_/B _21044_/B _21044_/C vssd1 vssd1 vccd1 vccd1 _21044_/X sky130_fd_sc_hd__or3_1
XFILLER_119_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19970__B _22923_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17093__B1 _17085_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13076__A _13304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11308__B _11308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21946_ _22037_/B _22122_/C _22037_/A vssd1 vssd1 vccd1 vccd1 _21946_/Y sky130_fd_sc_hd__nand3_1
XFILLER_55_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17396__A1 _15934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21877_ _21877_/A vssd1 vssd1 vccd1 vccd1 _22221_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11630_ _11647_/C _11647_/D vssd1 vssd1 vccd1 vccd1 _11630_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20828_ _20828_/A vssd1 vssd1 vccd1 vccd1 _20994_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20637__A _20637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11561_ _11568_/A vssd1 vssd1 vccd1 vccd1 _11561_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__20152__B1 _20125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20759_ _20759_/A _20759_/B vssd1 vssd1 vccd1 vccd1 _20891_/A sky130_fd_sc_hd__nand2_1
XFILLER_196_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17649__C _18303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18107__A _18107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ _13300_/A _13300_/B vssd1 vssd1 vccd1 vccd1 _13300_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14280_ _14280_/A _14280_/B _14280_/C vssd1 vssd1 vccd1 vccd1 _14281_/C sky130_fd_sc_hd__nand3_1
XFILLER_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11492_ _18682_/C vssd1 vssd1 vccd1 vccd1 _16078_/C sky130_fd_sc_hd__buf_4
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13231_ _13234_/B _13157_/A _13230_/X vssd1 vssd1 vccd1 vccd1 _13504_/B sky130_fd_sc_hd__a21oi_2
XFILLER_136_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22429_ _22714_/Q input53/X _22435_/S vssd1 vssd1 vccd1 vccd1 _22430_/A sky130_fd_sc_hd__mux2_1
XANTENNA__19845__B1 _19900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input65_A wb_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ _13162_/A _13504_/A _13162_/C vssd1 vssd1 vccd1 vccd1 _13384_/A sky130_fd_sc_hd__or3_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12113_ _16274_/A vssd1 vssd1 vccd1 vccd1 _16921_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14134__A1 _13736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11994__A _12107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15466__A _15557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17970_ _22903_/Q _17970_/B vssd1 vssd1 vccd1 vccd1 _17970_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14370__A _14370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ _21214_/A _21213_/A vssd1 vssd1 vccd1 vccd1 _13125_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17608__C1 _17502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19073__A1 _11625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12044_ _16477_/B vssd1 vssd1 vccd1 vccd1 _19197_/D sky130_fd_sc_hd__buf_2
X_16921_ _16921_/A vssd1 vssd1 vccd1 vccd1 _16921_/X sky130_fd_sc_hd__buf_2
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18777__A _19941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19640_ _19635_/Y _19638_/Y _19649_/B vssd1 vssd1 vccd1 vccd1 _19640_/X sky130_fd_sc_hd__a21o_1
XFILLER_172_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18281__C1 _19358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16852_ _16848_/X _16853_/B _16853_/C vssd1 vssd1 vccd1 vccd1 _16852_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_120_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15634__A1 _18512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15803_ _15803_/A vssd1 vssd1 vccd1 vccd1 _15803_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22903__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19571_ _19571_/A _19571_/B _22918_/Q vssd1 vssd1 vccd1 vccd1 _19574_/B sky130_fd_sc_hd__nand3_2
XFILLER_168_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16783_ _16515_/Y _16941_/A _16781_/Y _16782_/X vssd1 vssd1 vccd1 vccd1 _16792_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_19_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13995_ _13877_/Y _14686_/B _14808_/A _13881_/Y vssd1 vssd1 vccd1 vccd1 _13998_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_93_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18522_ _18915_/A _18916_/A vssd1 vssd1 vccd1 vccd1 _18522_/Y sky130_fd_sc_hd__nand2_1
X_15734_ _15752_/A _15752_/B _15752_/C _15825_/A _15825_/C vssd1 vssd1 vccd1 vccd1
+ _15734_/X sky130_fd_sc_hd__a32o_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12946_ _20249_/C _20584_/C _12950_/C _12950_/B vssd1 vssd1 vccd1 vccd1 _12954_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22380__A1 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18453_ _19199_/B _19199_/C _18453_/C vssd1 vssd1 vccd1 vccd1 _18453_/X sky130_fd_sc_hd__and3_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _15665_/A _15665_/B _15665_/C vssd1 vssd1 vccd1 vccd1 _15668_/A sky130_fd_sc_hd__and3_1
XANTENNA__15937__A2 _15792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20391__B1 _20263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ _22827_/Q vssd1 vssd1 vccd1 vccd1 _20870_/C sky130_fd_sc_hd__buf_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_655 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19128__A2 _18812_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _15903_/X _20255_/A _17647_/A _18814_/A _16177_/A vssd1 vssd1 vccd1 vccd1
+ _17404_/X sky130_fd_sc_hd__o32a_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _14727_/A _14721_/B _15005_/B _15006_/B vssd1 vssd1 vccd1 vccd1 _14616_/Y
+ sky130_fd_sc_hd__nand4_1
X_18384_ _18165_/A _18165_/B _18383_/Y _18310_/Y vssd1 vssd1 vccd1 vccd1 _18384_/Y
+ sky130_fd_sc_hd__a22oi_1
X_11828_ _11817_/Y _11822_/X _11811_/Y _11815_/Y vssd1 vssd1 vccd1 vccd1 _11829_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_61_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15596_ _15596_/A vssd1 vssd1 vccd1 vccd1 _15596_/Y sky130_fd_sc_hd__inv_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17335_ _17335_/A _17486_/C vssd1 vssd1 vccd1 vccd1 _17335_/Y sky130_fd_sc_hd__nand2_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14547_ _14547_/A _14547_/B _14547_/C vssd1 vssd1 vccd1 vccd1 _14661_/B sky130_fd_sc_hd__nand3_1
XFILLER_159_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11759_ _11703_/X _11752_/Y _11755_/Y _11758_/Y vssd1 vssd1 vccd1 vccd1 _11762_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17266_ _17299_/A _17299_/C vssd1 vssd1 vccd1 vccd1 _17266_/Y sky130_fd_sc_hd__nand2_1
X_14478_ _14478_/A _14478_/B _14478_/C vssd1 vssd1 vccd1 vccd1 _14611_/A sky130_fd_sc_hd__nand3_4
XANTENNA__16362__A2 _15645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16217_ _16217_/A vssd1 vssd1 vccd1 vccd1 _18192_/A sky130_fd_sc_hd__buf_2
X_19005_ _18891_/X _18893_/X _19085_/A vssd1 vssd1 vccd1 vccd1 _19009_/B sky130_fd_sc_hd__o21ai_1
XFILLER_174_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14373__A1 _18698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13429_ _13579_/A vssd1 vssd1 vccd1 vccd1 _13635_/A sky130_fd_sc_hd__clkbuf_2
X_17197_ _17197_/A _17197_/B _17197_/C vssd1 vssd1 vccd1 vccd1 _17197_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__18639__B2 _18546_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12065__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14373__B2 _22765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16148_ _16131_/A _16131_/B _16146_/Y _16147_/Y vssd1 vssd1 vccd1 vccd1 _16148_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_6_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12923__A2 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22912__D _22912_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15376__A _15382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16079_ _16080_/A _16080_/C _16080_/B vssd1 vssd1 vccd1 vccd1 _16081_/A sky130_fd_sc_hd__a21oi_1
XFILLER_170_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19907_ _19907_/A _19907_/B vssd1 vssd1 vccd1 vccd1 _19907_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19603__A3 _18131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11409__A _11712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19838_ _19838_/A vssd1 vssd1 vccd1 vccd1 _19987_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18811__A1 _12064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14428__A2 _14418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15823__B _16106_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 wb_adr_i[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
X_19769_ _19836_/A _19769_/B _19836_/C _19836_/D vssd1 vssd1 vccd1 vccd1 _19782_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_83_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13100__A2 _14380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21800_ _21671_/Y _21664_/X _21657_/Y _21648_/X vssd1 vssd1 vccd1 vccd1 _21803_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_22780_ _22812_/CLK _22780_/D vssd1 vssd1 vccd1 vccd1 _22780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14439__B _22967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_622 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21731_ _21730_/A _21730_/B _21730_/C _21730_/D vssd1 vssd1 vccd1 vccd1 _21777_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21841__A _21841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16935__A _19587_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16050__A1 _16613_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21560__B _21560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21662_ _21662_/A _21662_/B vssd1 vssd1 vccd1 vccd1 _21662_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20613_ _20613_/A _20613_/B _20613_/C vssd1 vssd1 vccd1 vccd1 _20620_/B sky130_fd_sc_hd__nand3_2
X_21593_ _21478_/X _21486_/A _21481_/B _21482_/Y vssd1 vssd1 vccd1 vccd1 _21771_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_131_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_bq_clk_i clkbuf_3_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_20544_ _20429_/C _20414_/X _20426_/X _20427_/Y vssd1 vssd1 vccd1 vccd1 _20544_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_192_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14364__A1 _16322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16670__A _16670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20475_ _20599_/A _20599_/B _20475_/C vssd1 vssd1 vccd1 vccd1 _20499_/D sky130_fd_sc_hd__nand3_1
XFILLER_69_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22214_ _22215_/A _22215_/B vssd1 vssd1 vccd1 vccd1 _22216_/A sky130_fd_sc_hd__nor2_1
XANTENNA__21634__B1 _21963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19981__A _19981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22145_ _22145_/A _22145_/B _22145_/C vssd1 vssd1 vccd1 vccd1 _22146_/A sky130_fd_sc_hd__nand3_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14667__A2 _14843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19055__A1 _18330_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13518__B _13521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22076_ _22073_/Y _22074_/Y _22075_/X vssd1 vssd1 vccd1 vccd1 _22163_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__22611__S _22619_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22926__CLK _22948_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11319__A _18107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21027_ _21027_/A _21027_/B vssd1 vssd1 vccd1 vccd1 _21030_/C sky130_fd_sc_hd__and2_1
XANTENNA__19460__D1 _19614_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12800_ _12792_/Y _12796_/Y _12799_/X vssd1 vssd1 vccd1 vccd1 _12863_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_663 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13780_ _14613_/A vssd1 vssd1 vccd1 vccd1 _15008_/C sky130_fd_sc_hd__buf_2
XANTENNA__11980__C _11980_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15452__C _16772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12731_ _12916_/A _12916_/B _12917_/A vssd1 vssd1 vccd1 vccd1 _12739_/A sky130_fd_sc_hd__o21ai_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21929_ _21929_/A _21929_/B vssd1 vssd1 vccd1 vccd1 _22935_/D sky130_fd_sc_hd__nor2_1
XFILLER_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16041__A1 _15936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20912__A2 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15450_ _15450_/A vssd1 vssd1 vccd1 vccd1 _15450_/X sky130_fd_sc_hd__buf_4
XANTENNA__14068__C _14868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12662_ _12913_/A vssd1 vssd1 vccd1 vccd1 _15746_/B sky130_fd_sc_hd__buf_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16592__A2 _16745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16564__B _16564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14401_ _22805_/Q _14397_/X _14398_/X _14391_/X _22773_/Q vssd1 vssd1 vccd1 vccd1
+ _14401_/X sky130_fd_sc_hd__a32o_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11989__A _15776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11613_ _12094_/D vssd1 vssd1 vccd1 vccd1 _15774_/B sky130_fd_sc_hd__buf_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18482__D _19168_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15381_ _20593_/B vssd1 vssd1 vccd1 vccd1 _17530_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_338 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12593_ _12588_/Y _20471_/C _16477_/C _12592_/Y vssd1 vssd1 vccd1 vccd1 _12601_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _17120_/A _17120_/B vssd1 vssd1 vccd1 vccd1 _17122_/B sky130_fd_sc_hd__nand2_2
XANTENNA__20086__B _20323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_822 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14332_ _11860_/C _14317_/X _14320_/X _14331_/X _12493_/A vssd1 vssd1 vccd1 vccd1
+ _14332_/X sky130_fd_sc_hd__a32o_1
X_11544_ _15624_/A vssd1 vssd1 vccd1 vccd1 _16106_/C sky130_fd_sc_hd__buf_4
XANTENNA__21873__B1 _22057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_343 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17051_ _16433_/C _16439_/Y _17076_/B _16440_/Y vssd1 vssd1 vccd1 vccd1 _17053_/A
+ sky130_fd_sc_hd__o211ai_1
X_14263_ _14512_/A _14269_/A _14263_/C _14276_/D vssd1 vssd1 vccd1 vccd1 _14279_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11475_ _11818_/A _17083_/A _11468_/Y _11474_/X _11565_/A vssd1 vssd1 vccd1 vccd1
+ _11894_/B sky130_fd_sc_hd__o221ai_4
XFILLER_109_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16002_ _16010_/A _16010_/B _16011_/A _16011_/B vssd1 vssd1 vccd1 vccd1 _16003_/C
+ sky130_fd_sc_hd__nand4_1
X_13214_ _13210_/A _13210_/B _13350_/A _13213_/X vssd1 vssd1 vccd1 vccd1 _13215_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_7_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1096 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14194_ _14230_/A vssd1 vssd1 vccd1 vccd1 _14953_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_1112 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21629__C _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _13145_/A vssd1 vssd1 vccd1 vccd1 _13157_/A sky130_fd_sc_hd__buf_2
XFILLER_152_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1099 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _17953_/A _17953_/B vssd1 vssd1 vccd1 vccd1 _18002_/C sky130_fd_sc_hd__nand2_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _13304_/B vssd1 vssd1 vccd1 vccd1 _13079_/A sky130_fd_sc_hd__inv_2
XFILLER_105_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16904_ _16899_/Y _17070_/A _16903_/X vssd1 vssd1 vccd1 vccd1 _16905_/B sky130_fd_sc_hd__a21boi_1
X_12027_ _12054_/A _12054_/B _12055_/A _12055_/B vssd1 vssd1 vccd1 vccd1 _12027_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11877__C1 _18259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17884_ _17883_/D _17883_/B _17929_/A _20975_/B vssd1 vssd1 vccd1 vccd1 _17885_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19623_ _19615_/X _19616_/X _19621_/Y _19622_/X vssd1 vssd1 vccd1 vccd1 _19709_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16835_ _17436_/A vssd1 vssd1 vccd1 vccd1 _19615_/C sky130_fd_sc_hd__buf_2
XFILLER_54_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19554_ _19551_/Y _19552_/Y _19553_/X vssd1 vssd1 vccd1 vccd1 _19555_/D sky130_fd_sc_hd__o21bai_1
X_16766_ _16766_/A vssd1 vssd1 vccd1 vccd1 _16954_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13094__A1 _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13978_ _13978_/A vssd1 vssd1 vccd1 vccd1 _14191_/A sky130_fd_sc_hd__buf_2
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18505_ _18319_/A _18500_/Y _18319_/C _18698_/A vssd1 vssd1 vccd1 vccd1 _18876_/B
+ sky130_fd_sc_hd__o211ai_4
X_15717_ _17128_/B _16720_/C _15403_/X _15423_/Y vssd1 vssd1 vccd1 vccd1 _15752_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12929_ _12929_/A vssd1 vssd1 vccd1 vccd1 _12930_/A sky130_fd_sc_hd__clkbuf_4
X_19485_ _19342_/A _19342_/B _19342_/C _19340_/A vssd1 vssd1 vccd1 vccd1 _19486_/B
+ sky130_fd_sc_hd__a31oi_4
X_16697_ _16697_/A _16697_/B vssd1 vssd1 vccd1 vccd1 _16698_/C sky130_fd_sc_hd__nand2_1
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12841__A1 _20255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12841__B2 _16300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16032__A1 _15966_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18436_ _18601_/A _18601_/B _18430_/A vssd1 vssd1 vccd1 vccd1 _18960_/B sky130_fd_sc_hd__a21oi_2
X_15648_ _15918_/A _16737_/A _15645_/X _15646_/X _16400_/A vssd1 vssd1 vccd1 vccd1
+ _15648_/X sky130_fd_sc_hd__o221a_1
XFILLER_34_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19506__C1 _17532_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11899__A _11899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15579_ _15465_/X _15466_/Y _15546_/A _16921_/A vssd1 vssd1 vccd1 vccd1 _15579_/X
+ sky130_fd_sc_hd__o22a_1
X_18367_ _18367_/A _18367_/B _18367_/C _18659_/D vssd1 vssd1 vccd1 vccd1 _18367_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_175_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17318_ _17318_/A _17318_/B vssd1 vssd1 vccd1 vccd1 _17320_/A sky130_fd_sc_hd__nand2_1
X_18298_ _17822_/A _18778_/A _18305_/D _18305_/A vssd1 vssd1 vccd1 vccd1 _18301_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14346__A1 _12320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17249_ _12696_/X _17403_/A _17142_/A vssd1 vssd1 vccd1 vccd1 _17249_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_147_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21616__B1 _21944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20260_ _20260_/A vssd1 vssd1 vccd1 vccd1 _20260_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19285__A1 _19443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16099__A1 _13022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16099__B2 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20191_ _20191_/A _20191_/B vssd1 vssd1 vccd1 vccd1 _20192_/B sky130_fd_sc_hd__xor2_2
XFILLER_89_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18848__C _18848_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15834__A _15834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_563 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22901_ _22951_/CLK _22901_/D vssd1 vssd1 vccd1 vccd1 _22901_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__17680__B1_N _17669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15553__B _19358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19025__B _19496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16271__A1 _15580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22832_ _22850_/CLK _22844_/Q vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_622 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22763_ _22807_/CLK _22763_/D vssd1 vssd1 vccd1 vccd1 _22763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21714_ _21714_/A vssd1 vssd1 vccd1 vccd1 _21801_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22694_ _22696_/CLK _22694_/D vssd1 vssd1 vccd1 vccd1 _22694_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21645_ _21645_/A _21645_/B _21645_/C _21645_/D vssd1 vssd1 vccd1 vccd1 _21645_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_75_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21576_ _21576_/A _21576_/B vssd1 vssd1 vccd1 vccd1 _21917_/B sky130_fd_sc_hd__nand2_2
XFILLER_123_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20527_ _20532_/A _20532_/B _20529_/A _20534_/A vssd1 vssd1 vccd1 vccd1 _20531_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15728__B _16781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20458_ _20456_/Y _20339_/Y _20347_/B _20457_/Y _20221_/Y vssd1 vssd1 vccd1 vccd1
+ _20458_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_180_346 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17287__B1 _17286_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20389_ _20378_/Y _20381_/Y _20388_/Y vssd1 vssd1 vccd1 vccd1 _20396_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__15298__C1 _18093_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16495__D1 _19507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19028__A1 _19012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22128_ _22128_/A _22219_/A _22128_/C vssd1 vssd1 vccd1 vccd1 _22170_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19216__A _19507_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14950_ _15061_/A _14013_/A _14013_/B _15002_/A _14951_/C vssd1 vssd1 vccd1 vccd1
+ _14952_/A sky130_fd_sc_hd__a32o_1
XFILLER_43_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1072 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22059_ _22122_/C _22262_/A _22223_/A _22062_/A vssd1 vssd1 vccd1 vccd1 _22059_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13901_ _13793_/Y _13745_/C _13833_/C vssd1 vssd1 vccd1 vccd1 _13902_/B sky130_fd_sc_hd__a21o_1
XFILLER_43_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input28_A wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881_ _14881_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14887_/C sky130_fd_sc_hd__nor2_1
XFILLER_130_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16620_ _16620_/A _16620_/B _16620_/C vssd1 vssd1 vccd1 vccd1 _16637_/A sky130_fd_sc_hd__nand3_2
XANTENNA__16262__B2 _15723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ _13737_/X _13746_/X _14074_/A vssd1 vssd1 vccd1 vccd1 _13837_/A sky130_fd_sc_hd__a21o_1
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14079__B _14489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16551_ _18680_/D _20092_/A _20092_/B vssd1 vssd1 vccd1 vccd1 _16714_/A sky130_fd_sc_hd__nand3_1
XFILLER_44_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13763_ _13763_/A vssd1 vssd1 vccd1 vccd1 _14203_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16575__A _20579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _15502_/A _15502_/B _15502_/C _15502_/D vssd1 vssd1 vccd1 vccd1 _15597_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_43_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12714_ _12522_/A _12522_/B _12928_/A vssd1 vssd1 vccd1 vccd1 _12714_/Y sky130_fd_sc_hd__a21oi_1
X_19270_ _19296_/A _19434_/A _19434_/B vssd1 vssd1 vccd1 vccd1 _19299_/B sky130_fd_sc_hd__nand3_1
X_16482_ _16482_/A _22967_/Q vssd1 vssd1 vccd1 vccd1 _16483_/B sky130_fd_sc_hd__and2_2
X_13694_ _14222_/A vssd1 vssd1 vccd1 vccd1 _14212_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15433_ _15433_/A _15682_/A vssd1 vssd1 vccd1 vccd1 _15859_/A sky130_fd_sc_hd__nand2_1
X_18221_ _18182_/A _18276_/B _18276_/A vssd1 vssd1 vccd1 vccd1 _18221_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12645_ _12645_/A _12769_/A _12645_/C vssd1 vssd1 vccd1 vccd1 _12645_/X sky130_fd_sc_hd__and3_1
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18152_ _18389_/A _18389_/B _18389_/C vssd1 vssd1 vccd1 vccd1 _18383_/B sky130_fd_sc_hd__nand3_2
XFILLER_8_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15364_ _20341_/B vssd1 vssd1 vccd1 vccd1 _20101_/B sky130_fd_sc_hd__buf_2
XANTENNA__12051__A2 _11762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16317__A2 _15905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12576_ _12576_/A vssd1 vssd1 vccd1 vccd1 _12576_/X sky130_fd_sc_hd__buf_4
XFILLER_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17103_ _17103_/A _17338_/B _17103_/C vssd1 vssd1 vccd1 vccd1 _17196_/B sky130_fd_sc_hd__nand3_1
X_14315_ _22514_/A _22514_/B vssd1 vssd1 vccd1 vccd1 _14411_/A sky130_fd_sc_hd__nor2_1
XANTENNA__14328__A1 _12470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18083_ _18082_/B _18082_/C _22908_/Q vssd1 vssd1 vccd1 vccd1 _18084_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__15919__A _15919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15525__B1 _16759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11527_ _11378_/X _11299_/X _11420_/C _11471_/C vssd1 vssd1 vccd1 vccd1 _12003_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_157_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15295_ _22884_/Q _22885_/Q _22886_/Q _15288_/A _22888_/Q vssd1 vssd1 vccd1 vccd1
+ _15296_/B sky130_fd_sc_hd__o41a_1
XFILLER_116_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17034_ _16853_/C _16848_/X _16740_/Y _16733_/Y vssd1 vssd1 vccd1 vccd1 _17036_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14246_ _14246_/A _14246_/B vssd1 vssd1 vccd1 vccd1 _14253_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11458_ _11324_/X _11675_/B _14429_/A vssd1 vssd1 vccd1 vccd1 _11505_/A sky130_fd_sc_hd__a21oi_2
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14177_ _14094_/B _14094_/C _14094_/A vssd1 vssd1 vccd1 vccd1 _14178_/A sky130_fd_sc_hd__a21o_1
XANTENNA__15357__C _16304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11389_ _18482_/A vssd1 vssd1 vccd1 vccd1 _18984_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12343__A _12378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19019__A1 _17421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ _21220_/A _13319_/A _13126_/X _21606_/A vssd1 vssd1 vccd1 vccd1 _13128_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_3_0_bq_clk_i_A clkbuf_2_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _19480_/A _19481_/A _18985_/C vssd1 vssd1 vccd1 vccd1 _18985_/Y sky130_fd_sc_hd__nand3_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _17935_/C _17974_/A _17872_/C _17840_/A vssd1 vssd1 vccd1 vccd1 _17991_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _22727_/Q vssd1 vssd1 vccd1 vccd1 _13095_/A sky130_fd_sc_hd__buf_2
XFILLER_87_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater126 _22888_/Q vssd1 vssd1 vccd1 vccd1 _22876_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater137 _22789_/CLK vssd1 vssd1 vccd1 vccd1 _22787_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17867_ _17866_/A _18007_/A _18007_/B vssd1 vssd1 vccd1 vccd1 _17868_/B sky130_fd_sc_hd__o21a_1
Xrepeater148 _22808_/CLK vssd1 vssd1 vccd1 vccd1 _22810_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater159 _22751_/CLK vssd1 vssd1 vccd1 vccd1 _22742_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15804__D _16067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_706 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19606_ _19317_/Y _19330_/B _19479_/C _19475_/Y vssd1 vssd1 vccd1 vccd1 _19610_/A
+ sky130_fd_sc_hd__a31o_1
X_16818_ _20608_/C vssd1 vssd1 vccd1 vccd1 _20928_/B sky130_fd_sc_hd__buf_2
X_17798_ _17705_/Y _17623_/Y _17607_/A _17708_/Y vssd1 vssd1 vccd1 vccd1 _17800_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19537_ _19538_/A _19538_/B _19538_/C vssd1 vssd1 vccd1 vccd1 _19537_/Y sky130_fd_sc_hd__a21oi_1
X_16749_ _16741_/Y _16749_/B _16749_/C vssd1 vssd1 vccd1 vccd1 _16853_/A sky130_fd_sc_hd__nand3b_4
XFILLER_35_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19468_ _17427_/X _19839_/D _19466_/Y _19467_/Y vssd1 vssd1 vccd1 vccd1 _19476_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__16556__A2 _17111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18419_ _18232_/X _18275_/X _18417_/Y _18418_/Y vssd1 vssd1 vccd1 vccd1 _18773_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_50_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19399_ _19399_/A _19399_/B _19399_/C vssd1 vssd1 vccd1 vccd1 _19408_/A sky130_fd_sc_hd__nand3_1
XFILLER_107_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21430_ _21430_/A _21565_/B vssd1 vssd1 vccd1 vccd1 _21431_/B sky130_fd_sc_hd__nand2_1
XFILLER_194_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21361_ _21183_/X _21212_/Y _21237_/A vssd1 vssd1 vccd1 vccd1 _21369_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__12593__A3 _16477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20312_ _20311_/B _20311_/C _20311_/A vssd1 vssd1 vccd1 vccd1 _20562_/A sky130_fd_sc_hd__a21o_1
Xinput70 x[10] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21292_ _21292_/A _22673_/Q _21292_/C vssd1 vssd1 vccd1 vccd1 _21294_/D sky130_fd_sc_hd__and3_1
XFILLER_116_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18466__C1 _17525_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20243_ _15326_/X _15325_/X _20128_/A _16257_/C vssd1 vssd1 vccd1 vccd1 _20244_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_66_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18859__B _19481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20174_ _20174_/A _20174_/B _20174_/C vssd1 vssd1 vccd1 vccd1 _20314_/C sky130_fd_sc_hd__nand3_4
XANTENNA__17284__A3 _17833_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12403__D _12403_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18769__B1 _18770_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15714__D _16772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12700__B _20579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17441__B1 _17880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__A _22842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22815_ _22815_/CLK _22815_/D vssd1 vssd1 vccd1 vccd1 _22815_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16395__A _20917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17339__A4 _17341_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22746_ _22746_/CLK _22746_/D vssd1 vssd1 vccd1 vccd1 _22746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19202__C _19504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22677_ _22944_/CLK _22677_/D vssd1 vssd1 vccd1 vccd1 _22677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12428__A _20359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12569__B1 _15363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12430_ _12334_/X _12350_/Y _12428_/Y vssd1 vssd1 vccd1 vccd1 _12430_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21628_ _21724_/A _21724_/C _21724_/D vssd1 vssd1 vccd1 vccd1 _21633_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12033__A2 _11736_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16842__B _16842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12361_ _12361_/A vssd1 vssd1 vccd1 vccd1 _12403_/D sky130_fd_sc_hd__clkinv_2
XFILLER_194_983 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21559_ _21559_/A _21559_/B vssd1 vssd1 vccd1 vccd1 _21561_/A sky130_fd_sc_hd__nand2_1
XFILLER_139_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18115__A _18115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14100_ _14032_/A _14039_/A _14099_/A vssd1 vssd1 vccd1 vccd1 _14100_/X sky130_fd_sc_hd__a21o_1
X_11312_ _22968_/Q vssd1 vssd1 vccd1 vccd1 _11713_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_165_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15080_ _15080_/A _15080_/B _15080_/C vssd1 vssd1 vccd1 vccd1 _15080_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__16180__B1 _15932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12292_ _12292_/A _12303_/A vssd1 vssd1 vccd1 vccd1 _16267_/A sky130_fd_sc_hd__nand2_2
XFILLER_181_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14031_ _14052_/A _14031_/B _14031_/C _14036_/B vssd1 vssd1 vccd1 vccd1 _14032_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_141_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13533__A2 _21805_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18770_ _18770_/A _18779_/B _18770_/C vssd1 vssd1 vccd1 vccd1 _18770_/X sky130_fd_sc_hd__and3_1
XANTENNA__21195__B _21195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15982_ _12968_/B _15981_/X _15901_/Y vssd1 vssd1 vccd1 vccd1 _16005_/A sky130_fd_sc_hd__o21ai_4
XFILLER_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15691__C1 _15690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17721_ _17721_/A _22900_/Q _17721_/C vssd1 vssd1 vccd1 vccd1 _17722_/B sky130_fd_sc_hd__nand3_1
XFILLER_121_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14933_ _14933_/A vssd1 vssd1 vccd1 vccd1 _15154_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17432__B1 _17238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17652_ _19585_/D _17652_/B vssd1 vssd1 vccd1 vccd1 _17652_/Y sky130_fd_sc_hd__nand2_2
X_14864_ _14571_/X _14583_/Y _14366_/X vssd1 vssd1 vccd1 vccd1 _14865_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__17983__A1 _21017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _16873_/A _16617_/C _16600_/X vssd1 vssd1 vccd1 vccd1 _16603_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15921__B _16157_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13815_ _22757_/Q vssd1 vssd1 vccd1 vccd1 _13815_/X sky130_fd_sc_hd__buf_2
X_17583_ _17580_/Y _17581_/Y _17582_/X _17524_/Y vssd1 vssd1 vccd1 vccd1 _17583_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15994__B1 _15649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14795_ _14685_/A _14685_/B _14695_/A vssd1 vssd1 vccd1 vccd1 _14884_/A sky130_fd_sc_hd__o21ai_2
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14818__A _14818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19322_ _19322_/A _19322_/B _19322_/C vssd1 vssd1 vccd1 vccd1 _19323_/A sky130_fd_sc_hd__nand3_1
XANTENNA__13722__A _22869_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16534_ _16534_/A _16534_/B vssd1 vssd1 vccd1 vccd1 _16536_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13746_ _13750_/B vssd1 vssd1 vccd1 vccd1 _13746_/X sky130_fd_sc_hd__buf_2
XFILLER_31_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19253_ _19148_/X _19150_/Y _19250_/Y _19252_/X vssd1 vssd1 vccd1 vccd1 _19253_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_92_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16465_ _16465_/A vssd1 vssd1 vccd1 vccd1 _20255_/A sky130_fd_sc_hd__clkbuf_4
X_13677_ _13677_/A _13677_/B _13677_/C vssd1 vssd1 vccd1 vccd1 _13678_/C sky130_fd_sc_hd__nand3_1
XFILLER_189_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18204_ _18204_/A vssd1 vssd1 vccd1 vccd1 _18402_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15416_ _15932_/A _15919_/A _15350_/Y _15415_/X vssd1 vssd1 vccd1 vccd1 _15703_/A
+ sky130_fd_sc_hd__o31a_1
X_12628_ _12628_/A _12628_/B vssd1 vssd1 vccd1 vccd1 _12630_/C sky130_fd_sc_hd__nand2_1
X_19184_ _19163_/X _19162_/Y _19155_/Y vssd1 vssd1 vccd1 vccd1 _19185_/B sky130_fd_sc_hd__o21ai_1
X_16396_ _20975_/B vssd1 vssd1 vccd1 vccd1 _21050_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_31_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18135_ _18135_/A vssd1 vssd1 vccd1 vccd1 _19464_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15649__A _16078_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15347_ _16450_/B _16450_/C _16313_/C vssd1 vssd1 vccd1 vccd1 _15347_/X sky130_fd_sc_hd__and3_1
XFILLER_191_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ _12769_/B vssd1 vssd1 vccd1 vccd1 _12645_/C sky130_fd_sc_hd__inv_2
XFILLER_145_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18066_ _18040_/A _18059_/Y _18063_/X _18067_/A vssd1 vssd1 vccd1 vccd1 _18066_/X
+ sky130_fd_sc_hd__o211a_1
X_15278_ _22880_/Q _15278_/B vssd1 vssd1 vccd1 vccd1 _22868_/D sky130_fd_sc_hd__xor2_1
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16710__A2 _16708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17017_ _17027_/A _17027_/B _17019_/A _17019_/B vssd1 vssd1 vccd1 vccd1 _17017_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_171_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18448__C1 _18200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14229_ _14238_/A _14238_/B _14239_/B vssd1 vssd1 vccd1 vccd1 _14236_/A sky130_fd_sc_hd__a21o_1
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12073__A _17039_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__A1 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__B2 _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18679__B _22798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22920__D _22920_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20270__A2 _20115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ _18968_/A _18968_/B vssd1 vssd1 vccd1 vccd1 _18972_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22547__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _17954_/A _17954_/B _17919_/C vssd1 vssd1 vccd1 vccd1 _17920_/A sky130_fd_sc_hd__or3_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18899_ _18899_/A _18899_/B _18899_/C vssd1 vssd1 vccd1 vccd1 _18900_/A sky130_fd_sc_hd__nand3_1
XANTENNA__15534__D _22964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20930_ _20930_/A _21017_/C vssd1 vssd1 vccd1 vccd1 _20930_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20861_ _20864_/B _20866_/A _20866_/B vssd1 vssd1 vccd1 vccd1 _20863_/B sky130_fd_sc_hd__nand3b_1
XFILLER_82_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22600_ _11430_/C input62/X _22608_/S vssd1 vssd1 vccd1 vccd1 _22601_/A sky130_fd_sc_hd__mux2_1
XANTENNA__20449__B _20449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19715__A2 _19792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20792_ _20792_/A _20792_/B _20792_/C vssd1 vssd1 vccd1 vccd1 _20792_/X sky130_fd_sc_hd__and3_1
XFILLER_179_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22531_ _22531_/A vssd1 vssd1 vccd1 vccd1 _22758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16943__A _18193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22462_ _13301_/X input65/X _22464_/S vssd1 vssd1 vccd1 vccd1 _22463_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_950 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21413_ _21251_/A _21251_/C _21251_/B _21299_/X vssd1 vssd1 vccd1 vccd1 _21416_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_194_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15559__A _16257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22393_ _22439_/S vssd1 vssd1 vccd1 vccd1 _22402_/S sky130_fd_sc_hd__buf_2
XANTENNA__18151__A1 _11800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21344_ _21348_/A _21848_/B _21733_/A _21344_/D vssd1 vssd1 vccd1 vccd1 _21344_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_190_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21275_ _13419_/A _13416_/B _21270_/X vssd1 vssd1 vccd1 vccd1 _21276_/C sky130_fd_sc_hd__o21a_1
XFILLER_150_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22830__D _22842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20226_ _20083_/X _20339_/A _20457_/B _20457_/A vssd1 vssd1 vccd1 vccd1 _20228_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17924__D _21081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15294__A _22886_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22667__CLK _22959_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20157_ _20154_/A _20154_/B _20155_/X _20156_/X vssd1 vssd1 vccd1 vccd1 _20158_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12711__A _20478_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20088_ _12329_/X _12803_/X _20086_/Y _20087_/Y vssd1 vssd1 vccd1 vccd1 _20088_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _11930_/A _11930_/B _11930_/C vssd1 vssd1 vccd1 vccd1 _11930_/X sky130_fd_sc_hd__and3_1
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18611__C1 _18200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _11861_/A vssd1 vssd1 vccd1 vccd1 _11861_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19167__B1 _11672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _13618_/A _13618_/B _13601_/A vssd1 vssd1 vccd1 vccd1 _13617_/B sky130_fd_sc_hd__a21oi_2
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14580_ _14602_/A _14602_/B _14602_/C vssd1 vssd1 vccd1 vccd1 _14580_/X sky130_fd_sc_hd__and3_1
XANTENNA__15460__C _15991_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ _11792_/A _11792_/B _18339_/C vssd1 vssd1 vccd1 vccd1 _11793_/B sky130_fd_sc_hd__nand3_2
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13531_ _13524_/X _13526_/X _13527_/Y _13530_/X vssd1 vssd1 vccd1 vccd1 _13538_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_159_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22729_ _22731_/CLK _22729_/D vssd1 vssd1 vccd1 vccd1 _22729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16853__A _16853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16250_ _16250_/A _16250_/B _16250_/C vssd1 vssd1 vccd1 vccd1 _16530_/A sky130_fd_sc_hd__nand3_2
X_13462_ _13185_/A _13185_/B _13577_/A vssd1 vssd1 vccd1 vccd1 _13563_/C sky130_fd_sc_hd__a21o_1
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13203__A1 _21185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15201_ _15169_/A _15169_/B _15181_/B _15174_/A _15200_/X vssd1 vssd1 vccd1 vccd1
+ _15203_/A sky130_fd_sc_hd__o311a_1
XFILLER_185_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12413_ _12413_/A vssd1 vssd1 vccd1 vccd1 _12413_/X sky130_fd_sc_hd__buf_6
XFILLER_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16181_ _15918_/X _20449_/B _16180_/X _16080_/C vssd1 vssd1 vccd1 vccd1 _16181_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__20806__C _20806_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13393_ _21234_/A _13338_/B _13354_/Y vssd1 vssd1 vccd1 vccd1 _13393_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_182_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15132_ _15132_/A _15132_/B vssd1 vssd1 vccd1 vccd1 _15132_/Y sky130_fd_sc_hd__nand2_1
XFILLER_182_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12344_ _16318_/A _12339_/X _12343_/Y vssd1 vssd1 vccd1 vccd1 _15320_/A sky130_fd_sc_hd__o21ai_1
XFILLER_181_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15188__B _15188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19940_ _19905_/A _19937_/B _19905_/C _19939_/Y vssd1 vssd1 vccd1 vccd1 _19949_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_181_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15063_ _15119_/D _15058_/A _15058_/B _15062_/Y _15059_/Y vssd1 vssd1 vccd1 vccd1
+ _15065_/B sky130_fd_sc_hd__a32o_1
XFILLER_175_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12275_ _12340_/D vssd1 vssd1 vccd1 vccd1 _12385_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14014_ _13904_/Y _13924_/A _13748_/X _14562_/A vssd1 vssd1 vccd1 vccd1 _14014_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12714__B1 _12928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19871_ _19804_/X _19736_/B _19735_/C _19807_/A vssd1 vssd1 vccd1 vccd1 _19872_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_136_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18822_ _18826_/A _18826_/B _18827_/A vssd1 vssd1 vccd1 vccd1 _18823_/C sky130_fd_sc_hd__a21boi_1
XFILLER_110_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18753_ _18753_/A _18753_/B _18753_/C vssd1 vssd1 vccd1 vccd1 _18763_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13436__B _21498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15965_ _20502_/A vssd1 vssd1 vccd1 vccd1 _17401_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17704_ _17704_/A _17704_/B vssd1 vssd1 vccd1 vccd1 _17781_/C sky130_fd_sc_hd__xor2_2
XANTENNA__15932__A _15932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14916_ _14916_/A _14916_/B _14916_/C _14916_/D vssd1 vssd1 vccd1 vccd1 _14919_/B
+ sky130_fd_sc_hd__nand4_1
X_18684_ _18684_/A vssd1 vssd1 vccd1 vccd1 _18862_/A sky130_fd_sc_hd__clkbuf_2
X_15896_ _15813_/Y _15900_/A _15778_/Y vssd1 vssd1 vccd1 vccd1 _15975_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__11674__C_N _11673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17635_ _17635_/A vssd1 vssd1 vccd1 vccd1 _17730_/A sky130_fd_sc_hd__buf_2
XFILLER_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14847_ _14847_/A _14847_/B vssd1 vssd1 vccd1 vccd1 _14848_/A sky130_fd_sc_hd__and2_1
XFILLER_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17566_ _11821_/X _17728_/A _17564_/Y _17565_/X vssd1 vssd1 vccd1 vccd1 _17574_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15370__C _16322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_720 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14778_ _14859_/A _14191_/C _14858_/A _14857_/B vssd1 vssd1 vccd1 vccd1 _14781_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19305_ _19255_/Y _19303_/Y _19253_/Y _19434_/B vssd1 vssd1 vccd1 vccd1 _19305_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_147_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16517_ _16517_/A _16517_/B vssd1 vssd1 vccd1 vccd1 _16517_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15719__B1 _15341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ _22756_/Q _22755_/Q vssd1 vssd1 vccd1 vccd1 _13738_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17497_ _17497_/A _17497_/B vssd1 vssd1 vccd1 vccd1 _17513_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12068__A _18810_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19236_ _19396_/A _19396_/B vssd1 vssd1 vccd1 vccd1 _19238_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16448_ _15335_/A _11702_/A _16256_/Y vssd1 vssd1 vccd1 vccd1 _16452_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__22915__D _22915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16482__B _22967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19167_ _14431_/A _15808_/X _11672_/A _19461_/B _19461_/C vssd1 vssd1 vccd1 vccd1
+ _19167_/Y sky130_fd_sc_hd__o2111ai_4
X_16379_ _16213_/Y _16214_/X _16636_/A _16378_/X vssd1 vssd1 vccd1 vccd1 _16386_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_191_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18118_ _18690_/A vssd1 vssd1 vccd1 vccd1 _19165_/A sky130_fd_sc_hd__buf_2
XFILLER_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19098_ _19254_/A _19254_/B _19098_/C vssd1 vssd1 vccd1 vccd1 _19098_/X sky130_fd_sc_hd__and3_1
XFILLER_105_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12515__B _22824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18049_ _18049_/A _18049_/B vssd1 vssd1 vccd1 vccd1 _18049_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12705__B1 _12967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21060_ _21061_/B _21061_/A vssd1 vssd1 vccd1 vccd1 _21097_/A sky130_fd_sc_hd__or2_1
XFILLER_28_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18202__B _18571_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20011_ _20035_/A _20057_/B _20057_/A _20010_/X vssd1 vssd1 vccd1 vccd1 _22905_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20243__A2 _15325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12531__A _22825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15655__C1 _15654_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16938__A _17133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21962_ _21606_/X _21853_/X _21957_/Y _21961_/X vssd1 vssd1 vccd1 vccd1 _21972_/B
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__12484__A2 _15774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_536 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20913_ _20913_/A vssd1 vssd1 vccd1 vccd1 _21083_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21893_ _21892_/B _21892_/C _21892_/A vssd1 vssd1 vccd1 vccd1 _21893_/X sky130_fd_sc_hd__a21o_1
XANTENNA__14458__A _15205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20844_ _20844_/A vssd1 vssd1 vccd1 vccd1 _21082_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15973__A3 _17312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20775_ _20559_/A _20667_/Y _20768_/Y _20770_/A vssd1 vssd1 vccd1 vccd1 _20775_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_80_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19687__C _19687_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18372__A1 _11345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18372__B2 _18371_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22514_ _22514_/A _22514_/B _22586_/C vssd1 vssd1 vccd1 vccd1 _22571_/A sky130_fd_sc_hd__and3_1
XFILLER_167_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16922__A2 _15792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22445_ _13659_/C input35/X _22453_/S vssd1 vssd1 vccd1 vccd1 _22446_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_216 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18124__A1 _12165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12706__A _16759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__A1 _11703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22376_ _12470_/X input57/X _22380_/S vssd1 vssd1 vccd1 vccd1 _22377_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1043 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21327_ _21318_/A _13633_/A _21323_/Y _21326_/X vssd1 vssd1 vccd1 vccd1 _21332_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_11_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12060_ _12059_/B _12247_/B _11693_/X _11565_/Y vssd1 vssd1 vccd1 vccd1 _12061_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_21258_ _22851_/Q vssd1 vssd1 vccd1 vccd1 _21689_/A sky130_fd_sc_hd__inv_2
XFILLER_132_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12172__A1 _12170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20209_ _20210_/A _20210_/B _20208_/X vssd1 vssd1 vccd1 vccd1 _20446_/B sky130_fd_sc_hd__o21ai_4
XFILLER_78_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14449__B1 _14448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21189_ _21473_/A _21188_/Y _22731_/Q vssd1 vssd1 vccd1 vccd1 _21480_/A sky130_fd_sc_hd__o21bai_2
XFILLER_131_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16848__A _16853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _15755_/A _15755_/B _15756_/B _15756_/C vssd1 vssd1 vccd1 vccd1 _15750_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12962_ _12963_/A _12963_/B _13003_/B vssd1 vssd1 vccd1 vccd1 _12962_/Y sky130_fd_sc_hd__a21boi_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input10_A wb_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18060__B1 _18023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _11566_/X _15936_/A _11392_/Y _11871_/X _11869_/X vssd1 vssd1 vccd1 vccd1
+ _11914_/B sky130_fd_sc_hd__o311a_1
X_14701_ _14571_/X _14583_/Y _14791_/B _14775_/D vssd1 vssd1 vccd1 vccd1 _14861_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_79_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15471__B _15586_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _15682_/A _15859_/A _15681_/C _15681_/D vssd1 vssd1 vccd1 vccd1 _15761_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _20182_/A _20183_/A _20182_/B vssd1 vssd1 vccd1 vccd1 _12894_/B sky130_fd_sc_hd__and3_1
XFILLER_61_804 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17420_ _17420_/A _17420_/B _17420_/C vssd1 vssd1 vccd1 vccd1 _17457_/D sky130_fd_sc_hd__nand3_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _15377_/A vssd1 vssd1 vccd1 vccd1 _15792_/B sky130_fd_sc_hd__clkbuf_4
X_14632_ _14635_/A _14635_/B _14635_/C vssd1 vssd1 vccd1 vccd1 _14632_/X sky130_fd_sc_hd__and3_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _17344_/Y _17494_/A _17206_/B vssd1 vssd1 vccd1 vccd1 _17351_/Y sky130_fd_sc_hd__a21boi_1
X_14563_ _14274_/A _14562_/X _14568_/A _14462_/Y _14463_/X vssd1 vssd1 vccd1 vccd1
+ _14602_/A sky130_fd_sc_hd__o32a_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_500 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11775_ _12018_/A _12165_/A _11774_/Y vssd1 vssd1 vccd1 vccd1 _11945_/A sky130_fd_sc_hd__o21ai_2
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16302_ _16302_/A vssd1 vssd1 vccd1 vccd1 _20605_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _21315_/B _13581_/A _13515_/A _13516_/D vssd1 vssd1 vccd1 vccd1 _13523_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15177__A1 _14845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17282_ _17282_/A vssd1 vssd1 vccd1 vccd1 _17293_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14494_ _14626_/A _14494_/B _14494_/C _14494_/D vssd1 vssd1 vccd1 vccd1 _14500_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_186_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19021_ _19014_/X _19015_/Y _19194_/A _17672_/A _19017_/Y vssd1 vssd1 vccd1 vccd1
+ _19022_/B sky130_fd_sc_hd__o2111ai_1
X_16233_ _16225_/A _16227_/A _16486_/C _17144_/C vssd1 vssd1 vccd1 vccd1 _16506_/A
+ sky130_fd_sc_hd__o211ai_4
X_13445_ _13465_/A _13465_/B _13169_/X vssd1 vssd1 vccd1 vccd1 _13455_/A sky130_fd_sc_hd__a21o_1
XFILLER_174_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12935__B1 _16937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22832__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16164_ _16174_/A _16169_/D _16163_/X vssd1 vssd1 vccd1 vccd1 _16166_/C sky130_fd_sc_hd__o21ai_1
X_13376_ _13376_/A vssd1 vssd1 vccd1 vccd1 _21522_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15115_ _15115_/A _15115_/B _15115_/C vssd1 vssd1 vccd1 vccd1 _15115_/Y sky130_fd_sc_hd__nand3_1
XFILLER_6_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12327_ _12340_/A _12284_/A _12319_/Y _12320_/Y vssd1 vssd1 vccd1 vccd1 _12418_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__20473__A2 _16745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16095_ _16090_/Y _16043_/C _16190_/B _16094_/X vssd1 vssd1 vccd1 vccd1 _16201_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18303__A _18303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19923_ _19809_/A _19809_/B _19919_/A _19823_/A vssd1 vssd1 vccd1 vccd1 _19923_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_138_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15046_ _15046_/A _15046_/B _15175_/D vssd1 vssd1 vccd1 vccd1 _15101_/A sky130_fd_sc_hd__or3b_1
X_12258_ _12258_/A _22909_/Q vssd1 vssd1 vccd1 vccd1 _12259_/B sky130_fd_sc_hd__and2_1
XFILLER_114_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14550__B _22876_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19854_ _17442_/X _19987_/C _19793_/A _19852_/Y _19853_/Y vssd1 vssd1 vccd1 vccd1
+ _19856_/B sky130_fd_sc_hd__o311a_1
XFILLER_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189_ _12189_/A _18208_/B vssd1 vssd1 vccd1 vccd1 _12189_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__21086__D _21086_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18805_ _18796_/X _18618_/A _18799_/Y _18804_/Y vssd1 vssd1 vccd1 vccd1 _18825_/A
+ sky130_fd_sc_hd__o211ai_4
Xclkbuf_4_3_0_bq_clk_i clkbuf_4_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _22937_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19785_ _19788_/B _19785_/B _19785_/C vssd1 vssd1 vccd1 vccd1 _19796_/A sky130_fd_sc_hd__nand3b_1
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16997_ _16997_/A _17313_/A _16997_/C vssd1 vssd1 vccd1 vccd1 _17001_/A sky130_fd_sc_hd__nand3_1
XFILLER_96_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18736_ _18736_/A _18736_/B _18736_/C vssd1 vssd1 vccd1 vccd1 _18743_/B sky130_fd_sc_hd__nand3_1
XFILLER_97_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15948_ _15937_/X _15942_/X _15947_/Y vssd1 vssd1 vccd1 vccd1 _15949_/B sky130_fd_sc_hd__o21ai_1
XFILLER_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18667_ _18670_/A _18827_/A _18664_/X _18666_/X vssd1 vssd1 vccd1 vccd1 _18735_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15879_ _15879_/A vssd1 vssd1 vccd1 vccd1 _15879_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15404__A2 _12607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13182__A _22735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17618_ _17615_/X _17719_/B _17617_/Y _17508_/Y vssd1 vssd1 vccd1 vccd1 _17619_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12218__A2 _12052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19788__B _19788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18598_ _18598_/A _18598_/B vssd1 vssd1 vccd1 vccd1 _18598_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17549_ _17541_/Y _17544_/Y _17663_/A _17663_/B vssd1 vssd1 vccd1 vccd1 _17552_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__17157__A2 _17270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13332__D _21739_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11977__A1 _15904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20560_ _20314_/Y _20189_/Y _20191_/A vssd1 vssd1 vccd1 vccd1 _20560_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__17739__D _20806_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19219_ _19227_/C _19227_/B vssd1 vssd1 vccd1 vccd1 _19219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_192_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18106__A1 _16921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20491_ _20455_/X _20459_/Y _20485_/Y _20490_/Y vssd1 vssd1 vccd1 vccd1 _20491_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_121_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22230_ _22172_/A _22037_/A _22037_/B _22231_/B _22231_/C vssd1 vssd1 vccd1 vccd1
+ _22232_/A sky130_fd_sc_hd__a32o_1
XFILLER_146_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19854__A1 _17442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17023__A1_N _16732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20743__A _20928_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22161_ _21908_/X _21911_/X _22024_/Y _22160_/Y vssd1 vssd1 vccd1 vccd1 _22161_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19309__A _19329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21112_ _21112_/A _21112_/B vssd1 vssd1 vccd1 vccd1 _21138_/C sky130_fd_sc_hd__xnor2_2
XFILLER_160_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22092_ _22092_/A _22092_/B _22680_/Q vssd1 vssd1 vccd1 vccd1 _22094_/A sky130_fd_sc_hd__and3_1
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21043_ _21023_/A _21023_/B _21030_/C vssd1 vssd1 vccd1 vccd1 _21061_/B sky130_fd_sc_hd__a21oi_2
XFILLER_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input2_A wb_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21724__D _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21945_ _22041_/C vssd1 vssd1 vccd1 vccd1 _22037_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__20259__B1_N _20263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20924__B1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17396__A2 _17822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16053__C1 _12988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13092__A _22842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11605__A _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21876_ _21876_/A vssd1 vssd1 vccd1 vccd1 _22221_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ _20827_/A _20827_/B _20827_/C _20827_/D vssd1 vssd1 vccd1 vccd1 _20828_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_126_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22855__CLK _22937_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11560_ _11668_/A _15539_/A _11560_/C vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__nand3_4
XFILLER_168_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20152__A1 _20143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20758_ _20758_/A _20758_/B vssd1 vssd1 vccd1 vccd1 _20890_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17649__D _18303_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18107__B _18107_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14906__A1 _14670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ _11709_/B vssd1 vssd1 vccd1 vccd1 _18453_/C sky130_fd_sc_hd__buf_4
XFILLER_195_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20689_ _20936_/B _20793_/C vssd1 vssd1 vccd1 vccd1 _20689_/Y sky130_fd_sc_hd__nand2_1
XFILLER_137_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13230_ _13234_/A vssd1 vssd1 vccd1 vccd1 _13230_/X sky130_fd_sc_hd__buf_2
XFILLER_155_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22428_ _22428_/A vssd1 vssd1 vccd1 vccd1 _22713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _13161_/A _21336_/C _13161_/C vssd1 vssd1 vccd1 vccd1 _13162_/C sky130_fd_sc_hd__and3_2
XFILLER_164_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22359_ _21700_/X _21701_/X _22352_/A vssd1 vssd1 vccd1 vccd1 _22359_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_3_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12112_ _12112_/A vssd1 vssd1 vccd1 vccd1 _16274_/A sky130_fd_sc_hd__buf_2
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14134__A2 _13833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13092_ _22842_/Q vssd1 vssd1 vccd1 vccd1 _13319_/A sky130_fd_sc_hd__clkinv_2
XANTENNA_input58_A wb_dat_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16920_ _16014_/A _17443_/A _16911_/X _16913_/X vssd1 vssd1 vccd1 vccd1 _16920_/Y
+ sky130_fd_sc_hd__o22ai_4
X_12043_ _12043_/A _15536_/A _12235_/B vssd1 vssd1 vccd1 vccd1 _16477_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13267__A _22847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19073__A2 _11626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17084__A1 _11636_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16851_ _16851_/A vssd1 vssd1 vccd1 vccd1 _16853_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__18281__B1 _18453_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17084__B2 _17083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15482__A _15482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15802_ _15793_/Y _15794_/X _15829_/A vssd1 vssd1 vccd1 vccd1 _15803_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__15634__A2 _15718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19570_ _19571_/A _19571_/B _22918_/Q vssd1 vssd1 vccd1 vccd1 _19574_/A sky130_fd_sc_hd__a21o_1
XFILLER_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16782_ _16782_/A vssd1 vssd1 vccd1 vccd1 _16782_/X sky130_fd_sc_hd__clkbuf_2
X_13994_ _14686_/B _14770_/A _14771_/A _13984_/Y _13986_/Y vssd1 vssd1 vccd1 vccd1
+ _13998_/A sky130_fd_sc_hd__a32o_1
X_18521_ _18490_/B _18490_/C _18490_/A vssd1 vssd1 vccd1 vccd1 _18916_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__11656__B1 _15435_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _15733_/A _15733_/B _15733_/C vssd1 vssd1 vccd1 vccd1 _15825_/C sky130_fd_sc_hd__nand3_2
XFILLER_19_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12945_ _20129_/B vssd1 vssd1 vccd1 vccd1 _20249_/C sky130_fd_sc_hd__clkbuf_4
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18452_ _12018_/X _16248_/X _18448_/Y vssd1 vssd1 vccd1 vccd1 _18452_/X sky130_fd_sc_hd__o21a_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _15664_/A vssd1 vssd1 vccd1 vccd1 _15666_/A sky130_fd_sc_hd__inv_2
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20391__A1 _12761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _15746_/B vssd1 vssd1 vccd1 vccd1 _12876_/X sky130_fd_sc_hd__buf_4
XFILLER_61_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15937__A3 _15792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _17403_/A vssd1 vssd1 vccd1 vccd1 _17647_/A sky130_fd_sc_hd__buf_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _14506_/Y _14612_/X _14892_/D _14614_/Y _14917_/C vssd1 vssd1 vccd1 vccd1
+ _14621_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_61_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18383_ _18383_/A _18383_/B vssd1 vssd1 vccd1 vccd1 _18383_/Y sky130_fd_sc_hd__nand2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11827_ _11687_/Y _11643_/Y _11689_/Y _11690_/Y vssd1 vssd1 vccd1 vccd1 _11829_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_15595_ _16287_/A _16287_/B _16286_/A vssd1 vssd1 vccd1 vccd1 _15672_/B sky130_fd_sc_hd__nand3_1
XFILLER_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17334_/A _17334_/B vssd1 vssd1 vccd1 vccd1 _17335_/A sky130_fd_sc_hd__nand2_1
XFILLER_14_572 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11745_/B _11757_/Y _11623_/X vssd1 vssd1 vccd1 vccd1 _11758_/Y sky130_fd_sc_hd__o21ai_1
X_14546_ _14547_/B _14547_/C _14547_/A vssd1 vssd1 vccd1 vccd1 _14548_/A sky130_fd_sc_hd__a21oi_1
XFILLER_92_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_594 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16898__A1 _17502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17265_ _17146_/Y _17264_/Y _17180_/A _17180_/C vssd1 vssd1 vccd1 vccd1 _17299_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_147_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14477_ _13986_/B _14568_/A _14131_/X _14468_/Y _15069_/A vssd1 vssd1 vccd1 vccd1
+ _14478_/C sky130_fd_sc_hd__o2111ai_4
X_11689_ _11689_/A vssd1 vssd1 vccd1 vccd1 _11689_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19004_ _19085_/A _19085_/B _19086_/A _19086_/B vssd1 vssd1 vccd1 vccd1 _19004_/Y
+ sky130_fd_sc_hd__nand4_4
XANTENNA__19445__B1_N _22917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16216_ _16216_/A _16216_/B vssd1 vssd1 vccd1 vccd1 _16530_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15570__A1 _15580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13428_ _13428_/A _13428_/B vssd1 vssd1 vccd1 vccd1 _13433_/C sky130_fd_sc_hd__nand2_1
X_17196_ _17196_/A _17196_/B _17200_/B _17200_/C vssd1 vssd1 vccd1 vccd1 _17197_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_127_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19774__D _19774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16147_ _16137_/C _16137_/A _16137_/B _16143_/Y vssd1 vssd1 vccd1 vccd1 _16147_/Y
+ sky130_fd_sc_hd__a31oi_1
X_13359_ _13359_/A vssd1 vssd1 vccd1 vccd1 _13359_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14561__A _15182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16078_ _16129_/C _16078_/B _16078_/C vssd1 vssd1 vccd1 vccd1 _16080_/B sky130_fd_sc_hd__and3_1
XANTENNA__12136__A1 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19906_ _19905_/A _19937_/B _19905_/C _19939_/A vssd1 vssd1 vccd1 vccd1 _19907_/B
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__17872__A _21083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15029_ _15088_/A _15030_/B _15030_/C vssd1 vssd1 vccd1 vccd1 _15031_/B sky130_fd_sc_hd__a21o_1
XFILLER_130_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13884__A1 _13851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18687__B _18876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19837_ _19837_/A _19837_/B vssd1 vssd1 vccd1 vccd1 _19856_/A sky130_fd_sc_hd__and2_1
XFILLER_151_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18811__A2 _16758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16488__A _16488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19768_ _19842_/A _19768_/B _19768_/C _19768_/D vssd1 vssd1 vccd1 vccd1 _19836_/D
+ sky130_fd_sc_hd__nand4_4
Xinput2 wb_adr_i[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__15823__C _19614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18719_ _11511_/X _18718_/X _18869_/A _18862_/A vssd1 vssd1 vccd1 vccd1 _18722_/B
+ sky130_fd_sc_hd__o211ai_2
X_19699_ _15522_/X _15521_/X _15523_/X _19695_/A vssd1 vssd1 vccd1 vccd1 _19699_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21174__A3 _13162_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22878__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21730_ _21730_/A _21730_/B _21730_/C _21730_/D vssd1 vssd1 vccd1 vccd1 _21732_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_92_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17679__A_N _17669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16050__A2 _20745_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21661_ _21654_/X _21642_/Y _21618_/Y _21624_/Y _21647_/Y vssd1 vssd1 vccd1 vccd1
+ _21661_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18208__A _18208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20612_ _20685_/A _15723_/X _15939_/A _20611_/Y _20606_/Y vssd1 vssd1 vccd1 vccd1
+ _20613_/C sky130_fd_sc_hd__o221ai_2
XFILLER_33_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21592_ _21587_/Y _21589_/Y _21591_/Y vssd1 vssd1 vccd1 vccd1 _21771_/A sky130_fd_sc_hd__o21bai_1
XANTENNA__21331__B1 _21591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20543_ _20658_/B _20658_/C vssd1 vssd1 vccd1 vccd1 _20543_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15561__A1 _12111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20474_ _20587_/A _20462_/A _20579_/C _16344_/A _20581_/A vssd1 vssd1 vccd1 vccd1
+ _20475_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_152_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22213_ _22200_/Y _21932_/Y _22166_/Y vssd1 vssd1 vccd1 vccd1 _22213_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_192_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22144_ _22142_/A _22142_/B _22143_/X vssd1 vssd1 vccd1 vccd1 _22156_/B sky130_fd_sc_hd__a21o_1
XFILLER_134_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14667__A3 _14843_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19055__A2 _18203_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22075_ _22075_/A _22075_/B vssd1 vssd1 vccd1 vccd1 _22075_/X sky130_fd_sc_hd__and2_1
XFILLER_86_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21026_ _21027_/A _21027_/B vssd1 vssd1 vccd1 vccd1 _21030_/B sky130_fd_sc_hd__nor2_1
XANTENNA__19460__C1 _19614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11319__B _18985_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15452__D _15997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _12602_/Y _12613_/Y _12601_/Y vssd1 vssd1 vccd1 vccd1 _12917_/A sky130_fd_sc_hd__o21ai_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21928_ _21925_/Y _21927_/X _21922_/Y vssd1 vssd1 vccd1 vccd1 _21929_/B sky130_fd_sc_hd__a21oi_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16041__A2 _15932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12661_ _15810_/C vssd1 vssd1 vccd1 vccd1 _12913_/A sky130_fd_sc_hd__buf_2
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _21964_/A _21725_/Y _21958_/A _21852_/Y _21854_/X vssd1 vssd1 vccd1 vccd1
+ _21859_/X sky130_fd_sc_hd__o311a_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18118__A _18690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16564__C _16996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11612_ _18648_/D vssd1 vssd1 vccd1 vccd1 _18665_/A sky130_fd_sc_hd__clkbuf_4
X_14400_ _22772_/Q _14322_/X _14396_/X _22740_/Q _14399_/X vssd1 vssd1 vccd1 vccd1
+ _14400_/X sky130_fd_sc_hd__a221o_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _15415_/C vssd1 vssd1 vccd1 vccd1 _16062_/A sky130_fd_sc_hd__clkbuf_4
X_12592_ _12592_/A _12592_/B vssd1 vssd1 vccd1 vccd1 _12592_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20086__C _20463_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14331_ _22369_/D vssd1 vssd1 vccd1 vccd1 _14331_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11543_ _11541_/X _18371_/A _11533_/A vssd1 vssd1 vccd1 vccd1 _11645_/A sky130_fd_sc_hd__o21ai_2
XFILLER_184_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17050_ _16882_/X _16637_/Y _16638_/Y _16895_/A _16644_/C vssd1 vssd1 vccd1 vccd1
+ _17050_/X sky130_fd_sc_hd__a32o_1
X_14262_ _14261_/C _14261_/B _14272_/A vssd1 vssd1 vccd1 vccd1 _14263_/C sky130_fd_sc_hd__a21bo_1
XFILLER_184_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11474_ _11542_/A vssd1 vssd1 vccd1 vccd1 _11474_/X sky130_fd_sc_hd__buf_4
XFILLER_137_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16001_ _16045_/B _15986_/Y _15995_/Y _16046_/A vssd1 vssd1 vccd1 vccd1 _16003_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_100_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13213_ _13434_/A vssd1 vssd1 vccd1 vccd1 _13213_/X sky130_fd_sc_hd__buf_2
XFILLER_87_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14193_ _14222_/A _14494_/C _14195_/D _14195_/A vssd1 vssd1 vccd1 vccd1 _14198_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13144_ _13144_/A vssd1 vssd1 vccd1 vccd1 _13161_/A sky130_fd_sc_hd__buf_2
XFILLER_83_1018 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17952_ _17957_/A _17957_/B vssd1 vssd1 vccd1 vccd1 _17953_/B sky130_fd_sc_hd__or2_1
XFILLER_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _22729_/Q vssd1 vssd1 vccd1 vccd1 _13304_/B sky130_fd_sc_hd__buf_2
XFILLER_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16903_ _16702_/B _16663_/Y _16700_/B _16675_/Y vssd1 vssd1 vccd1 vccd1 _16903_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12026_ _12088_/A vssd1 vssd1 vccd1 vccd1 _12055_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_78_553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11877__B1 _11349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17883_ _19839_/B _17883_/B _21044_/B _17883_/D vssd1 vssd1 vccd1 vccd1 _17885_/A
+ sky130_fd_sc_hd__or4_1
X_19622_ _18107_/B _18107_/C _19772_/B _19621_/B _19621_/C vssd1 vssd1 vccd1 vccd1
+ _19622_/X sky130_fd_sc_hd__a32o_1
X_16834_ _16834_/A _17189_/B vssd1 vssd1 vccd1 vccd1 _16840_/A sky130_fd_sc_hd__nand2_1
XFILLER_120_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13725__A _13725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18006__B1 _22905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19553_ _19455_/C _19418_/C _19455_/A _19454_/X vssd1 vssd1 vccd1 vccd1 _19553_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11629__B1 _17312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16765_ _16489_/X _16496_/X _16507_/X _16506_/X vssd1 vssd1 vccd1 vccd1 _16768_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13977_ _22858_/D _14911_/C _14911_/A _14002_/B _14002_/C vssd1 vssd1 vccd1 vccd1
+ _14009_/C sky130_fd_sc_hd__a32o_1
X_18504_ _18876_/A vssd1 vssd1 vccd1 vccd1 _18706_/B sky130_fd_sc_hd__buf_2
XFILLER_19_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15716_ _15406_/X _15404_/X _15711_/A _15403_/X _17128_/B vssd1 vssd1 vccd1 vccd1
+ _15752_/B sky130_fd_sc_hd__o2111ai_4
XANTENNA__15940__A _15940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19484_ _19636_/A _19636_/B vssd1 vssd1 vccd1 vccd1 _19486_/A sky130_fd_sc_hd__nand2_1
XFILLER_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _12928_/A vssd1 vssd1 vccd1 vccd1 _12928_/X sky130_fd_sc_hd__buf_2
X_16696_ _16692_/X _16693_/Y _16694_/Y _16695_/X vssd1 vssd1 vccd1 vccd1 _16697_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_34_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12841__A2 _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19769__D _19836_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18435_ _18435_/A _18435_/B vssd1 vssd1 vccd1 vccd1 _22891_/D sky130_fd_sc_hd__xnor2_1
X_15647_ _15647_/A vssd1 vssd1 vccd1 vccd1 _16400_/A sky130_fd_sc_hd__buf_2
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12859_ _12859_/A _12859_/B vssd1 vssd1 vccd1 vccd1 _20120_/B sky130_fd_sc_hd__nand2_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19506__B1 _17532_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18366_ _11744_/X _18123_/Y _18154_/X vssd1 vssd1 vccd1 vccd1 _18366_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__11899__B _11899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15578_ _15566_/X _15571_/Y _15574_/X _15577_/X vssd1 vssd1 vccd1 vccd1 _15583_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17317_ _17520_/A _17520_/D vssd1 vssd1 vccd1 vccd1 _17318_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14529_ _13957_/A _14527_/Y _14528_/Y vssd1 vssd1 vccd1 vccd1 _14530_/B sky130_fd_sc_hd__a21oi_1
X_18297_ _18293_/X _18294_/X _18295_/Y _18296_/Y vssd1 vssd1 vccd1 vccd1 _18305_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__16771__A _16771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17248_ _16778_/X _16779_/X _17405_/A _17406_/A vssd1 vssd1 vccd1 vccd1 _17257_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_388 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17179_ _17173_/C _17173_/D _17178_/Y vssd1 vssd1 vccd1 vccd1 _17184_/A sky130_fd_sc_hd__a21o_1
XFILLER_155_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16099__A2 _16098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14722__C _14722_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20190_ _20189_/A _20186_/Y _20189_/Y vssd1 vssd1 vccd1 vccd1 _20191_/B sky130_fd_sc_hd__o21ai_2
XFILLER_143_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12109__A1 _15714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18698__A _18698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13306__B1 _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18848__D _18848_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17752__D _20972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18796__A1 _11474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22900_ _22951_/CLK _22900_/D vssd1 vssd1 vccd1 vccd1 _22900_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_5_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15553__C _15774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16011__A _16011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19025__C _19496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16271__A2 _15933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22831_ _22850_/CLK _22843_/Q vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19322__A _19322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22762_ _22762_/CLK _22762_/D vssd1 vssd1 vccd1 vccd1 _22762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_634 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12832__A2 _12827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21713_ _21713_/A _22851_/Q _21713_/C vssd1 vssd1 vccd1 vccd1 _21714_/A sky130_fd_sc_hd__and3_1
XFILLER_52_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22693_ _22693_/CLK _22693_/D vssd1 vssd1 vccd1 vccd1 _22693_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21644_ _21504_/A _21504_/B _21504_/C _21501_/B _21501_/A vssd1 vssd1 vccd1 vccd1
+ _21649_/A sky130_fd_sc_hd__a32oi_4
XFILLER_36_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18880__B _18880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21575_ _21551_/A _21551_/B _21421_/A vssd1 vssd1 vccd1 vccd1 _21576_/B sky130_fd_sc_hd__o21a_1
XFILLER_138_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20526_ _20526_/A _20526_/B _20526_/C vssd1 vssd1 vccd1 vccd1 _20534_/A sky130_fd_sc_hd__nand3_2
XANTENNA__22833__D _22845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16731__B1 _20793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15297__A _15297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20457_ _20457_/A _20457_/B vssd1 vssd1 vccd1 vccd1 _20457_/Y sky130_fd_sc_hd__nand2_1
XFILLER_137_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15728__C _16308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20388_ _20388_/A _20388_/B _20388_/C vssd1 vssd1 vccd1 vccd1 _20388_/Y sky130_fd_sc_hd__nand3_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15298__B1 _14430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16495__C1 _16100_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22127_ _22128_/A _22219_/A _22128_/C vssd1 vssd1 vccd1 vccd1 _22129_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22058_ _22058_/A vssd1 vssd1 vccd1 vccd1 _22223_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19216__B _19496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21009_ _21009_/A vssd1 vssd1 vccd1 vccd1 _21082_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13900_ _13810_/A _13833_/B _13810_/B _14571_/A _13815_/X vssd1 vssd1 vccd1 vccd1
+ _13902_/A sky130_fd_sc_hd__a311o_1
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14880_ _14880_/A _14880_/B _14880_/C vssd1 vssd1 vccd1 vccd1 _14880_/X sky130_fd_sc_hd__and3_1
XFILLER_43_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13831_ _13831_/A vssd1 vssd1 vccd1 vccd1 _14074_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16550_ _12827_/X _15617_/X _11779_/C _11779_/B _20675_/A vssd1 vssd1 vccd1 vccd1
+ _16550_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_56_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13762_ _13948_/A _13949_/A vssd1 vssd1 vccd1 vccd1 _13763_/A sky130_fd_sc_hd__nand2_1
XFILLER_189_915 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15501_ _15501_/A vssd1 vssd1 vccd1 vccd1 _15502_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12713_ _20255_/B vssd1 vssd1 vccd1 vccd1 _12928_/A sky130_fd_sc_hd__buf_2
X_16481_ _16481_/A _16481_/B _16481_/C _16481_/D vssd1 vssd1 vccd1 vccd1 _16483_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13693_ _14199_/A vssd1 vssd1 vccd1 vccd1 _14222_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18220_ _18276_/A _18277_/A _18276_/B vssd1 vssd1 vccd1 vccd1 _18220_/Y sky130_fd_sc_hd__nand3_1
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15432_ _15517_/A _15512_/B _15512_/C _15700_/B _15431_/Y vssd1 vssd1 vccd1 vccd1
+ _15433_/A sky130_fd_sc_hd__a32oi_4
XFILLER_176_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12644_ _12645_/A _12769_/A _12645_/C vssd1 vssd1 vccd1 vccd1 _12644_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18151_ _11800_/X _12167_/X _18139_/X _18137_/Y _18141_/Y vssd1 vssd1 vccd1 vccd1
+ _18389_/C sky130_fd_sc_hd__o221ai_4
X_15363_ _15369_/A _16322_/B _15363_/C vssd1 vssd1 vccd1 vccd1 _20341_/B sky130_fd_sc_hd__nand3_1
X_12575_ _16947_/A _20101_/C _12988_/B _12420_/X vssd1 vssd1 vccd1 vccd1 _12583_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_168_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17102_ _17103_/A _17338_/B _17103_/C vssd1 vssd1 vccd1 vccd1 _17196_/A sky130_fd_sc_hd__a21o_1
XFILLER_15_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14314_ _22586_/D _22586_/B vssd1 vssd1 vccd1 vccd1 _22514_/B sky130_fd_sc_hd__and2b_1
X_18082_ _22908_/Q _18082_/B _18082_/C vssd1 vssd1 vccd1 vccd1 _18084_/A sky130_fd_sc_hd__nand3b_1
XFILLER_172_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15525__A1 _12209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11526_ _11526_/A vssd1 vssd1 vccd1 vccd1 _15797_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15294_ _22886_/Q _15294_/B vssd1 vssd1 vccd1 vccd1 _22874_/D sky130_fd_sc_hd__xor2_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17033_ _17033_/A _17033_/B _17033_/C vssd1 vssd1 vccd1 vccd1 _17040_/A sky130_fd_sc_hd__nand3_1
XFILLER_144_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11457_ _11659_/B vssd1 vssd1 vccd1 vccd1 _11675_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14245_ _14245_/A _14245_/B vssd1 vssd1 vccd1 vccd1 _14282_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17278__A1 _16275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14176_ _14285_/C _14285_/A _14285_/B vssd1 vssd1 vccd1 vccd1 _14180_/A sky130_fd_sc_hd__a21boi_1
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11388_ _11404_/B _11423_/A _11404_/D _11404_/A _11727_/C vssd1 vssd1 vccd1 vccd1
+ _18482_/A sky130_fd_sc_hd__o311ai_4
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12343__B _12343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15357__D _18985_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _21351_/A _21351_/B vssd1 vssd1 vccd1 vccd1 _21606_/A sky130_fd_sc_hd__nand2_2
XANTENNA__15935__A _15935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19019__A2 _17422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18984_ _18984_/A _18984_/B _19480_/A _19481_/A vssd1 vssd1 vccd1 vccd1 _18984_/Y
+ sky130_fd_sc_hd__nand4_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _19987_/A _21082_/C _17935_/C _17974_/A vssd1 vssd1 vccd1 vccd1 _17991_/A
+ sky130_fd_sc_hd__or4_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _22735_/Q vssd1 vssd1 vccd1 vccd1 _21307_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12009_ _12009_/A vssd1 vssd1 vccd1 vccd1 _12009_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_61_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16469__C _16842_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater127 _22877_/Q vssd1 vssd1 vccd1 vccd1 _15279_/A sky130_fd_sc_hd__clkbuf_1
X_17866_ _17866_/A _18007_/A _18007_/B vssd1 vssd1 vccd1 vccd1 _17868_/A sky130_fd_sc_hd__nor3_1
Xrepeater138 _22791_/CLK vssd1 vssd1 vccd1 vccd1 _22789_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_16_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater149 _22807_/CLK vssd1 vssd1 vccd1 vccd1 _22808_/CLK sky130_fd_sc_hd__clkbuf_1
X_19605_ _19605_/A _19605_/B _19605_/C vssd1 vssd1 vccd1 vccd1 _19605_/Y sky130_fd_sc_hd__nand3_1
X_16817_ _20605_/A vssd1 vssd1 vccd1 vccd1 _20928_/A sky130_fd_sc_hd__buf_2
XFILLER_66_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17797_ _17797_/A _18007_/A vssd1 vssd1 vccd1 vccd1 _22961_/D sky130_fd_sc_hd__nor2_1
XFILLER_94_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19536_ _19536_/A _19536_/B _19536_/C _19536_/D vssd1 vssd1 vccd1 vccd1 _19540_/B
+ sky130_fd_sc_hd__nand4_1
X_16748_ _16738_/X _16736_/Y _16747_/X _16723_/X vssd1 vssd1 vccd1 vccd1 _16749_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_59_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22918__D _22918_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19467_ _11737_/X _11738_/X _15810_/A _19618_/A _19323_/X vssd1 vssd1 vccd1 vccd1
+ _19467_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16679_ _16406_/A _16406_/B _15881_/A _16686_/A vssd1 vssd1 vccd1 vccd1 _16683_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18981__A _19694_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18418_ _18416_/A _18417_/A _18216_/B _18216_/A vssd1 vssd1 vccd1 vccd1 _18418_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_34_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19398_ _19398_/A _19458_/B _19398_/C vssd1 vssd1 vccd1 vccd1 _19399_/C sky130_fd_sc_hd__nand3_1
XFILLER_22_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22916__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18349_ _18349_/A _18349_/B vssd1 vssd1 vccd1 vccd1 _18351_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16932__C _16932_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15516__A1 _15755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21360_ _21393_/A _21388_/A vssd1 vssd1 vccd1 vccd1 _21379_/A sky130_fd_sc_hd__nand2_1
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16713__B1 _16712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20311_ _20311_/A _20311_/B _20311_/C vssd1 vssd1 vccd1 vccd1 _20313_/A sky130_fd_sc_hd__nand3_1
XANTENNA__20454__C _20454_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput60 wb_dat_i[3] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_4
X_21291_ _21292_/C _21292_/A _22673_/Q vssd1 vssd1 vccd1 vccd1 _21294_/C sky130_fd_sc_hd__a21oi_2
Xinput71 x[11] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18466__B1 _19046_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20242_ _20242_/A vssd1 vssd1 vccd1 vccd1 _20242_/X sky130_fd_sc_hd__buf_2
XFILLER_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20273__B1 _20398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20173_ _20182_/B _20182_/A _20183_/A vssd1 vssd1 vccd1 vccd1 _20174_/C sky130_fd_sc_hd__a21boi_1
XFILLER_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15295__A3 _22886_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21285__C _21285_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12502__A1 _12500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18875__B _18876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17441__A1 _17442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17441__B2 _16015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19718__B1 _19788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15580__A _15580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22814_ _22815_/CLK _22814_/D vssd1 vssd1 vccd1 vccd1 _22814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17729__C1 _17922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22745_ _22746_/CLK _22745_/D vssd1 vssd1 vccd1 vccd1 _22745_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15204__B1 _15205_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19202__D _19202_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11613__A _12094_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22676_ _22943_/CLK _22676_/D vssd1 vssd1 vccd1 vccd1 _22676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16952__B1 _12930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22617__S _22619_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12569__A1 _12470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21627_ _13344_/X _13345_/X _21853_/A vssd1 vssd1 vccd1 vccd1 _21631_/A sky130_fd_sc_hd__a21o_1
XANTENNA__15507__A1 _15580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16842__C _16842_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12360_ _12457_/A _12687_/B vssd1 vssd1 vccd1 vccd1 _12374_/A sky130_fd_sc_hd__nand2_1
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21558_ _21558_/A vssd1 vssd1 vccd1 vccd1 _21930_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_87 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_995 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11311_ _11404_/A vssd1 vssd1 vccd1 vccd1 _11311_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20509_ _16778_/X _16779_/X _20505_/Y _20913_/A _20503_/Y vssd1 vssd1 vccd1 vccd1
+ _20511_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_10_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16180__A1 _15890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12291_ _12421_/A _12822_/A _12385_/A _12384_/A vssd1 vssd1 vccd1 vccd1 _12292_/A
+ sky130_fd_sc_hd__nand4_4
X_21489_ _21489_/A _21872_/A vssd1 vssd1 vccd1 vccd1 _21490_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16180__B2 _16179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14030_ _14052_/C _14052_/B vssd1 vssd1 vccd1 vccd1 _14036_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21757__A _21757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12163__B _18093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15755__A _15755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18472__A3 _17442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18131__A _18328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input40_A wb_dat_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15981_ _18512_/A vssd1 vssd1 vccd1 vccd1 _15981_/X sky130_fd_sc_hd__buf_4
XANTENNA__21195__C _21195_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15691__B1 _16498_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17720_ _17720_/A _17720_/B _17720_/C vssd1 vssd1 vccd1 vccd1 _17795_/A sky130_fd_sc_hd__nand3_1
XANTENNA__17970__A _22903_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14932_ _14932_/A vssd1 vssd1 vccd1 vccd1 _14996_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_102_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22588__A _22656_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17651_ _19689_/C vssd1 vssd1 vccd1 vccd1 _19585_/D sky130_fd_sc_hd__buf_2
XANTENNA__18090__D1 _15690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14863_ _14863_/A _14863_/B _14863_/C vssd1 vssd1 vccd1 vccd1 _14865_/A sky130_fd_sc_hd__nand3_4
XFILLER_21_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17983__A2 _21017_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16602_ _16602_/A _16602_/B _16602_/C vssd1 vssd1 vccd1 vccd1 _16617_/C sky130_fd_sc_hd__nand3_1
XFILLER_17_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13814_ _13814_/A _13814_/B vssd1 vssd1 vccd1 vccd1 _14126_/A sky130_fd_sc_hd__nand2_2
XFILLER_91_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17582_ _17627_/A _17581_/B _17553_/A _17580_/A vssd1 vssd1 vccd1 vccd1 _17582_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15921__C _17652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14794_ _14685_/B _14862_/A _14935_/A _13873_/X _14793_/Y vssd1 vssd1 vccd1 vccd1
+ _14884_/C sky130_fd_sc_hd__o2111ai_4
X_19321_ _19317_/Y _19319_/Y _19320_/X vssd1 vssd1 vccd1 vccd1 _19321_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_44_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16533_ _16250_/A _16532_/Y _16529_/B _16529_/C vssd1 vssd1 vccd1 vccd1 _16534_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__22939__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13745_ _13736_/C _13745_/B _13745_/C vssd1 vssd1 vccd1 vccd1 _13750_/B sky130_fd_sc_hd__nand3b_1
XFILLER_73_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19252_ _19251_/Y _19248_/Y _19249_/Y vssd1 vssd1 vccd1 vccd1 _19252_/X sky130_fd_sc_hd__a21o_1
XFILLER_149_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16464_ _16469_/B vssd1 vssd1 vccd1 vccd1 _16842_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13676_ _13617_/B _13617_/A _13609_/Y vssd1 vssd1 vccd1 vccd1 _13678_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18203_ _18203_/A _18203_/B _18203_/C _18282_/A vssd1 vssd1 vccd1 vccd1 _18204_/A
+ sky130_fd_sc_hd__or4_2
X_15415_ _20675_/A _20675_/B _15415_/C vssd1 vssd1 vccd1 vccd1 _15415_/X sky130_fd_sc_hd__and3_2
XFILLER_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19183_ _19530_/A _19343_/A _19240_/C _19240_/D vssd1 vssd1 vccd1 vccd1 _19237_/C
+ sky130_fd_sc_hd__nand4_4
X_12627_ _15586_/C _20502_/C _12557_/A _12557_/B vssd1 vssd1 vccd1 vccd1 _12628_/B
+ sky130_fd_sc_hd__a22o_1
X_16395_ _20917_/B vssd1 vssd1 vccd1 vccd1 _20975_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_129_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18145__C1 _15988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14834__A _14834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18134_ _18690_/A _18483_/B vssd1 vssd1 vccd1 vccd1 _18135_/A sky130_fd_sc_hd__nand2_2
XFILLER_89_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15346_ _15633_/B vssd1 vssd1 vccd1 vccd1 _16450_/B sky130_fd_sc_hd__buf_2
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12558_ _20514_/A _12671_/A _12790_/A _12672_/A _12628_/A vssd1 vssd1 vccd1 vccd1
+ _12769_/B sky130_fd_sc_hd__o41a_2
XFILLER_157_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18065_ _18065_/A _18065_/B _18065_/C vssd1 vssd1 vccd1 vccd1 _18067_/A sky130_fd_sc_hd__and3_1
XFILLER_117_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11509_ _12090_/C vssd1 vssd1 vccd1 vccd1 _18512_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15277_ _15279_/A _22878_/Q _22879_/Q _15288_/C vssd1 vssd1 vccd1 vccd1 _15278_/B
+ sky130_fd_sc_hd__o31a_1
X_12489_ _12484_/Y _12487_/X _12358_/X _12488_/Y vssd1 vssd1 vccd1 vccd1 _12489_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_144_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17016_ _16732_/Y _16742_/Y _16726_/Y _17025_/A _17025_/B vssd1 vssd1 vccd1 vccd1
+ _17019_/B sky130_fd_sc_hd__o2111ai_4
XANTENNA__18448__B1 _18107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21047__A2 _17839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14228_ _14273_/A _15154_/B _14226_/A vssd1 vssd1 vccd1 vccd1 _14243_/B sky130_fd_sc_hd__a21oi_1
XFILLER_172_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12073__B _19046_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15665__A _15665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21452__C1 _21805_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _14272_/C _14857_/A _14161_/C _14161_/B vssd1 vssd1 vccd1 vccd1 _14159_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18967_ _22914_/Q _18967_/B vssd1 vssd1 vccd1 vccd1 _18968_/B sky130_fd_sc_hd__or2_1
XFILLER_140_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12801__B _20605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17880__A _17880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17918_ _18007_/C _17918_/B vssd1 vssd1 vccd1 vccd1 _22963_/D sky130_fd_sc_hd__xnor2_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18898_ _18895_/X _19022_/C _18901_/A _19009_/A vssd1 vssd1 vccd1 vccd1 _18899_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_6_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17849_ _17775_/X _17847_/Y _17848_/Y vssd1 vssd1 vccd1 vccd1 _17849_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_93_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15434__B1 _12758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20860_ _20793_/Y _20860_/B _20860_/C vssd1 vssd1 vccd1 vccd1 _20866_/B sky130_fd_sc_hd__nand3b_2
XFILLER_93_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19519_ _19581_/A _19521_/C _19516_/Y _19518_/X vssd1 vssd1 vccd1 vccd1 _19532_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__19715__A3 _19615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20791_ _12928_/X _17435_/A _20790_/Y vssd1 vssd1 vccd1 vccd1 _20791_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11433__A _11942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22530_ _13799_/X input63/X _22536_/S vssd1 vssd1 vccd1 vccd1 _22531_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22437__S _22439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12248__B _12250_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22461_ _22461_/A vssd1 vssd1 vccd1 vccd1 _22727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21412_ _21251_/X _21299_/X _21417_/B _21553_/A vssd1 vssd1 vccd1 vccd1 _21415_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_182_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_962 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15559__B _15559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22392_ _22392_/A vssd1 vssd1 vccd1 vccd1 _22697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18151__A2 _12167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21343_ _21343_/A vssd1 vssd1 vccd1 vccd1 _21733_/A sky130_fd_sc_hd__buf_2
XFILLER_194_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21274_ _21265_/Y _21266_/Y _21263_/Y _21257_/Y vssd1 vssd1 vccd1 vccd1 _21419_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_118_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20481__A _20579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15575__A _18848_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20225_ _20093_/B _20219_/Y _20090_/Y vssd1 vssd1 vccd1 vccd1 _20228_/A sky130_fd_sc_hd__o21a_1
XFILLER_150_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20156_ _12788_/B _12792_/C _20143_/Y _20144_/Y vssd1 vssd1 vccd1 vccd1 _20156_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13807__B _14270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20087_ _16294_/X _16293_/X _20466_/B _16302_/A vssd1 vssd1 vccd1 vccd1 _20087_/Y
+ sky130_fd_sc_hd__o211ai_2
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21746__B1 _22057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17414__A1 _15941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18611__B1 _17380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12239__B1 _12240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11860_ _11860_/A _11860_/B _11860_/C vssd1 vssd1 vccd1 vccd1 _11861_/A sky130_fd_sc_hd__and3_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19167__A1 _14431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20359__C _20359_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _11969_/A vssd1 vssd1 vccd1 vccd1 _11791_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_710 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20989_ _20989_/A _20992_/C vssd1 vssd1 vccd1 vccd1 _20990_/B sky130_fd_sc_hd__nor2_1
X_13530_ _13563_/A _13563_/B _13563_/C _13528_/X _13529_/Y vssd1 vssd1 vccd1 vccd1
+ _13530_/X sky130_fd_sc_hd__a32o_2
XFILLER_129_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22728_ _22728_/CLK _22728_/D vssd1 vssd1 vccd1 vccd1 _22728_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13261__C _21724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16853__B _16853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13461_ _13461_/A _13461_/B vssd1 vssd1 vccd1 vccd1 _13461_/Y sky130_fd_sc_hd__nor2_1
X_22659_ _22659_/A vssd1 vssd1 vccd1 vccd1 _22949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ _15200_/A _15200_/B vssd1 vssd1 vccd1 vccd1 _15200_/X sky130_fd_sc_hd__xor2_1
XANTENNA__21693__A_N _21688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ _16328_/A vssd1 vssd1 vccd1 vccd1 _15369_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16180_ _15890_/X _15936_/X _15932_/X _16179_/X vssd1 vssd1 vccd1 vccd1 _16180_/X
+ sky130_fd_sc_hd__o22a_1
X_13392_ _13392_/A _13392_/B _13392_/C vssd1 vssd1 vccd1 vccd1 _13495_/A sky130_fd_sc_hd__nand3_2
XFILLER_12_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15131_ _15132_/B _15132_/A vssd1 vssd1 vccd1 vccd1 _15133_/A sky130_fd_sc_hd__nor2_1
XFILLER_154_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12343_ _12378_/A _12343_/B vssd1 vssd1 vccd1 vccd1 _12343_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15062_ _15062_/A _15114_/D _15114_/C _15070_/A vssd1 vssd1 vccd1 vccd1 _15062_/Y
+ sky130_fd_sc_hd__nand4_1
X_12274_ _22693_/Q vssd1 vssd1 vccd1 vccd1 _12300_/A sky130_fd_sc_hd__inv_2
XFILLER_4_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12714__A1 _12522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14013_ _14013_/A _14013_/B vssd1 vssd1 vccd1 vccd1 _14562_/A sky130_fd_sc_hd__nand2_1
XFILLER_49_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19870_ _19867_/X _19894_/A _19836_/D _19836_/Y vssd1 vssd1 vccd1 vccd1 _19921_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17102__B1 _17103_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12902__A _20130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17653__A1 _15941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18821_ _19651_/A _19334_/B _18664_/B _18666_/X vssd1 vssd1 vccd1 vccd1 _18826_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18752_ _18568_/A _18608_/Y _18568_/B vssd1 vssd1 vccd1 vccd1 _18753_/C sky130_fd_sc_hd__o21ai_1
X_15964_ _15964_/A _15964_/B vssd1 vssd1 vccd1 vccd1 _15964_/Y sky130_fd_sc_hd__nand2_2
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17703_ _17855_/A _17855_/B vssd1 vssd1 vccd1 vccd1 _17704_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__21201__A2 _21195_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14915_ _14916_/A _14916_/B _14916_/C _14916_/D vssd1 vssd1 vccd1 vccd1 _14919_/A
+ sky130_fd_sc_hd__a22o_1
X_18683_ _11415_/A _18855_/A _18682_/Y vssd1 vssd1 vccd1 vccd1 _18684_/A sky130_fd_sc_hd__o21ai_2
X_15895_ _15813_/Y _15900_/A _15778_/Y _15975_/B vssd1 vssd1 vccd1 vccd1 _15924_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__15416__B1 _15415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17634_ _17634_/A vssd1 vssd1 vccd1 vccd1 _17635_/A sky130_fd_sc_hd__buf_2
X_14846_ _14552_/X _14845_/C _14845_/A vssd1 vssd1 vccd1 vccd1 _14847_/B sky130_fd_sc_hd__o21ai_1
XFILLER_64_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17565_ _17427_/X _16737_/X _16276_/X _17091_/A vssd1 vssd1 vccd1 vccd1 _17565_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14777_ _15058_/A _15058_/B _14777_/C vssd1 vssd1 vccd1 vccd1 _14857_/B sky130_fd_sc_hd__and3_1
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11989_ _15776_/A vssd1 vssd1 vccd1 vccd1 _15893_/A sky130_fd_sc_hd__buf_4
XFILLER_95_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19304_ _19253_/Y _19255_/Y _19303_/Y vssd1 vssd1 vccd1 vccd1 _19304_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16516_ _18203_/C _12696_/X _16476_/X _16515_/Y _16479_/A vssd1 vssd1 vccd1 vccd1
+ _16517_/B sky130_fd_sc_hd__o221ai_1
XFILLER_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15719__A1 _11912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13728_ _13728_/A _14110_/B _14834_/C vssd1 vssd1 vccd1 vccd1 _14079_/A sky130_fd_sc_hd__and3_2
XFILLER_56_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17496_ _17375_/Y _17376_/Y _17495_/X vssd1 vssd1 vccd1 vccd1 _17726_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__15719__B2 _12009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19235_ _19400_/A _19244_/A _19246_/B vssd1 vssd1 vccd1 vccd1 _19396_/B sky130_fd_sc_hd__nand3_1
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16447_ _16447_/A _20323_/B vssd1 vssd1 vccd1 vccd1 _16816_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13659_ _13660_/A _13659_/B _13659_/C _21938_/B vssd1 vssd1 vccd1 vccd1 _13665_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19166_ _19168_/C vssd1 vssd1 vccd1 vccd1 _19461_/C sky130_fd_sc_hd__buf_2
XFILLER_118_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16378_ _16704_/A _16704_/B _16366_/Y _16374_/Y vssd1 vssd1 vccd1 vccd1 _16378_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_129_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18117_ _18126_/A _18128_/C _18319_/C vssd1 vssd1 vccd1 vccd1 _18690_/A sky130_fd_sc_hd__nand3_2
X_15329_ _15329_/A vssd1 vssd1 vccd1 vccd1 _15329_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17875__A _17875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19097_ _19104_/A _19254_/C _19097_/C vssd1 vssd1 vccd1 vccd1 _19097_/X sky130_fd_sc_hd__and3_1
XANTENNA__19793__C _19793_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18048_ _18048_/A _18048_/B _18048_/C vssd1 vssd1 vccd1 vccd1 _18048_/X sky130_fd_sc_hd__and3_1
XFILLER_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12705__A1 _12968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15395__A _20323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12705__B2 _12727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20779__A1 _15941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20010_ _20010_/A _20057_/B vssd1 vssd1 vccd1 vccd1 _20010_/X sky130_fd_sc_hd__or2b_1
XFILLER_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19999_ _20024_/A _19999_/B vssd1 vssd1 vccd1 vccd1 _19999_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16938__B _19490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21961_ _21376_/X _21958_/X _21960_/Y vssd1 vssd1 vccd1 vccd1 _21961_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20912_ _21009_/A _17733_/A _20919_/A vssd1 vssd1 vccd1 vccd1 _20916_/B sky130_fd_sc_hd__o21ai_1
XFILLER_27_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15958__A1 _15937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21892_ _21892_/A _21892_/B _21892_/C vssd1 vssd1 vccd1 vccd1 _21892_/Y sky130_fd_sc_hd__nand3_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13969__B1 _13968_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20843_ _20843_/A vssd1 vssd1 vccd1 vccd1 _20843_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_710 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19968__C _22924_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20774_ _20774_/A vssd1 vssd1 vccd1 vccd1 _22915_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__20703__A1 _12968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19687__D _19687_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18372__A2 _11351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13285__B1_N _13475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22513_ _22513_/A vssd1 vssd1 vccd1 vccd1 _22751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16922__A3 _16921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22444_ _22512_/S vssd1 vssd1 vccd1 vccd1 _22453_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__22456__A1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14394__B1 _14370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20786__A1_N _20210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22375_ _22375_/A vssd1 vssd1 vccd1 vccd1 _22689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21326_ _21324_/X _21325_/Y _21478_/A vssd1 vssd1 vccd1 vccd1 _21326_/X sky130_fd_sc_hd__o21a_1
XFILLER_159_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21257_ _21266_/B _21261_/B _21254_/X _21256_/Y vssd1 vssd1 vccd1 vccd1 _21257_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__13818__A _22868_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12172__A2 _12171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20208_ _16267_/X _16266_/X _20359_/B _16268_/X vssd1 vssd1 vccd1 vccd1 _20208_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_145_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21188_ _21188_/A _21188_/B _21188_/C vssd1 vssd1 vccd1 vccd1 _21188_/Y sky130_fd_sc_hd__nor3_1
XFILLER_89_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20139_ _20155_/B _20155_/C _20155_/A vssd1 vssd1 vccd1 vccd1 _20149_/C sky130_fd_sc_hd__nand3b_1
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12961_ _12997_/A _12963_/D vssd1 vssd1 vccd1 vccd1 _13003_/B sky130_fd_sc_hd__nand2_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _22765_/Q vssd1 vssd1 vccd1 vccd1 _14775_/D sky130_fd_sc_hd__inv_2
XFILLER_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _11912_/A vssd1 vssd1 vccd1 vccd1 _15936_/A sky130_fd_sc_hd__buf_4
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _15680_/A _15680_/B _15680_/C vssd1 vssd1 vccd1 vccd1 _15681_/D sky130_fd_sc_hd__nand3_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15471__C _15528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _20182_/A _20183_/A _20182_/B vssd1 vssd1 vccd1 vccd1 _12894_/A sky130_fd_sc_hd__a21oi_2
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _14622_/X _14635_/B _14635_/C vssd1 vssd1 vccd1 vccd1 _14631_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__20089__C _20341_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11843_ _12059_/B _12247_/B _11899_/A vssd1 vssd1 vccd1 vccd1 _11927_/A sky130_fd_sc_hd__a21o_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _17350_/A _17350_/B _17350_/C vssd1 vssd1 vccd1 vccd1 _17494_/A sky130_fd_sc_hd__nand3_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14562_ _14562_/A vssd1 vssd1 vccd1 vccd1 _14562_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _19197_/A _11949_/D vssd1 vssd1 vccd1 vccd1 _11774_/Y sky130_fd_sc_hd__nand2_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16296_/Y _16299_/Y _15797_/X _17443_/A vssd1 vssd1 vccd1 vccd1 _16301_/Y
+ sky130_fd_sc_hd__o2bb2ai_4
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13513_ _13513_/A _13513_/B _13521_/B _13519_/B vssd1 vssd1 vccd1 vccd1 _13515_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17281_ _18659_/D _17281_/B _20678_/B _18839_/B vssd1 vssd1 vccd1 vccd1 _17282_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14493_ _14491_/C _14963_/A _14963_/B _14486_/A _14494_/B vssd1 vssd1 vccd1 vccd1
+ _14500_/B sky130_fd_sc_hd__a32o_1
XFILLER_110_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19020_ _19026_/A _19020_/B vssd1 vssd1 vccd1 vccd1 _19022_/A sky130_fd_sc_hd__nand2_1
X_16232_ _16770_/A _16771_/A vssd1 vssd1 vccd1 vccd1 _17137_/A sky130_fd_sc_hd__nand2_1
XFILLER_110_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13444_ _13215_/A _13215_/B _13475_/B _13475_/C vssd1 vssd1 vccd1 vccd1 _13468_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__22447__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19312__A1 _19000_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12935__A1 _15804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16163_ _16169_/C _16111_/A _16111_/B vssd1 vssd1 vccd1 vccd1 _16163_/X sky130_fd_sc_hd__a21o_1
X_13375_ _13375_/A vssd1 vssd1 vccd1 vccd1 _21522_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15114_ _15114_/A _15114_/B _15114_/C _15114_/D vssd1 vssd1 vccd1 vccd1 _15119_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_155_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12326_ _12401_/A _12402_/A _12288_/A vssd1 vssd1 vccd1 vccd1 _12576_/A sky130_fd_sc_hd__a21oi_4
X_16094_ _16024_/A _16090_/B _16092_/Y _16093_/X vssd1 vssd1 vccd1 vccd1 _16094_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__21670__A2 _13162_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22106__A _22106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_997 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18303__B _18303_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19922_ _19922_/A _19922_/B vssd1 vssd1 vccd1 vccd1 _19922_/X sky130_fd_sc_hd__xor2_1
X_15045_ _15045_/A vssd1 vssd1 vccd1 vccd1 _22679_/D sky130_fd_sc_hd__clkbuf_1
X_12257_ _22909_/Q _12258_/A vssd1 vssd1 vccd1 vccd1 _18266_/A sky130_fd_sc_hd__nor2_1
XFILLER_107_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12632__A _15901_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19853_ _19909_/A _19909_/B _19851_/A _19851_/B vssd1 vssd1 vccd1 vccd1 _19853_/Y
+ sky130_fd_sc_hd__o211ai_2
X_12188_ _12188_/A _12188_/B _12188_/C vssd1 vssd1 vccd1 vccd1 _12225_/A sky130_fd_sc_hd__nand3_1
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18804_ _18804_/A _18804_/B vssd1 vssd1 vccd1 vccd1 _18804_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19784_ _19784_/A _19787_/B _19784_/C vssd1 vssd1 vccd1 vccd1 _19785_/C sky130_fd_sc_hd__nand3_1
X_16996_ _16996_/A vssd1 vssd1 vccd1 vccd1 _17313_/A sky130_fd_sc_hd__buf_2
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_bq_clk_i_A bq_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18735_ _18735_/A _18735_/B _18741_/C _18741_/D vssd1 vssd1 vccd1 vccd1 _18736_/C
+ sky130_fd_sc_hd__nand4_1
X_15947_ _15875_/B _15856_/Y _16024_/C _15946_/X vssd1 vssd1 vccd1 vccd1 _15947_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22383__A0 _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16477__C _16477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18666_ _19507_/A _18666_/B _18839_/B _19507_/D vssd1 vssd1 vccd1 vccd1 _18666_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15878_ _16209_/C _16208_/A _15951_/A _15877_/X vssd1 vssd1 vccd1 vccd1 _15879_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_37_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16601__A2 _16602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17617_ _17500_/Y _17501_/X _17616_/Y vssd1 vssd1 vccd1 vccd1 _17617_/Y sky130_fd_sc_hd__o21ai_1
X_14829_ _14828_/B _14828_/C _14764_/Y vssd1 vssd1 vccd1 vccd1 _14829_/X sky130_fd_sc_hd__a21bo_1
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18597_ _12250_/D _18236_/Y _18240_/Y _18772_/A vssd1 vssd1 vccd1 vccd1 _18598_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12218__A3 _19772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14612__A1 _13820_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12079__A _12079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17548_ _17731_/A _17388_/X _17382_/Y _17546_/X _17678_/A vssd1 vssd1 vccd1 vccd1
+ _17663_/B sky130_fd_sc_hd__o311a_1
XANTENNA__11426__A1 _18292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11977__A2 _15905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17479_ _17479_/A _17479_/B _17479_/C _17479_/D vssd1 vssd1 vccd1 vccd1 _17479_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17562__B1 _16016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14294__A _14843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11711__A _22959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19218_ _19218_/A _19218_/B vssd1 vssd1 vccd1 vccd1 _19227_/B sky130_fd_sc_hd__nand2_1
X_20490_ _20487_/X _20488_/X _20489_/Y vssd1 vssd1 vccd1 vccd1 _20490_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_146_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18106__A2 _12116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19149_ _19149_/A _19149_/B _19149_/C vssd1 vssd1 vccd1 vccd1 _19149_/X sky130_fd_sc_hd__and3_1
XFILLER_9_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17314__B1 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22160_ _22160_/A _22160_/B vssd1 vssd1 vccd1 vccd1 _22160_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21111_ _21088_/A _21088_/B _21091_/A vssd1 vssd1 vccd1 vccd1 _21112_/B sky130_fd_sc_hd__o21bai_2
XFILLER_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13638__A _21866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22091_ _22088_/Y _22284_/C _22145_/C vssd1 vssd1 vccd1 vccd1 _22092_/B sky130_fd_sc_hd__a21o_1
XFILLER_132_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16014__A _16014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21042_ _21008_/A _21008_/B _21031_/B vssd1 vssd1 vccd1 vccd1 _21062_/B sky130_fd_sc_hd__o21a_1
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18290__A1 _17636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17093__A2 _17083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22374__A0 _12528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21944_ _21944_/A vssd1 vssd1 vccd1 vccd1 _22122_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__20924__B2 _17922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21875_ _21875_/A _21875_/B _21875_/C vssd1 vssd1 vccd1 vccd1 _21882_/A sky130_fd_sc_hd__nand3_2
XFILLER_36_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22836__D _22848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20826_ _20830_/A _20830_/C _20830_/B vssd1 vssd1 vccd1 vccd1 _20840_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__12614__B1 _12602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20757_ _20758_/A _20830_/A _20759_/B _20759_/A vssd1 vssd1 vccd1 vccd1 _20761_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_11_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18107__C _18107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11490_ _18167_/A vssd1 vssd1 vccd1 vccd1 _18797_/C sky130_fd_sc_hd__buf_4
XFILLER_195_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20688_ _20793_/B vssd1 vssd1 vccd1 vccd1 _20936_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16108__A1 _16586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22427_ _22713_/Q input52/X _22435_/S vssd1 vssd1 vccd1 vccd1 _22428_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19845__A2 _20012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13590__A1 _21445_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15316__C1 _12003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13160_ _13456_/A vssd1 vssd1 vccd1 vccd1 _13504_/A sky130_fd_sc_hd__clkinv_2
XFILLER_151_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22358_ _22358_/A _22358_/B vssd1 vssd1 vccd1 vccd1 _22944_/D sky130_fd_sc_hd__nor2_1
XFILLER_191_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18123__B _19168_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12111_ _12111_/A vssd1 vssd1 vccd1 vccd1 _12111_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13091_ _21315_/B vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__clkbuf_2
X_21309_ _21738_/A _21476_/C _21739_/C vssd1 vssd1 vccd1 vccd1 _21482_/A sky130_fd_sc_hd__nand3_1
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22289_ _22684_/Q _22289_/B vssd1 vssd1 vccd1 vccd1 _22297_/B sky130_fd_sc_hd__nor2_1
XFILLER_156_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12042_ _16242_/A _22658_/B vssd1 vssd1 vccd1 vccd1 _12235_/B sky130_fd_sc_hd__nand2_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20663__A1_N _20827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20612__B1 _15939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18281__A1 _11859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16850_ _16734_/X _16735_/X _16849_/Y _16739_/Y vssd1 vssd1 vccd1 vccd1 _16853_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_133_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17084__A2 _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15801_ _15801_/A _15801_/B _15801_/C vssd1 vssd1 vccd1 vccd1 _15829_/A sky130_fd_sc_hd__nand3_1
XFILLER_19_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16781_ _20133_/A _16781_/B _18192_/A _18193_/A vssd1 vssd1 vccd1 vccd1 _16781_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_92_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13993_ _22866_/Q vssd1 vssd1 vccd1 vccd1 _14686_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_92_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18520_ _18520_/A _18520_/B vssd1 vssd1 vccd1 vccd1 _18726_/B sky130_fd_sc_hd__nand2_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _15427_/X _16039_/A _15406_/X _15404_/X _15403_/X vssd1 vssd1 vccd1 vccd1
+ _15733_/C sky130_fd_sc_hd__o221ai_4
X_12944_ _12705_/X _12737_/D _12942_/Y _12943_/X vssd1 vssd1 vccd1 vccd1 _12944_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20915__A1 _20123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18451_ _18451_/A _18451_/B vssd1 vssd1 vccd1 vccd1 _18451_/Y sky130_fd_sc_hd__nor2_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15663_ _15673_/B _16213_/A vssd1 vssd1 vccd1 vccd1 _15667_/A sky130_fd_sc_hd__nand2_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12875_ _12886_/B _12776_/A _16160_/C _20452_/C vssd1 vssd1 vccd1 vccd1 _12875_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17792__B1 _22901_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16594__A _16594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20391__A2 _16179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17402_ _15934_/A _17400_/X _17247_/X _17401_/Y vssd1 vssd1 vccd1 vccd1 _17402_/Y
+ sky130_fd_sc_hd__o22ai_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14614_ _13950_/X _13905_/Y _14619_/A _14503_/X vssd1 vssd1 vccd1 vccd1 _14614_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_60_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18382_ _18408_/C vssd1 vssd1 vccd1 vccd1 _18396_/C sky130_fd_sc_hd__buf_2
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _11811_/Y _11815_/Y _11761_/Y _11762_/X vssd1 vssd1 vccd1 vccd1 _11829_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__12605__B1 _12938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15594_ _15577_/X _15477_/B _15566_/X _15571_/Y _15574_/C vssd1 vssd1 vccd1 vccd1
+ _16286_/A sky130_fd_sc_hd__o2111ai_4
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_359 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17333_ _17486_/A _17486_/B _17333_/C _17333_/D vssd1 vssd1 vccd1 vccd1 _17333_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_144_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20679__B1 _20685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14561_/C _14044_/Y _14098_/B _14098_/A vssd1 vssd1 vccd1 vccd1 _14547_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_81_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11757_ _12062_/A _12165_/A _18133_/A vssd1 vssd1 vccd1 vccd1 _11757_/Y sky130_fd_sc_hd__nor3_1
XFILLER_18_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17264_ _16956_/Y _16949_/Y _17149_/B _17149_/A vssd1 vssd1 vccd1 vccd1 _17264_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_174_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14476_ _14693_/A vssd1 vssd1 vccd1 vccd1 _15069_/A sky130_fd_sc_hd__buf_2
XFILLER_146_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20844__A _20844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11688_ _11643_/Y _11649_/Y _11687_/Y vssd1 vssd1 vccd1 vccd1 _11842_/B sky130_fd_sc_hd__a21bo_1
X_19003_ _19179_/C _19007_/B _19001_/Y _19002_/Y vssd1 vssd1 vccd1 vccd1 _19086_/B
+ sky130_fd_sc_hd__o22ai_4
X_16215_ _16215_/A _16215_/B vssd1 vssd1 vccd1 vccd1 _16216_/B sky130_fd_sc_hd__nand2_1
XANTENNA__15938__A _15938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13427_ _13521_/A _21212_/C _13521_/C vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__nand3_1
X_17195_ _17027_/B _17027_/C _17187_/X vssd1 vssd1 vccd1 vccd1 _17197_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__15570__A2 _16039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15307__C1 _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16146_ _16141_/X _16140_/Y _16137_/Y _16132_/Y vssd1 vssd1 vccd1 vccd1 _16146_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_13358_ _13358_/A _13358_/B _13358_/C vssd1 vssd1 vccd1 vccd1 _13359_/A sky130_fd_sc_hd__nand3_1
XFILLER_142_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12309_ _12292_/A _12520_/B _12413_/A vssd1 vssd1 vccd1 vccd1 _12447_/A sky130_fd_sc_hd__a21o_1
XFILLER_142_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16077_ _15972_/X _16110_/B _16068_/Y _16055_/Y vssd1 vssd1 vccd1 vccd1 _16082_/A
+ sky130_fd_sc_hd__a22o_1
X_13289_ _13289_/A _13484_/B vssd1 vssd1 vccd1 vccd1 _13290_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19905_ _19905_/A _19937_/B _19905_/C _19939_/A vssd1 vssd1 vccd1 vccd1 _19907_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_170_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15028_ _15028_/A _15028_/B vssd1 vssd1 vccd1 vccd1 _15030_/C sky130_fd_sc_hd__nor2_1
XANTENNA__17872__B _21083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16807__C1 _18093_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13884__A2 _13851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19836_ _19836_/A _20012_/A _19836_/C _19836_/D vssd1 vssd1 vccd1 vccd1 _19836_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_122_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17591__C _20936_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16488__B _17139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15392__B _15665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19767_ _19695_/A _17822_/A _17817_/A _19176_/X vssd1 vssd1 vccd1 vccd1 _19836_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_7_1071 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16979_ _16978_/A _16978_/B _16939_/Y _16945_/X vssd1 vssd1 vccd1 vccd1 _16980_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__18984__A _18984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 wb_adr_i[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18718_ _19176_/A vssd1 vssd1 vccd1 vccd1 _18718_/X sky130_fd_sc_hd__buf_2
X_19698_ _19698_/A _19698_/B _19698_/C vssd1 vssd1 vccd1 vccd1 _19789_/A sky130_fd_sc_hd__nand3_1
XFILLER_80_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18649_ _12157_/X _12158_/X _17421_/A _17422_/A vssd1 vssd1 vccd1 vccd1 _18649_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15794__C1 _15834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21660_ _21650_/A _21650_/B _21650_/C _21659_/X vssd1 vssd1 vccd1 vccd1 _21660_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_52_668 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20611_ _20611_/A _20611_/B vssd1 vssd1 vccd1 vccd1 _20611_/Y sky130_fd_sc_hd__nand2_1
X_21591_ _21738_/A _21591_/B _22041_/C vssd1 vssd1 vccd1 vccd1 _21591_/Y sky130_fd_sc_hd__nand3_1
XFILLER_177_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12537__A _22823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11441__A _15714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20542_ _20545_/A _20420_/C _20426_/X _20427_/Y vssd1 vssd1 vccd1 vccd1 _20658_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_20_543 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20473_ _12734_/X _16745_/A _20495_/A vssd1 vssd1 vccd1 vccd1 _20599_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__15561__A2 _15569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22212_ _22212_/A _22212_/B _22212_/C vssd1 vssd1 vccd1 vccd1 _22212_/Y sky130_fd_sc_hd__nor3_1
XFILLER_118_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22143_ _22164_/A _22159_/B vssd1 vssd1 vccd1 vccd1 _22143_/X sky130_fd_sc_hd__and2_1
XFILLER_69_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22074_ _22072_/A _22072_/B _22068_/C _22068_/D vssd1 vssd1 vccd1 vccd1 _22074_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_102_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22595__A0 _11860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21025_ _21086_/C _17816_/B _20969_/A _20967_/Y vssd1 vssd1 vccd1 vccd1 _21027_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19460__B1 _11672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14199__A _14199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22822__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21927_ _22678_/Q _21927_/B _21927_/C vssd1 vssd1 vccd1 vccd1 _21927_/X sky130_fd_sc_hd__or3_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _15586_/C vssd1 vssd1 vccd1 vccd1 _15810_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__16041__A3 _20728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21858_ _21850_/Y _21852_/Y _21854_/X vssd1 vssd1 vccd1 vccd1 _21858_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11611_/A _11611_/B vssd1 vssd1 vccd1 vccd1 _18648_/D sky130_fd_sc_hd__nand2_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16329__A1 _16435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20809_ _20804_/Y _20884_/B _20808_/Y vssd1 vssd1 vccd1 vccd1 _20810_/C sky130_fd_sc_hd__a21oi_1
XFILLER_169_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12591_ _15631_/A _12493_/Y _12610_/A _20134_/A vssd1 vssd1 vccd1 vccd1 _12592_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_168_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21789_ _21847_/B _21789_/B vssd1 vssd1 vccd1 vccd1 _21789_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ _14361_/A vssd1 vssd1 vccd1 vccd1 _14330_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_196_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11542_ _11542_/A vssd1 vssd1 vccd1 vccd1 _18371_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20086__D _20456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14261_ _14272_/A _14261_/B _14261_/C vssd1 vssd1 vccd1 vccd1 _14269_/A sky130_fd_sc_hd__nand3b_1
X_11473_ _18093_/A _18093_/B vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__nand2_2
XANTENNA__18134__A _18690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16000_ _16000_/A _16000_/B _16000_/C vssd1 vssd1 vccd1 vccd1 _16046_/A sky130_fd_sc_hd__nand3_1
XANTENNA_input70_A x[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13212_ _21398_/A _13517_/A vssd1 vssd1 vccd1 vccd1 _13434_/A sky130_fd_sc_hd__nand2_1
XFILLER_136_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14192_ _14510_/C _14210_/A _14911_/C _14191_/B _14489_/C vssd1 vssd1 vccd1 vccd1
+ _14195_/A sky130_fd_sc_hd__a32o_1
XFILLER_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13143_ _13143_/A _13143_/B vssd1 vssd1 vccd1 vccd1 _13144_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17951_ _17949_/A _17919_/C _17950_/A vssd1 vssd1 vccd1 vccd1 _17957_/B sky130_fd_sc_hd__o21a_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _21213_/A _13519_/B _21214_/A vssd1 vssd1 vccd1 vccd1 _13120_/B sky130_fd_sc_hd__nand3_2
X_16902_ _22893_/Q _16702_/Y _16899_/Y _17070_/A _16901_/Y vssd1 vssd1 vccd1 vccd1
+ _16905_/A sky130_fd_sc_hd__o2111a_1
XANTENNA__15493__A _19197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12025_ _12025_/A _12025_/B _12025_/C vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__nand3_2
X_17882_ _17882_/A _19896_/B _17882_/C vssd1 vssd1 vccd1 vccd1 _17883_/D sky130_fd_sc_hd__and3_1
XFILLER_120_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19621_ _19985_/C _19621_/B _19621_/C _19793_/C vssd1 vssd1 vccd1 vccd1 _19621_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_120_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_727 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16833_ _16906_/A _16906_/B _16906_/C vssd1 vssd1 vccd1 vccd1 _16866_/B sky130_fd_sc_hd__nand3_2
XFILLER_120_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15473__D1 _17246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__A1 _11625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19552_ _19552_/A _19552_/B _19552_/C vssd1 vssd1 vccd1 vccd1 _19552_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__19203__B1 _19211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764_ _15546_/X _16758_/X _16773_/A vssd1 vssd1 vccd1 vccd1 _16768_/A sky130_fd_sc_hd__o21ai_2
XFILLER_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13976_ _14475_/A _14475_/B _13975_/Y vssd1 vssd1 vccd1 vccd1 _14002_/C sky130_fd_sc_hd__a21o_2
XANTENNA__16017__B1 _16016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21010__B1 _20514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15715_ _16554_/C _16191_/A _15775_/B _15714_/X vssd1 vssd1 vccd1 vccd1 _15752_/A
+ sky130_fd_sc_hd__a31o_1
X_18503_ _18698_/B _18678_/D vssd1 vssd1 vccd1 vccd1 _18876_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12927_ _12772_/X _12774_/X _12689_/X _12712_/Y _20793_/B vssd1 vssd1 vccd1 vccd1
+ _12927_/X sky130_fd_sc_hd__o221a_1
X_19483_ _19630_/A _19630_/C _19630_/D vssd1 vssd1 vccd1 vccd1 _19636_/B sky130_fd_sc_hd__nand3_2
X_16695_ _22890_/Q _22889_/Q _16695_/C _16695_/D vssd1 vssd1 vccd1 vccd1 _16695_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18434_ _18434_/A _18434_/B vssd1 vssd1 vccd1 vccd1 _18435_/B sky130_fd_sc_hd__nand2_1
X_15646_ _15646_/A vssd1 vssd1 vccd1 vccd1 _15646_/X sky130_fd_sc_hd__buf_4
XFILLER_61_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12858_ _12863_/A _12863_/B _12843_/X _12851_/Y _12862_/B vssd1 vssd1 vccd1 vccd1
+ _12867_/A sky130_fd_sc_hd__o221ai_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19506__A1 _12170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18365_ _18365_/A _18995_/A vssd1 vssd1 vccd1 vccd1 _18365_/Y sky130_fd_sc_hd__nor2_1
X_11809_ _11809_/A _11809_/B vssd1 vssd1 vccd1 vccd1 _11814_/B sky130_fd_sc_hd__nor2_1
X_15577_ _19012_/D _17672_/A _20390_/C _15577_/D vssd1 vssd1 vccd1 vccd1 _15577_/X
+ sky130_fd_sc_hd__and4_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12789_/A vssd1 vssd1 vccd1 vccd1 _20241_/A sky130_fd_sc_hd__buf_2
XFILLER_109_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17081_/A _17591_/B _17085_/Y vssd1 vssd1 vccd1 vccd1 _17520_/D sky130_fd_sc_hd__o21ai_4
XFILLER_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11801__A1 _11800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14528_ _13937_/C _13937_/D _13947_/A vssd1 vssd1 vccd1 vccd1 _14528_/Y sky130_fd_sc_hd__a21oi_2
X_18296_ _18296_/A _18296_/B vssd1 vssd1 vccd1 vccd1 _18296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17247_ _17247_/A vssd1 vssd1 vccd1 vccd1 _17247_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14459_ _14103_/B _14103_/A _14103_/C vssd1 vssd1 vccd1 vccd1 _14661_/C sky130_fd_sc_hd__a21bo_4
XFILLER_179_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18044__A _18044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17178_ _17178_/A _17178_/B vssd1 vssd1 vccd1 vccd1 _17178_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16129_ _16129_/A _20390_/C _16129_/C _16192_/D vssd1 vssd1 vccd1 vccd1 _16131_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_6_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12109__A2 _18510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22845__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15059__A1 _14503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18796__A2 _15545_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19819_ _18246_/A _18246_/B _19761_/Y _19880_/C vssd1 vssd1 vccd1 vccd1 _19822_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13635__B _21878_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16011__B _16011_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22830_ _22850_/CLK _22842_/Q vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_602 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19322__B _19322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16559__A1 _15797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22761_ _22761_/CLK _22761_/D vssd1 vssd1 vccd1 vccd1 _22761_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21712_ _21815_/B _21702_/B _21574_/A _21707_/B vssd1 vssd1 vccd1 vccd1 _21821_/A
+ sky130_fd_sc_hd__a211o_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22692_ _22693_/CLK _22692_/D vssd1 vssd1 vccd1 vccd1 _22692_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12575__A1_N _16947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21643_ _21636_/X _21654_/C _21642_/Y vssd1 vssd1 vccd1 vccd1 _21662_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21574_ _21574_/A _21707_/B vssd1 vssd1 vccd1 vccd1 _21834_/A sky130_fd_sc_hd__nor2_1
XFILLER_123_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20525_ _20491_/Y _20501_/X _20623_/A _20623_/B vssd1 vssd1 vccd1 vccd1 _20526_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_122_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16731__A1 _16564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16731__B2 _16106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_676 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20456_ _20477_/A _20456_/B _20456_/C _20576_/B vssd1 vssd1 vccd1 vccd1 _20456_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_174_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18889__A _19316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17793__A _22901_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20387_ _20362_/Y _20367_/Y _20337_/A _20403_/B vssd1 vssd1 vccd1 vccd1 _20388_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15298__A1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15298__B2 _15808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22126_ _22129_/A _22129_/B _22124_/Y _22125_/X vssd1 vssd1 vccd1 vccd1 _22135_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_122_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22057_ _22182_/A _22057_/B _22182_/C vssd1 vssd1 vccd1 vccd1 _22190_/D sky130_fd_sc_hd__and3_1
XANTENNA__22032__A2 _21522_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19984__A1 _19419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21008_ _21008_/A _21008_/B vssd1 vssd1 vccd1 vccd1 _21008_/X sky130_fd_sc_hd__or2_1
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16798__A1 _15840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13830_ _13819_/Y _13824_/X _13829_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_29_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13761_ _13766_/B _13761_/B vssd1 vssd1 vccd1 vccd1 _13949_/A sky130_fd_sc_hd__nand2_2
X_22959_ _22959_/CLK _22959_/D vssd1 vssd1 vccd1 vccd1 _22959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15500_ _15500_/A _15500_/B vssd1 vssd1 vccd1 vccd1 _15596_/A sky130_fd_sc_hd__nor2_1
XFILLER_71_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12712_ _12689_/A _17401_/B _12711_/X _12681_/X vssd1 vssd1 vccd1 vccd1 _12712_/Y
+ sky130_fd_sc_hd__a31oi_2
X_16480_ _15504_/X _17379_/A _16476_/X _16513_/A _16479_/X vssd1 vssd1 vccd1 vccd1
+ _16480_/X sky130_fd_sc_hd__o311a_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _13776_/B vssd1 vssd1 vccd1 vccd1 _14199_/A sky130_fd_sc_hd__buf_2
XFILLER_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15431_ _15707_/B _15700_/C vssd1 vssd1 vccd1 vccd1 _15431_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12643_ _12745_/B _12643_/B vssd1 vssd1 vccd1 vccd1 _12755_/B sky130_fd_sc_hd__nand2_1
XFILLER_169_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18150_ _18150_/A _18150_/B vssd1 vssd1 vccd1 vccd1 _18389_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15362_ _16323_/A _16323_/B _16323_/C _15362_/D vssd1 vssd1 vccd1 vccd1 _15369_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_157_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12574_ _12574_/A vssd1 vssd1 vccd1 vccd1 _12988_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_169_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17101_ _17001_/C _17001_/A _17001_/B _17006_/C _16727_/X vssd1 vssd1 vccd1 vccd1
+ _17103_/C sky130_fd_sc_hd__a32o_2
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14313_ _14351_/A vssd1 vssd1 vccd1 vccd1 _14313_/X sky130_fd_sc_hd__clkbuf_2
X_18081_ _18077_/A _18057_/B _18079_/A vssd1 vssd1 vccd1 vccd1 _18081_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_183_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11525_ _18482_/A _18482_/B vssd1 vssd1 vccd1 vccd1 _11526_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15525__A2 _12211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15293_ _22884_/Q _22885_/Q _15288_/A _22888_/Q vssd1 vssd1 vccd1 vccd1 _15294_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__12905__A _20133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17032_ _16873_/C _16858_/A _16856_/Y vssd1 vssd1 vccd1 vccd1 _17033_/C sky130_fd_sc_hd__a21oi_1
XFILLER_183_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14244_ _14253_/A _14246_/A _14246_/B vssd1 vssd1 vccd1 vccd1 _14245_/B sky130_fd_sc_hd__a21bo_1
X_11456_ _11727_/C _11407_/B _15435_/B vssd1 vssd1 vccd1 vccd1 _11504_/A sky130_fd_sc_hd__a21o_1
XFILLER_7_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17278__A2 _16708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14175_ _14172_/A _14175_/B _14175_/C vssd1 vssd1 vccd1 vccd1 _14285_/B sky130_fd_sc_hd__nand3b_1
XFILLER_139_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11387_ _11411_/A vssd1 vssd1 vccd1 vccd1 _11727_/C sky130_fd_sc_hd__buf_2
XANTENNA__22868__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13126_ _13126_/A vssd1 vssd1 vccd1 vccd1 _13126_/X sky130_fd_sc_hd__clkbuf_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _18983_/A vssd1 vssd1 vccd1 vccd1 _19156_/D sky130_fd_sc_hd__buf_2
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17934_ _17928_/X _17885_/A _17932_/Y vssd1 vssd1 vccd1 vccd1 _17974_/A sky130_fd_sc_hd__a21oi_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13067_/A _13067_/B _13057_/C _13112_/C vssd1 vssd1 vccd1 vccd1 _13096_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_87_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12008_ _12008_/A vssd1 vssd1 vccd1 vccd1 _12009_/A sky130_fd_sc_hd__clkbuf_4
X_17865_ _17850_/Y _17851_/X _17864_/Y vssd1 vssd1 vccd1 vccd1 _18007_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__16789__A1 _17636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater128 _22875_/Q vssd1 vssd1 vccd1 vccd1 _22863_/D sky130_fd_sc_hd__buf_2
Xrepeater139 _22761_/CLK vssd1 vssd1 vccd1 vccd1 _22791_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
X_19604_ _19591_/Y _19594_/Y _19598_/Y _19602_/Y _19603_/X vssd1 vssd1 vccd1 vccd1
+ _19605_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16816_ _16816_/A _16911_/A vssd1 vssd1 vccd1 vccd1 _16816_/Y sky130_fd_sc_hd__nor2_1
X_17796_ _17795_/A _17795_/B _17795_/C vssd1 vssd1 vccd1 vccd1 _18007_/A sky130_fd_sc_hd__a21oi_4
XFILLER_19_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19727__A1 _19605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19535_ _19510_/Y _19513_/Y _19538_/C _19538_/A vssd1 vssd1 vccd1 vccd1 _19536_/D
+ sky130_fd_sc_hd__o211ai_2
XFILLER_35_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16747_ _15932_/X _16746_/X _16727_/X _16732_/B vssd1 vssd1 vccd1 vccd1 _16747_/X
+ sky130_fd_sc_hd__o31a_1
X_13959_ _13959_/A vssd1 vssd1 vccd1 vccd1 _14510_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16678_ _15881_/Y _16212_/Y _16406_/Y vssd1 vssd1 vccd1 vccd1 _16683_/B sky130_fd_sc_hd__o21ai_1
X_19466_ _14432_/A _15808_/X _11672_/X _19694_/D _19465_/Y vssd1 vssd1 vccd1 vccd1
+ _19466_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18417_ _18417_/A _18417_/B _18417_/C vssd1 vssd1 vccd1 vccd1 _18417_/Y sky130_fd_sc_hd__nand3_1
XFILLER_179_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15629_ _16563_/A _16563_/B vssd1 vssd1 vccd1 vccd1 _16361_/A sky130_fd_sc_hd__and2_1
X_19397_ _19239_/X _19242_/Y _19396_/Y vssd1 vssd1 vccd1 vccd1 _19399_/B sky130_fd_sc_hd__o21ai_1
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18348_ _18348_/A _19165_/A _18483_/B vssd1 vssd1 vccd1 vccd1 _18349_/B sky130_fd_sc_hd__and3_1
XFILLER_159_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_660 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16932__D _20502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18279_ _18279_/A _18279_/B vssd1 vssd1 vccd1 vccd1 _18572_/C sky130_fd_sc_hd__nand2_1
XFILLER_190_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20310_ _20553_/A _20553_/B _20309_/A _20314_/B vssd1 vssd1 vccd1 vccd1 _20311_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput50 wb_dat_i[23] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
X_21290_ _21294_/B _21558_/A _21288_/Y _21289_/Y vssd1 vssd1 vccd1 vccd1 _21292_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_162_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput61 wb_dat_i[4] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_4
Xinput72 x[1] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20241_ _20241_/A vssd1 vssd1 vccd1 vccd1 _20685_/A sky130_fd_sc_hd__buf_2
XFILLER_162_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20751__B _20751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20172_ _12886_/A _12878_/X _12781_/B _20165_/Y _20181_/B vssd1 vssd1 vccd1 vccd1
+ _20174_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17118__A _20781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12502__A2 _12501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19333__A _19687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18875__C _18875_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_760 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19718__B2 _19719_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22813_ _22813_/CLK _22813_/D vssd1 vssd1 vccd1 vccd1 _22813_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19052__B _19694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17729__B1 _17442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22744_ _22744_/CLK _22744_/D vssd1 vssd1 vccd1 vccd1 _22744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16952__A1 _15546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22675_ _22948_/CLK _22675_/D vssd1 vssd1 vccd1 vccd1 _22675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16952__B2 _18814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12428__C _20359_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21626_ _21493_/Y _21610_/A _21499_/X vssd1 vssd1 vccd1 vccd1 _21716_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__21828__A2 _22674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18154__B1 _15981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15507__A2 _12735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21557_ _21560_/A _21576_/A _21838_/A _21556_/Y vssd1 vssd1 vccd1 vccd1 _21566_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ _22956_/Q vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__buf_4
XFILLER_166_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20508_ _20508_/A vssd1 vssd1 vccd1 vccd1 _20913_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12290_ _22693_/Q _22692_/Q vssd1 vssd1 vccd1 vccd1 _12822_/A sky130_fd_sc_hd__nor2_4
XFILLER_153_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16180__A2 _15936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21488_ _21478_/X _21874_/C _21874_/A _21872_/A _21482_/Y vssd1 vssd1 vccd1 vccd1
+ _21488_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_153_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20439_ _20439_/A _20439_/B _22932_/Q vssd1 vssd1 vccd1 vccd1 _20562_/C sky130_fd_sc_hd__nand3_1
XFILLER_106_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16468__B1 _16842_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12163__C _15714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21476__C _21476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18131__B _18131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22109_ _21376_/X _21594_/Y _22108_/Y vssd1 vssd1 vccd1 vccd1 _22109_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_121_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15980_ _15797_/X _15890_/A _15780_/B _15901_/Y _15900_/Y vssd1 vssd1 vccd1 vccd1
+ _16045_/B sky130_fd_sc_hd__o221ai_4
XFILLER_110_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15691__A1 _14431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14931_ _14880_/A _14880_/B _14877_/C _14887_/C vssd1 vssd1 vccd1 vccd1 _14947_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_130_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18090__C1 _11666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17650_ _17645_/Y _17648_/Y _17649_/X vssd1 vssd1 vccd1 vccd1 _17654_/B sky130_fd_sc_hd__a21bo_1
X_14862_ _14862_/A _14932_/A vssd1 vssd1 vccd1 vccd1 _14862_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16586__B _16586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17983__A3 _19945_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16601_ _16602_/A _16602_/B _16602_/C _16600_/X vssd1 vssd1 vccd1 vccd1 _16601_/Y
+ sky130_fd_sc_hd__a31oi_1
X_13813_ _13826_/A _13826_/B _13826_/C vssd1 vssd1 vccd1 vccd1 _13814_/B sky130_fd_sc_hd__a21bo_2
XFILLER_180_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17581_ _17627_/A _17581_/B _17628_/A vssd1 vssd1 vccd1 vccd1 _17581_/Y sky130_fd_sc_hd__nand3_1
X_14793_ _14793_/A _14793_/B vssd1 vssd1 vccd1 vccd1 _14793_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16532_ _16532_/A _16532_/B vssd1 vssd1 vccd1 vccd1 _16532_/Y sky130_fd_sc_hd__nand2_1
X_19320_ _19320_/A _19490_/C _19490_/D vssd1 vssd1 vccd1 vccd1 _19320_/X sky130_fd_sc_hd__and3_1
XFILLER_73_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13744_ _13773_/A vssd1 vssd1 vccd1 vccd1 _13745_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19590__C1 _18718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19251_ _19239_/X _19242_/Y _19396_/C _19238_/A vssd1 vssd1 vccd1 vccd1 _19251_/Y
+ sky130_fd_sc_hd__o211ai_4
X_16463_ _16463_/A _16463_/B _16463_/C vssd1 vssd1 vccd1 vccd1 _16469_/B sky130_fd_sc_hd__nand3_1
X_13675_ _13677_/A _13677_/B _13677_/C vssd1 vssd1 vccd1 vccd1 _13678_/A sky130_fd_sc_hd__a21o_1
X_18202_ _18571_/B _18571_/C vssd1 vssd1 vccd1 vccd1 _18402_/B sky130_fd_sc_hd__nand2_1
X_15414_ _20092_/B vssd1 vssd1 vccd1 vccd1 _20675_/B sky130_fd_sc_hd__buf_2
XFILLER_19_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19182_ _19190_/A _19190_/B _19182_/C vssd1 vssd1 vccd1 vccd1 _19240_/D sky130_fd_sc_hd__nand3_2
Xclkbuf_0_bq_clk_i bq_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_bq_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_12626_ _20134_/C vssd1 vssd1 vccd1 vccd1 _20502_/C sky130_fd_sc_hd__clkbuf_2
X_16394_ _20793_/C vssd1 vssd1 vccd1 vccd1 _20917_/B sky130_fd_sc_hd__buf_2
XANTENNA__18145__B1 _18896_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14834__B _15186_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18306__B _18572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18133_ _18133_/A vssd1 vssd1 vccd1 vccd1 _18365_/A sky130_fd_sc_hd__clkbuf_2
X_15345_ _15331_/Y _15329_/A _15426_/B _15344_/X vssd1 vssd1 vccd1 vccd1 _15345_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_8_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12557_ _12557_/A _12557_/B _16486_/C _20134_/C vssd1 vssd1 vccd1 vccd1 _12628_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__22690__CLK _22690_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18064_ _17946_/A _17996_/A _18036_/B _18035_/B _18033_/A vssd1 vssd1 vccd1 vccd1
+ _18065_/C sky130_fd_sc_hd__o32a_1
XANTENNA__13509__B2 _22108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11508_ _11493_/Y _11501_/Y _11507_/X vssd1 vssd1 vccd1 vccd1 _11551_/B sky130_fd_sc_hd__a21bo_1
X_15276_ _22876_/D vssd1 vssd1 vccd1 vccd1 _15288_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12488_ _12417_/X _12425_/X _12346_/Y _12357_/Y vssd1 vssd1 vccd1 vccd1 _12488_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17015_ _17006_/Y _17008_/Y _17010_/X vssd1 vssd1 vccd1 vccd1 _17025_/B sky130_fd_sc_hd__a21o_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18448__A1 _17381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14227_ _15114_/D vssd1 vssd1 vccd1 vccd1 _15154_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__19418__A _19418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11439_ _14429_/A _11435_/X _11438_/Y vssd1 vssd1 vccd1 vccd1 _15633_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__21047__A3 _17839_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14182__B2 _13924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14158_ _14230_/A vssd1 vssd1 vccd1 vccd1 _14857_/A sky130_fd_sc_hd__buf_2
XFILLER_113_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13109_ _22724_/Q vssd1 vssd1 vccd1 vccd1 _13112_/D sky130_fd_sc_hd__inv_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ _18967_/B _22914_/Q vssd1 vssd1 vccd1 vccd1 _18968_/A sky130_fd_sc_hd__nand2_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _14167_/A _14167_/B _14167_/C vssd1 vssd1 vccd1 vccd1 _14089_/Y sky130_fd_sc_hd__a21oi_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21683__A _21683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17917_ _17866_/A _18007_/A _17864_/Y _17851_/X _17850_/Y vssd1 vssd1 vccd1 vccd1
+ _17918_/B sky130_fd_sc_hd__o32ai_4
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12496__A1 _15631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18897_ _18897_/A vssd1 vssd1 vccd1 vccd1 _19009_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18620__A1 _12064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17848_ _17775_/X _17799_/B _17860_/B vssd1 vssd1 vccd1 vccd1 _17848_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_187_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17779_ _17625_/A _17625_/B _17702_/A _17702_/B _17778_/Y vssd1 vssd1 vccd1 vccd1
+ _17779_/X sky130_fd_sc_hd__a41o_1
XANTENNA__14297__A input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19518_ _17083_/X _18980_/C _19981_/A _19321_/Y _19324_/X vssd1 vssd1 vccd1 vccd1
+ _19518_/X sky130_fd_sc_hd__o32a_1
XFILLER_35_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20790_ _16579_/X _16580_/X _20793_/A _17462_/A vssd1 vssd1 vccd1 vccd1 _20790_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19449_ _19449_/A _19449_/B _22917_/Q vssd1 vssd1 vccd1 vccd1 _19449_/Y sky130_fd_sc_hd__nand3_1
XFILLER_179_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17401__A _17401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22460_ _13095_/X input64/X _22464_/S vssd1 vssd1 vccd1 vccd1 _22461_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21411_ _21411_/A vssd1 vssd1 vccd1 vccd1 _21553_/A sky130_fd_sc_hd__buf_2
XFILLER_176_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22391_ _12378_/C input66/X _22391_/S vssd1 vssd1 vccd1 vccd1 _22392_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20494__A1 _12697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21342_ _21348_/A _21344_/D _21767_/A _21341_/X vssd1 vssd1 vccd1 vccd1 _21342_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__21691__B1 _21809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21273_ _21257_/Y _21261_/Y _21263_/Y vssd1 vssd1 vccd1 vccd1 _21281_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20481__B _20579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20246__A1 _20685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20224_ _20224_/A _20224_/B _20224_/C vssd1 vssd1 vccd1 vccd1 _20236_/B sky130_fd_sc_hd__nand3_4
XANTENNA__19047__B _19047_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11931__B1 _11762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20155_ _20155_/A _20155_/B _20155_/C vssd1 vssd1 vccd1 vccd1 _20155_/X sky130_fd_sc_hd__and3_1
XFILLER_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13807__C _14892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13133__C1 _13055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20086_ _20086_/A _20323_/B _20463_/C _20456_/C vssd1 vssd1 vccd1 vccd1 _20086_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17414__A2 _17388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18611__A1 _12170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14228__A2 _15154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19167__A2 _15808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11792_/A _11792_/B _11790_/C vssd1 vssd1 vccd1 vccd1 _11969_/A sky130_fd_sc_hd__nand3_2
XANTENNA__20706__C1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20988_ _21008_/A _21008_/B vssd1 vssd1 vccd1 vccd1 _20992_/C sky130_fd_sc_hd__xor2_1
XANTENNA__11998__B1 _15893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22727_ _22728_/CLK _22727_/D vssd1 vssd1 vccd1 vccd1 _22727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13460_ _13460_/A _13460_/B vssd1 vssd1 vccd1 vccd1 _13537_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22658_ _22658_/A _22658_/B vssd1 vssd1 vccd1 vccd1 _22659_/A sky130_fd_sc_hd__and2_1
XFILLER_139_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19885__A_N _22922_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12411_ _12411_/A vssd1 vssd1 vccd1 vccd1 _12967_/A sky130_fd_sc_hd__buf_2
X_21609_ _21609_/A _21609_/B _22229_/C vssd1 vssd1 vccd1 vccd1 _21610_/B sky130_fd_sc_hd__nand3_2
XFILLER_51_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13391_ _13391_/A _13391_/B vssd1 vssd1 vccd1 vccd1 _13392_/C sky130_fd_sc_hd__nand2_1
X_22589_ _18953_/C input35/X _22597_/S vssd1 vssd1 vccd1 vccd1 _22590_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16689__B1 _22891_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15130_ _15145_/A _15145_/B vssd1 vssd1 vccd1 vccd1 _15132_/A sky130_fd_sc_hd__xnor2_1
XFILLER_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21682__B1 _21687_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12342_ _12361_/A vssd1 vssd1 vccd1 vccd1 _12343_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_193_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15061_ _15061_/A vssd1 vssd1 vccd1 vccd1 _15119_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_107_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12273_ _12387_/A _12273_/B _12300_/B vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__nand3_2
XFILLER_182_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14670__A _14670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20237__A1 _20678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14012_ _14034_/A _14034_/B _14035_/A _14523_/A vssd1 vssd1 vccd1 vccd1 _14031_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13911__A1 _13814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12714__A2 _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17981__A _21044_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18820_ _19061_/A vssd1 vssd1 vccd1 vccd1 _19651_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13286__A _13340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17653__A2 _17822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22599__A _22656_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18751_ _18725_/X _18732_/Y _18737_/X _18748_/B vssd1 vssd1 vccd1 vccd1 _18753_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15963_ _15949_/A _15947_/Y _15959_/X _15962_/X vssd1 vssd1 vccd1 vccd1 _15964_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__13436__D _21739_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17702_ _17702_/A _17702_/B vssd1 vssd1 vccd1 vccd1 _17855_/B sky130_fd_sc_hd__nand2_2
X_14914_ _14972_/A _14972_/B _14914_/C vssd1 vssd1 vccd1 vccd1 _14916_/D sky130_fd_sc_hd__or3_1
XFILLER_64_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15894_ _15890_/X _16098_/A _15900_/B _15900_/A vssd1 vssd1 vccd1 vccd1 _15894_/X
+ sky130_fd_sc_hd__o22a_1
X_18682_ _18857_/A _18858_/A _18682_/C vssd1 vssd1 vccd1 vccd1 _18682_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__15416__A1 _15932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17633_ _19844_/D _17882_/C _17833_/A _19774_/D vssd1 vssd1 vccd1 vccd1 _17633_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14845_ _14845_/A _14845_/B _14845_/C vssd1 vssd1 vccd1 vccd1 _14847_/A sky130_fd_sc_hd__or3_1
XFILLER_91_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11534__A _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15006__A _15006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_510 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17564_ _17564_/A _17564_/B vssd1 vssd1 vccd1 vccd1 _17564_/Y sky130_fd_sc_hd__nor2_1
X_14776_ _14869_/A _22766_/Q _14869_/B vssd1 vssd1 vccd1 vccd1 _14858_/A sky130_fd_sc_hd__nand3_2
XFILLER_16_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11988_ _11988_/A vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__buf_4
X_19303_ _19303_/A _19303_/B vssd1 vssd1 vccd1 vccd1 _19303_/Y sky130_fd_sc_hd__nand2_1
X_16515_ _16515_/A _18192_/A _18193_/A vssd1 vssd1 vccd1 vccd1 _16515_/Y sky130_fd_sc_hd__nand3_2
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13727_ _13727_/A vssd1 vssd1 vccd1 vccd1 _14834_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_44_593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17495_ _17497_/A _17497_/B vssd1 vssd1 vccd1 vccd1 _17495_/X sky130_fd_sc_hd__and2_1
XANTENNA__15719__A2 _15723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14845__A _14845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17221__A _22895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19234_ _19246_/A _19400_/B vssd1 vssd1 vccd1 vccd1 _19396_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16446_ _15589_/X _16474_/A _16247_/B _16221_/Y vssd1 vssd1 vccd1 vccd1 _16734_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_13658_ _13658_/A _13658_/B _13658_/C vssd1 vssd1 vccd1 vccd1 _13659_/B sky130_fd_sc_hd__nand3_1
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _20461_/C vssd1 vssd1 vccd1 vccd1 _12973_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16377_ _16377_/A _16377_/B _16377_/C vssd1 vssd1 vccd1 vccd1 _16704_/B sky130_fd_sc_hd__nand3_1
XANTENNA__18669__A1 _17427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19165_ _19165_/A vssd1 vssd1 vccd1 vccd1 _19461_/B sky130_fd_sc_hd__clkbuf_4
X_13589_ _13576_/X _13578_/X _13587_/Y _13588_/X vssd1 vssd1 vccd1 vccd1 _13589_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_118_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20476__A1 _20579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15328_ _12090_/C _12921_/A _15327_/Y vssd1 vssd1 vccd1 vccd1 _15344_/A sky130_fd_sc_hd__o21ai_1
X_18116_ _18116_/A _18116_/B _18677_/A _18116_/D vssd1 vssd1 vccd1 vccd1 _18126_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__20476__B2 _16304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12953__A2 _16100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19096_ _19096_/A vssd1 vssd1 vccd1 vccd1 _19254_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_118_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18047_ _18049_/A _18049_/B _18046_/Y vssd1 vssd1 vccd1 vccd1 _18069_/C sky130_fd_sc_hd__o21ai_2
X_15259_ _15259_/A _15259_/B _15259_/C vssd1 vssd1 vccd1 vccd1 _15260_/B sky130_fd_sc_hd__nor3_2
XFILLER_126_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12705__A2 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20779__A2 _20123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11709__A _16257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19998_ _19998_/A _19998_/B vssd1 vssd1 vccd1 vccd1 _19999_/B sky130_fd_sc_hd__or2_1
XFILLER_113_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18949_ _18945_/A _18945_/B _18945_/C _18952_/C vssd1 vssd1 vccd1 vccd1 _18950_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_101_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12250__D _12250_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16938__C _19490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13924__A _13924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21960_ _21185_/X _21187_/X _22182_/B _22229_/A vssd1 vssd1 vccd1 vccd1 _21960_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__16300__A _16300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20911_ _20123_/X _17440_/A _17460_/A _20910_/Y vssd1 vssd1 vccd1 vccd1 _20919_/A
+ sky130_fd_sc_hd__o31ai_1
XFILLER_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15958__A2 _15942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21891_ _21891_/A _21891_/B vssd1 vssd1 vccd1 vccd1 _21892_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_655 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11444__A _19061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13969__A1 _13904_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20842_ _20890_/B _20830_/A _20890_/C vssd1 vssd1 vccd1 vccd1 _20842_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__14630__A2 _14512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20773_ _20773_/A _20773_/B vssd1 vssd1 vccd1 vccd1 _20774_/A sky130_fd_sc_hd__and2_1
XANTENNA__20703__A2 _16746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17131__A _19587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18372__A3 _16276_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22512_ _22751_/Q input59/X _22512_/S vssd1 vssd1 vccd1 vccd1 _22513_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22443_ _22499_/A vssd1 vssd1 vccd1 vccd1 _22512_/S sky130_fd_sc_hd__buf_2
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22374_ _12528_/A input46/X _22380_/S vssd1 vssd1 vccd1 vccd1 _22375_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15586__A _16770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21325_ _21609_/A _21595_/B vssd1 vssd1 vccd1 vccd1 _21325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15894__A1 _15890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21256_ _21683_/A _21299_/B _21260_/B vssd1 vssd1 vccd1 vccd1 _21256_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__22929__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20207_ _20463_/A _20463_/B _20207_/C vssd1 vssd1 vccd1 vccd1 _20210_/B sky130_fd_sc_hd__nand3_4
XFILLER_131_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21187_ _21187_/A vssd1 vssd1 vccd1 vccd1 _21187_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14449__A2 _16879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20138_ _20132_/X _20142_/B _20137_/X vssd1 vssd1 vccd1 vccd1 _20155_/A sky130_fd_sc_hd__a21o_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13121__A2 _21750_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20069_ _20069_/A _22828_/Q vssd1 vssd1 vccd1 vccd1 _20835_/A sky130_fd_sc_hd__and2_1
XFILLER_86_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12960_ _12960_/A _12960_/B vssd1 vssd1 vccd1 vccd1 _12963_/D sky130_fd_sc_hd__nand2_1
XFILLER_180_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_674 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _11911_/A vssd1 vssd1 vccd1 vccd1 _11912_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18060__A2 _17839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_538 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12891_/A vssd1 vssd1 vccd1 vccd1 _20182_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15471__D _15901_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_655 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _15061_/A _14512_/A _14512_/B _14629_/X vssd1 vssd1 vccd1 vccd1 _14635_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11842_/A _11842_/B _11842_/C vssd1 vssd1 vccd1 vccd1 _12247_/B sky130_fd_sc_hd__nand3_2
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _15182_/A _14561_/B _14561_/C _14561_/D vssd1 vssd1 vccd1 vccd1 _14561_/Y
+ sky130_fd_sc_hd__nor4_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11770_/X _11771_/X _18679_/C _11605_/A vssd1 vssd1 vccd1 vccd1 _11949_/D
+ sky130_fd_sc_hd__a31oi_4
XFILLER_14_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18137__A _19197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16300_/A vssd1 vssd1 vccd1 vccd1 _17443_/A sky130_fd_sc_hd__clkbuf_4
X_13512_ _13552_/A _13512_/B vssd1 vssd1 vccd1 vccd1 _13614_/C sky130_fd_sc_hd__nor2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _17280_/A vssd1 vssd1 vccd1 vccd1 _18659_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__14909__B1 _15082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14492_ _14500_/A _14611_/A _14490_/Y _14491_/X vssd1 vssd1 vccd1 vccd1 _14492_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ _12772_/A _12774_/A _16225_/X _16227_/X _17144_/C vssd1 vssd1 vccd1 vccd1
+ _16231_/X sky130_fd_sc_hd__o221a_2
XANTENNA__14385__A1 _18258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13443_ _13443_/A _13475_/A vssd1 vssd1 vccd1 vccd1 _13468_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14385__B2 _14863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16880__A _17039_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16162_ _16154_/X _16157_/X _16161_/Y vssd1 vssd1 vccd1 vccd1 _16162_/X sky130_fd_sc_hd__o21ba_1
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12935__A2 _20593_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13374_ _13426_/A vssd1 vssd1 vccd1 vccd1 _13579_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_943 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15113_ _15114_/A _15154_/A _15186_/A _15154_/B vssd1 vssd1 vccd1 vccd1 _15113_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14137__A1 _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12325_ _12368_/D _12324_/X _12320_/A vssd1 vssd1 vccd1 vccd1 _12577_/A sky130_fd_sc_hd__a21o_2
XFILLER_181_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16093_ _16093_/A _16093_/B _16134_/B vssd1 vssd1 vccd1 vccd1 _16093_/X sky130_fd_sc_hd__and3_1
XFILLER_177_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12913__A _12913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21670__A3 _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15885__A1 _15812_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19921_ _19921_/A _19921_/B vssd1 vssd1 vccd1 vccd1 _19921_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18303__C _18303_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15044_ _15044_/A _15044_/B vssd1 vssd1 vccd1 vccd1 _15045_/A sky130_fd_sc_hd__and2_1
X_12256_ _12256_/A vssd1 vssd1 vccd1 vccd1 _12258_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19852_ _19852_/A _19909_/C vssd1 vssd1 vccd1 vccd1 _19852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12726__A2_N _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12187_ _12183_/Y _12184_/Y _12185_/Y _12186_/Y vssd1 vssd1 vccd1 vccd1 _12188_/C
+ sky130_fd_sc_hd__o22ai_2
XFILLER_110_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18803_ _19202_/D _19353_/B _19353_/C vssd1 vssd1 vccd1 vccd1 _18804_/B sky130_fd_sc_hd__and3_1
XFILLER_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19783_ _19781_/B _19783_/B _19848_/B vssd1 vssd1 vccd1 vccd1 _19784_/C sky130_fd_sc_hd__nand3b_1
XFILLER_110_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16995_ _16709_/Y _16998_/A _16994_/Y vssd1 vssd1 vccd1 vccd1 _16997_/A sky130_fd_sc_hd__o21ai_1
XFILLER_95_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18734_ _18527_/Y _18557_/A _18729_/A vssd1 vssd1 vccd1 vccd1 _18736_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15946_ _15883_/A _15875_/A _15874_/B vssd1 vssd1 vccd1 vccd1 _15946_/X sky130_fd_sc_hd__a21o_1
XFILLER_77_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22383__A1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18665_ _18665_/A vssd1 vssd1 vccd1 vccd1 _19507_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15877_ _15759_/Y _15873_/X _15875_/Y _15876_/X vssd1 vssd1 vccd1 vccd1 _15877_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17616_ _17616_/A _17616_/B _17616_/C vssd1 vssd1 vccd1 vccd1 _17616_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__16601__A3 _16602_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21680__B _21680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14828_ _14764_/Y _14828_/B _14828_/C vssd1 vssd1 vccd1 vccd1 _14828_/Y sky130_fd_sc_hd__nand3b_1
X_18596_ _18970_/A _18596_/B vssd1 vssd1 vccd1 vccd1 _18606_/A sky130_fd_sc_hd__nand2_1
XFILLER_184_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17547_ _17531_/D _17678_/A _17546_/X vssd1 vssd1 vccd1 vccd1 _17663_/A sky130_fd_sc_hd__a21oi_1
X_14759_ _14661_/C _14549_/B _14758_/Y _14662_/Y vssd1 vssd1 vccd1 vccd1 _14759_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_177_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17478_ _17466_/B _17467_/X _17318_/A _17318_/B vssd1 vssd1 vccd1 vccd1 _17479_/D
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17562__A1 _17442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17562__B2 _16746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19217_ _19059_/Y _19215_/X _19216_/Y vssd1 vssd1 vccd1 vccd1 _19218_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__14376__A1 _22702_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11711__B _22960_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16429_ _16429_/A vssd1 vssd1 vccd1 vccd1 _16444_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18185__A_N _18278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19148_ _19148_/A _19148_/B _19148_/C vssd1 vssd1 vccd1 vccd1 _19148_/X sky130_fd_sc_hd__and3_1
XFILLER_192_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11430__C _11430_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17314__B2 _17007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18511__B1 _15774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19854__A3 _19793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19079_ _19079_/A vssd1 vssd1 vccd1 vccd1 _19254_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21110_ _21086_/C _21086_/B _21086_/D _21086_/A _21109_/X vssd1 vssd1 vccd1 vccd1
+ _21112_/A sky130_fd_sc_hd__a32oi_4
XFILLER_160_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22090_ _22090_/A _22090_/B vssd1 vssd1 vccd1 vccd1 _22145_/C sky130_fd_sc_hd__nand2_1
XFILLER_160_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21041_ _21041_/A _21041_/B vssd1 vssd1 vccd1 vccd1 _22920_/D sky130_fd_sc_hd__xor2_1
XFILLER_119_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18510__A _18510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17093__A3 _17460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22374__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21943_ _22041_/A vssd1 vssd1 vccd1 vccd1 _22037_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21874_ _21874_/A _22058_/A _21874_/C vssd1 vssd1 vccd1 vccd1 _21875_/C sky130_fd_sc_hd__and3_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20825_ _20759_/A _20759_/B _20890_/A vssd1 vssd1 vccd1 vccd1 _20830_/C sky130_fd_sc_hd__a21boi_1
XFILLER_78_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20756_ _20547_/X _20445_/Y _20652_/Y _20660_/A _20755_/Y vssd1 vssd1 vccd1 vccd1
+ _20759_/A sky130_fd_sc_hd__a41oi_4
XANTENNA__14367__A1 _22796_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11621__B _12154_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14367__B2 _14366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16761__C1 _17251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20687_ _21009_/A _15935_/A _20671_/Y _20717_/A _20608_/Y vssd1 vssd1 vccd1 vccd1
+ _20713_/B sky130_fd_sc_hd__o311a_1
XFILLER_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22426_ _22426_/A vssd1 vssd1 vccd1 vccd1 _22435_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19845__A3 _20012_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13590__A2 _21489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22357_ _22356_/B _22356_/C _22356_/A vssd1 vssd1 vccd1 vccd1 _22358_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ _12110_/A _12110_/B _12110_/C vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__nand3_4
X_21308_ _21312_/C vssd1 vssd1 vccd1 vccd1 _21739_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ _22843_/Q vssd1 vssd1 vccd1 vccd1 _21315_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_123_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22288_ _22325_/A vssd1 vssd1 vccd1 vccd1 _22297_/A sky130_fd_sc_hd__inv_2
XFILLER_6_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12041_ _22660_/B vssd1 vssd1 vccd1 vccd1 _12043_/A sky130_fd_sc_hd__inv_2
XFILLER_105_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21239_ _21239_/A _21239_/B _21239_/C vssd1 vssd1 vccd1 vccd1 _21247_/C sky130_fd_sc_hd__nand3_2
XFILLER_85_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20612__A1 _20685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18281__A2 _11861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17084__A3 _17875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15800_ _15780_/Y _15975_/B _15778_/Y vssd1 vssd1 vccd1 vccd1 _15801_/C sky130_fd_sc_hd__o21ai_1
XFILLER_59_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16780_ _18445_/A _18797_/B _17246_/A vssd1 vssd1 vccd1 vccd1 _16941_/A sky130_fd_sc_hd__nand3_2
XANTENNA__15482__C _15482_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13992_ _13992_/A _13992_/B _13992_/C vssd1 vssd1 vccd1 vccd1 _14009_/B sky130_fd_sc_hd__nand3_2
XFILLER_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ _15731_/A _15731_/B vssd1 vssd1 vccd1 vccd1 _15733_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12943_ _12950_/B _12708_/A _12700_/Y vssd1 vssd1 vccd1 vccd1 _12943_/X sky130_fd_sc_hd__a21o_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16875__A _17313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20915__A2 _17880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _18450_/A _18450_/B vssd1 vssd1 vccd1 vccd1 _18458_/C sky130_fd_sc_hd__nand2_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _15662_/A _15662_/B _15662_/C vssd1 vssd1 vccd1 vccd1 _16213_/A sky130_fd_sc_hd__nand3_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12874_ _12777_/X _12781_/X _12868_/X _20169_/A vssd1 vssd1 vccd1 vccd1 _12874_/Y
+ sky130_fd_sc_hd__o211ai_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17401_ _17401_/A _17401_/B _17401_/C _17401_/D vssd1 vssd1 vccd1 vccd1 _17401_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _12083_/A vssd1 vssd1 vccd1 vccd1 _11837_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14613_ _14613_/A vssd1 vssd1 vccd1 vccd1 _14892_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_92_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15593_ _15566_/A _15571_/Y _15581_/X _15579_/X vssd1 vssd1 vccd1 vccd1 _16287_/B
+ sky130_fd_sc_hd__o2bb2ai_2
X_18381_ _18381_/A _18381_/B _18381_/C vssd1 vssd1 vccd1 vccd1 _18408_/C sky130_fd_sc_hd__nand3_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12605__A1 _15799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12605__B2 _20456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12908__A _15558_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _17177_/A _17177_/B _17177_/C _17200_/A vssd1 vssd1 vccd1 vccd1 _17332_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_144_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14544_/A _14544_/B _14544_/C vssd1 vssd1 vccd1 vccd1 _14547_/C sky130_fd_sc_hd__nand3_1
XANTENNA__20679__B2 _15919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11756_ _11756_/A vssd1 vssd1 vccd1 vccd1 _12165_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17263_ _17298_/B _17298_/C _17298_/A vssd1 vssd1 vccd1 vccd1 _17299_/A sky130_fd_sc_hd__a21o_1
X_14475_ _14475_/A _14475_/B vssd1 vssd1 vccd1 vccd1 _14693_/A sky130_fd_sc_hd__nand2_1
XFILLER_186_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11687_ _12083_/B _11687_/B vssd1 vssd1 vccd1 vccd1 _11687_/Y sky130_fd_sc_hd__nor2_1
X_19002_ _19002_/A _19002_/B vssd1 vssd1 vccd1 vccd1 _19002_/Y sky130_fd_sc_hd__nor2_1
X_16214_ _15666_/A _15668_/X _15673_/B vssd1 vssd1 vccd1 vccd1 _16214_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13426_ _13426_/A _21351_/C vssd1 vssd1 vccd1 vccd1 _13428_/A sky130_fd_sc_hd__nand2_1
X_17194_ _17196_/A _17196_/B _17200_/B _17200_/C vssd1 vssd1 vccd1 vccd1 _17197_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16145_ _16145_/A _16145_/B _16145_/C vssd1 vssd1 vccd1 vccd1 _16145_/Y sky130_fd_sc_hd__nand3_1
XFILLER_155_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15307__B1 _15557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ _21234_/A _13338_/B _13315_/X _13354_/B vssd1 vssd1 vccd1 vccd1 _13358_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_182_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12308_ _22703_/Q vssd1 vssd1 vccd1 vccd1 _12520_/B sky130_fd_sc_hd__buf_2
XANTENNA__14561__C _14561_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16076_ _16047_/A _16047_/B _16074_/Y _16075_/X vssd1 vssd1 vccd1 vccd1 _16076_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_142_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13288_ _13288_/A _13288_/B _13288_/C vssd1 vssd1 vccd1 vccd1 _13484_/B sky130_fd_sc_hd__nand3_2
X_19904_ _19846_/B _19850_/B _19901_/X _19902_/X vssd1 vssd1 vccd1 vccd1 _19939_/A
+ sky130_fd_sc_hd__a211oi_2
X_15027_ _15107_/C _15026_/C _15026_/B vssd1 vssd1 vccd1 vccd1 _15028_/B sky130_fd_sc_hd__a21oi_1
X_12239_ _12241_/C _12241_/A _12240_/A _12240_/B vssd1 vssd1 vccd1 vccd1 _18236_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_69_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_714 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16807__B1 _15690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19835_ _19817_/B _19817_/C _19817_/A vssd1 vssd1 vccd1 vccd1 _19835_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17591__D _19482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16488__C _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19766_ _19836_/C _19842_/A _18030_/A _18028_/A _19705_/B vssd1 vssd1 vccd1 vccd1
+ _19807_/A sky130_fd_sc_hd__a41oi_4
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16978_ _16978_/A _16978_/B _17158_/A _17158_/B vssd1 vssd1 vccd1 vccd1 _16980_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__15491__C1 _17234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18984__B _18984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput4 wb_adr_i[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
X_18717_ _18681_/A _18684_/A _18862_/B vssd1 vssd1 vccd1 vccd1 _18722_/A sky130_fd_sc_hd__a21bo_1
X_15929_ _15853_/B _15843_/Y _15945_/B _15945_/C vssd1 vssd1 vccd1 vccd1 _16043_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19697_ _19768_/B _19697_/B _19774_/D _19697_/D vssd1 vssd1 vccd1 vccd1 _19698_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_655 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19161__A _19161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18648_ _19011_/A _18648_/B _19016_/A _18648_/D vssd1 vssd1 vccd1 vccd1 _18659_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_188_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18579_ _18761_/A _18570_/A _18574_/X vssd1 vssd1 vccd1 vccd1 _18582_/A sky130_fd_sc_hd__a21o_1
XFILLER_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20610_ _20606_/Y _20608_/Y _20609_/X vssd1 vssd1 vccd1 vccd1 _20613_/B sky130_fd_sc_hd__a21o_1
X_21590_ _21739_/C vssd1 vssd1 vccd1 vccd1 _22041_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13222__B1_N _13475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14349__A1 _12107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14349__B2 _12378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20541_ _20653_/A _20538_/B _20540_/X _20536_/X vssd1 vssd1 vccd1 vccd1 _20658_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20472_ _20471_/Y _20456_/Y _20468_/X vssd1 vssd1 vccd1 vccd1 _20599_/A sky130_fd_sc_hd__a21oi_1
XFILLER_119_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22211_ _22211_/A _22211_/B vssd1 vssd1 vccd1 vccd1 _22939_/D sky130_fd_sc_hd__xnor2_1
XFILLER_69_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22142_ _22142_/A _22142_/B _22164_/A _22159_/B vssd1 vssd1 vccd1 vccd1 _22156_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_106_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12272__B _12519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19336__A _19336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22073_ _22073_/A _22073_/B _22068_/C vssd1 vssd1 vccd1 vccd1 _22073_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_161_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22595__A1 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21024_ _21050_/C vssd1 vssd1 vccd1 vccd1 _21086_/C sky130_fd_sc_hd__buf_2
XANTENNA__19460__A1 _14432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11319__D _16308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17006__D _17006_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21926_ _22678_/Q _21927_/B _21927_/C _21922_/Y _21925_/Y vssd1 vssd1 vccd1 vccd1
+ _21929_/A sky130_fd_sc_hd__o311a_1
XFILLER_71_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11618__A_N _22790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16041__A4 _15935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15785__B1 _16465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21857_ _21857_/A _21857_/B _21857_/C vssd1 vssd1 vccd1 vccd1 _21865_/A sky130_fd_sc_hd__nand3_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1019 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12728__A _20207_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _18115_/D _11980_/A _11980_/B _11616_/C vssd1 vssd1 vccd1 vccd1 _11611_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_187_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20808_ _20806_/Y _20804_/Y _20178_/A _15935_/X vssd1 vssd1 vccd1 vccd1 _20808_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12590_ _15559_/C _15559_/D _20461_/C vssd1 vssd1 vccd1 vccd1 _12592_/A sky130_fd_sc_hd__nand3_2
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21788_ _21790_/A _21790_/B _21786_/Y _21787_/Y vssd1 vssd1 vccd1 vccd1 _21847_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_196_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21322__A2 _21591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11541_ _11541_/A vssd1 vssd1 vccd1 vccd1 _11541_/X sky130_fd_sc_hd__buf_6
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20739_ _20631_/B _20631_/C _20631_/A _20735_/Y vssd1 vssd1 vccd1 vccd1 _20739_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_169_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20664__B _20827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14260_ _14131_/X _14181_/C _14181_/A _14259_/X _14201_/X vssd1 vssd1 vccd1 vccd1
+ _14261_/B sky130_fd_sc_hd__a32o_1
X_11472_ _11587_/A vssd1 vssd1 vccd1 vccd1 _18093_/B sky130_fd_sc_hd__buf_2
XFILLER_13_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18134__B _18483_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ _13504_/A vssd1 vssd1 vccd1 vccd1 _13350_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22409_ _22705_/Q input43/X _22413_/S vssd1 vssd1 vccd1 vccd1 _22410_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14191_ _14191_/A _14191_/B _14191_/C _14595_/B vssd1 vssd1 vccd1 vccd1 _14195_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11574__A1 _19619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13142_ _13110_/Y _13234_/C _13112_/C vssd1 vssd1 vccd1 vccd1 _13147_/A sky130_fd_sc_hd__a21o_1
XFILLER_3_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input63_A wb_dat_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15774__A _18328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17950_ _17950_/A _17950_/B vssd1 vssd1 vccd1 vccd1 _17957_/A sky130_fd_sc_hd__nor2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _13073_/A _13097_/A _13301_/A vssd1 vssd1 vccd1 vccd1 _21214_/A sky130_fd_sc_hd__nand3_2
XFILLER_105_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16901_ _16682_/Y _16685_/A _16675_/Y _16698_/Y vssd1 vssd1 vccd1 vccd1 _16901_/Y
+ sky130_fd_sc_hd__o211ai_2
X_12024_ _12024_/A _12024_/B vssd1 vssd1 vccd1 vccd1 _12025_/C sky130_fd_sc_hd__nand2_1
XANTENNA__15493__B _19197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17881_ _19585_/D _21019_/B _21019_/A vssd1 vssd1 vccd1 vccd1 _17882_/A sky130_fd_sc_hd__and3_1
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19620_ _17436_/A _20012_/B _20012_/C _19618_/A _19614_/A vssd1 vssd1 vccd1 vccd1
+ _19621_/C sky130_fd_sc_hd__a32o_1
X_16832_ _16845_/A _17189_/B _16830_/Y _16831_/X vssd1 vssd1 vccd1 vccd1 _16906_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15473__C1 _19016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19551_ _19545_/C _19545_/B _19545_/A vssd1 vssd1 vccd1 vccd1 _19551_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__19203__A1 _12064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16763_ _16494_/A _16760_/X _16766_/A vssd1 vssd1 vccd1 vccd1 _16773_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11629__A2 _11626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ _14112_/A _14963_/B _14110_/B _13975_/D vssd1 vssd1 vccd1 vccd1 _13975_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16017__A1 _16015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16017__B2 _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18502_ _22797_/Q vssd1 vssd1 vccd1 vccd1 _18678_/D sky130_fd_sc_hd__inv_2
XANTENNA__21010__A1 _12671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15714_ _15714_/A _15714_/B _16515_/A _16772_/A vssd1 vssd1 vccd1 vccd1 _15714_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_46_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21010__B2 _21082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19482_ _19482_/A _20012_/B _20012_/C vssd1 vssd1 vccd1 vccd1 _19630_/D sky130_fd_sc_hd__and3_1
XFILLER_20_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ _12926_/A _12926_/B _12926_/C vssd1 vssd1 vccd1 vccd1 _12933_/A sky130_fd_sc_hd__nand3_1
X_16694_ _22889_/Q _16424_/A _22890_/Q vssd1 vssd1 vccd1 vccd1 _16694_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18433_ _18432_/B _18432_/C _18432_/A vssd1 vssd1 vccd1 vccd1 _18434_/B sky130_fd_sc_hd__a21o_1
XFILLER_94_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15645_ _16332_/A vssd1 vssd1 vccd1 vccd1 _15645_/X sky130_fd_sc_hd__buf_4
XANTENNA__14579__B2 _14942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12857_ _12857_/A vssd1 vssd1 vccd1 vccd1 _12862_/B sky130_fd_sc_hd__clkbuf_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12638__A _16498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19506__A2 _12171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11542__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18364_ _18471_/C _18471_/B _18471_/A vssd1 vssd1 vccd1 vccd1 _18387_/A sky130_fd_sc_hd__nand3_2
X_11808_ _11630_/Y _11807_/Y _11647_/A vssd1 vssd1 vccd1 vccd1 _12035_/B sky130_fd_sc_hd__o21ai_2
X_15576_ _16912_/A vssd1 vssd1 vccd1 vccd1 _17672_/A sky130_fd_sc_hd__buf_4
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _16489_/A _12788_/B _12788_/C _20502_/C vssd1 vssd1 vccd1 vccd1 _12792_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22510__A1 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17523_/A _17520_/C vssd1 vssd1 vccd1 vccd1 _17318_/A sky130_fd_sc_hd__nand2_1
XFILLER_42_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11739_ _11625_/X _11626_/X _11737_/X _11738_/X _15458_/A vssd1 vssd1 vccd1 vccd1
+ _11739_/Y sky130_fd_sc_hd__o221ai_1
X_14527_ _13942_/Y _13911_/X _13903_/Y _13937_/C _13937_/D vssd1 vssd1 vccd1 vccd1
+ _14527_/Y sky130_fd_sc_hd__o2111ai_4
X_18295_ _18636_/A _17526_/X _18281_/Y _12216_/X _18289_/Y vssd1 vssd1 vccd1 vccd1
+ _18295_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__11801__A2 _11639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17246_ _17246_/A _17532_/C _17532_/D vssd1 vssd1 vccd1 vccd1 _17247_/A sky130_fd_sc_hd__nand3_1
X_14458_ _15205_/B vssd1 vssd1 vccd1 vccd1 _14987_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1048 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13409_ _13572_/B vssd1 vssd1 vccd1 vccd1 _13664_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_17177_ _17177_/A _17177_/B _17177_/C vssd1 vssd1 vccd1 vccd1 _17200_/B sky130_fd_sc_hd__nand3_2
XFILLER_116_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14389_ _22801_/Q _14381_/X _14382_/X _14331_/X _22705_/Q vssd1 vssd1 vccd1 vccd1
+ _14389_/X sky130_fd_sc_hd__a32o_1
XFILLER_183_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16128_ _16143_/A _16143_/B vssd1 vssd1 vccd1 vccd1 _16186_/B sky130_fd_sc_hd__nand2_1
XFILLER_182_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19690__A1 _12207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16059_ _16059_/A vssd1 vssd1 vccd1 vccd1 _16060_/A sky130_fd_sc_hd__buf_2
XFILLER_143_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19818_ _19823_/A _19818_/B vssd1 vssd1 vccd1 vccd1 _19880_/C sky130_fd_sc_hd__nand2_1
XFILLER_116_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19749_ _19761_/A _19761_/B _19761_/D _19760_/A _19760_/B vssd1 vssd1 vccd1 vccd1
+ _19749_/X sky130_fd_sc_hd__a32o_1
XANTENNA__13932__A _22873_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22760_ _22762_/CLK _22760_/D vssd1 vssd1 vccd1 vccd1 _22760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19322__C _19322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16559__A2 _15378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21711_ _21711_/A _21711_/B vssd1 vssd1 vccd1 vccd1 _22933_/D sky130_fd_sc_hd__xnor2_1
X_22691_ _22693_/CLK _22691_/D vssd1 vssd1 vccd1 vccd1 _22691_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13778__C1 _14503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21642_ _21654_/B _21641_/A _21654_/A vssd1 vssd1 vccd1 vccd1 _21642_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21573_ _21573_/A _21573_/B vssd1 vssd1 vccd1 vccd1 _22932_/D sky130_fd_sc_hd__xnor2_1
XFILLER_166_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20524_ _20513_/Y _20515_/X _20491_/Y _20501_/X vssd1 vssd1 vccd1 vccd1 _20526_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_192_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21299__C _21683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20455_ _20340_/Y _20343_/Y _20344_/Y _20347_/Y vssd1 vssd1 vccd1 vccd1 _20455_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20386_ _20397_/B _20386_/B vssd1 vssd1 vccd1 vccd1 _20388_/B sky130_fd_sc_hd__nand2_1
XFILLER_161_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15298__A2 _12774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22125_ _22128_/A _22219_/A _22128_/C vssd1 vssd1 vccd1 vccd1 _22125_/X sky130_fd_sc_hd__and3_1
XFILLER_134_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22056_ _21579_/A _21473_/Y _22055_/Y vssd1 vssd1 vccd1 vccd1 _22262_/A sky130_fd_sc_hd__a21oi_4
XFILLER_102_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21007_ _21067_/D _21007_/B _21007_/C vssd1 vssd1 vccd1 vccd1 _21037_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19984__A2 _20012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16798__A2 _15903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13811__A_N _13826_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13760_ _22754_/Q vssd1 vssd1 vccd1 vccd1 _13761_/B sky130_fd_sc_hd__clkbuf_4
X_22958_ _22964_/CLK _22958_/D vssd1 vssd1 vccd1 vccd1 _22958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21909_ _21909_/A _21909_/B vssd1 vssd1 vccd1 vccd1 _21909_/Y sky130_fd_sc_hd__nand2_1
X_12711_ _20478_/C vssd1 vssd1 vccd1 vccd1 _12711_/X sky130_fd_sc_hd__clkbuf_2
X_13691_ _13707_/B vssd1 vssd1 vccd1 vccd1 _13776_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_71_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22889_ _22952_/CLK _22889_/D vssd1 vssd1 vccd1 vccd1 _22889_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15430_ _15430_/A _15430_/B _15430_/C vssd1 vssd1 vccd1 vccd1 _15700_/C sky130_fd_sc_hd__nand3_2
X_12642_ _12745_/A _12745_/C vssd1 vssd1 vccd1 vccd1 _12643_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15361_ _20341_/A vssd1 vssd1 vccd1 vccd1 _20101_/A sky130_fd_sc_hd__buf_2
X_12573_ _22821_/Q vssd1 vssd1 vccd1 vccd1 _20101_/C sky130_fd_sc_hd__buf_4
XFILLER_178_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16368__A1_N _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17100_ _17310_/A _17341_/C _17098_/Y _17099_/X vssd1 vssd1 vccd1 vccd1 _17338_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_11_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11524_ _11430_/B _18116_/A _18482_/B _18482_/A _12003_/B vssd1 vssd1 vccd1 vccd1
+ _11581_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14312_ _14410_/A vssd1 vssd1 vccd1 vccd1 _14351_/A sky130_fd_sc_hd__clkbuf_2
X_18080_ _18080_/A vssd1 vssd1 vccd1 vccd1 _18080_/Y sky130_fd_sc_hd__inv_2
X_15292_ _22885_/Q _15292_/B vssd1 vssd1 vccd1 vccd1 _22873_/D sky130_fd_sc_hd__xnor2_1
XFILLER_141_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17031_ _17036_/A _17036_/B _17031_/C vssd1 vssd1 vccd1 vccd1 _17033_/B sky130_fd_sc_hd__nand3_1
X_14243_ _14243_/A _14243_/B vssd1 vssd1 vccd1 vccd1 _14246_/B sky130_fd_sc_hd__nor2_1
XANTENNA__17984__A _19419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11455_ _18203_/A vssd1 vssd1 vccd1 vccd1 _11818_/A sky130_fd_sc_hd__buf_2
XFILLER_125_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20267__C1 _20234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14174_ _14165_/X _14166_/Y _14169_/X _14090_/Y _14170_/X vssd1 vssd1 vccd1 vccd1
+ _14175_/C sky130_fd_sc_hd__o221ai_1
XANTENNA__19672__A1 _19293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11386_ _11386_/A vssd1 vssd1 vccd1 vccd1 _11503_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_194_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15289__A2 _15271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13125_ _13125_/A vssd1 vssd1 vccd1 vccd1 _21220_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18982_ _17083_/A _18889_/X _18890_/X _19772_/B _17313_/D vssd1 vssd1 vccd1 vccd1
+ _18982_/X sky130_fd_sc_hd__o311a_2
XFILLER_113_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12921__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17933_ _19941_/A _17883_/B _21044_/B _17928_/X _17932_/Y vssd1 vssd1 vccd1 vccd1
+ _17935_/C sky130_fd_sc_hd__o311a_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _22725_/Q vssd1 vssd1 vccd1 vccd1 _13112_/C sky130_fd_sc_hd__clkinv_2
XFILLER_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13736__B _13736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ _11972_/Y _11976_/Y _11986_/X _12006_/Y vssd1 vssd1 vccd1 vccd1 _12007_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_87_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17864_ _17849_/Y _17854_/X _17863_/X vssd1 vssd1 vccd1 vccd1 _17864_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__18632__C1 _18953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater129 _22871_/Q vssd1 vssd1 vccd1 vccd1 _22859_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__16789__A2 _16179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_bq_clk_i clkbuf_3_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_19603_ _18131_/B _19769_/B _18131_/C _19602_/B _19602_/A vssd1 vssd1 vccd1 vccd1
+ _19603_/X sky130_fd_sc_hd__a32o_1
XFILLER_93_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16815_ _19461_/A _15960_/A _17131_/B _18839_/B vssd1 vssd1 vccd1 vccd1 _16815_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_94_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17795_ _17795_/A _17795_/B _17795_/C vssd1 vssd1 vccd1 vccd1 _17797_/A sky130_fd_sc_hd__and3_1
X_19534_ _19538_/A _19538_/B _19538_/C vssd1 vssd1 vccd1 vccd1 _19536_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13752__A _14808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16746_ _17091_/A vssd1 vssd1 vccd1 vccd1 _16746_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13958_ _14506_/C vssd1 vssd1 vccd1 vccd1 _14911_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19465_ _19465_/A _19614_/B _19614_/C vssd1 vssd1 vccd1 vccd1 _19465_/Y sky130_fd_sc_hd__nand3_1
X_12909_ _20207_/C vssd1 vssd1 vccd1 vccd1 _20481_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16677_ _22892_/Q vssd1 vssd1 vccd1 vccd1 _16685_/A sky130_fd_sc_hd__clkinv_4
XFILLER_61_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13889_ _13881_/Y _13883_/Y _13884_/X vssd1 vssd1 vccd1 vccd1 _13889_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_62_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18416_ _18416_/A vssd1 vssd1 vccd1 vccd1 _18417_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ _20471_/B vssd1 vssd1 vccd1 vccd1 _16563_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_195_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19396_ _19396_/A _19396_/B _19396_/C vssd1 vssd1 vccd1 vccd1 _19396_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__14421__B1 _14413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18347_ _18137_/Y _18139_/X _18141_/Y _18150_/B vssd1 vssd1 vccd1 vccd1 _18351_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_15559_ _16257_/A _15559_/B _15559_/C _15559_/D vssd1 vssd1 vccd1 vccd1 _15559_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_187_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19360__B1 _19176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_672 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18278_ _18278_/A _18278_/B vssd1 vssd1 vccd1 vccd1 _18279_/B sky130_fd_sc_hd__nand2_1
XFILLER_174_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17229_ _17229_/A _17603_/C vssd1 vssd1 vccd1 vccd1 _17229_/Y sky130_fd_sc_hd__nor2_1
Xinput40 wb_dat_i[14] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_2
Xinput51 wb_dat_i[24] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 wb_dat_i[5] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput73 x[2] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
X_20240_ _20240_/A _20240_/B _20240_/C vssd1 vssd1 vccd1 vccd1 _20266_/A sky130_fd_sc_hd__nand3_2
XFILLER_157_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17674__B1 _19793_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20171_ _12781_/B _12886_/X _20165_/Y _20181_/B vssd1 vssd1 vccd1 vccd1 _20174_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19317__C _19461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22962__CLK _22964_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16229__A1 _14429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19614__A _19614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17977__A1 _21050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17441__A3 _17110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18875__D _18875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13662__A _13662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22812_ _22812_/CLK _22812_/D vssd1 vssd1 vccd1 vccd1 _22812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19052__C _19346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17729__A1 _17806_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22743_ _22743_/CLK _22743_/D vssd1 vssd1 vccd1 vccd1 _22743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16401__A1 _16397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15204__A2 _15205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22674_ _22943_/CLK _22674_/D vssd1 vssd1 vccd1 vccd1 _22674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21625_ _21449_/A _21449_/B _21460_/C vssd1 vssd1 vccd1 vccd1 _21654_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__20926__C _20936_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18154__A1 _12157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21556_ _21556_/A vssd1 vssd1 vccd1 vccd1 _21556_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21103__B _22942_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20507_ _20511_/A _20511_/B _20504_/X _20506_/Y vssd1 vssd1 vccd1 vccd1 _20519_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15101__B _15101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21487_ _21185_/X _21187_/X _22229_/A vssd1 vssd1 vccd1 vccd1 _21872_/A sky130_fd_sc_hd__o21a_1
XFILLER_5_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12726__B1 _12721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22860__D _22872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20438_ _20439_/A _20439_/B _22932_/Q vssd1 vssd1 vccd1 vccd1 _20563_/A sky130_fd_sc_hd__a21o_1
XANTENNA__19654__A1 _19652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20369_ _20250_/C _20611_/A _20511_/A _20370_/D vssd1 vssd1 vccd1 vccd1 _20371_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_171_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18131__C _18131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22108_ _22221_/A _22221_/B _22108_/C vssd1 vssd1 vccd1 vccd1 _22108_/Y sky130_fd_sc_hd__nand3_2
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15691__A2 _15808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22039_ _21853_/X _21958_/X _22037_/Y _22038_/X vssd1 vssd1 vccd1 vccd1 _22039_/Y
+ sky130_fd_sc_hd__o211ai_2
X_14930_ _14930_/A _14930_/B vssd1 vssd1 vccd1 vccd1 _14961_/A sky130_fd_sc_hd__and2_1
XFILLER_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input26_A wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ _14861_/A _14868_/B _14861_/C vssd1 vssd1 vccd1 vccd1 _14932_/A sky130_fd_sc_hd__nand3_2
XFILLER_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16600_ _16354_/A _16310_/Y _16354_/C vssd1 vssd1 vccd1 vccd1 _16600_/X sky130_fd_sc_hd__o21a_1
XANTENNA__16586__C _17313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13812_ _22767_/Q vssd1 vssd1 vccd1 vccd1 _13826_/B sky130_fd_sc_hd__buf_2
XFILLER_91_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17580_ _17580_/A vssd1 vssd1 vccd1 vccd1 _17580_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14792_ _14792_/A _14792_/B vssd1 vssd1 vccd1 vccd1 _14935_/A sky130_fd_sc_hd__nand2_2
X_16531_ _16283_/A _16283_/B _16288_/C _16530_/X vssd1 vssd1 vccd1 vccd1 _16531_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13743_ _22767_/Q vssd1 vssd1 vccd1 vccd1 _13773_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19250_ _19192_/Y _19238_/Y _19248_/Y _19249_/Y vssd1 vssd1 vccd1 vccd1 _19250_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_31_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16462_ _16257_/Y _16816_/A _16452_/X _15694_/A _20608_/A vssd1 vssd1 vccd1 vccd1
+ _16463_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_177_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ _13674_/A _13674_/B _13674_/C vssd1 vssd1 vccd1 vccd1 _13674_/Y sky130_fd_sc_hd__nand3_1
XFILLER_73_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18201_ _18199_/Y _18200_/Y _17632_/A _12050_/B _18195_/Y vssd1 vssd1 vccd1 vccd1
+ _18571_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_31_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15413_ _20092_/A vssd1 vssd1 vccd1 vccd1 _20675_/A sky130_fd_sc_hd__buf_2
X_19181_ _19190_/A _19190_/B _19182_/C vssd1 vssd1 vccd1 vccd1 _19240_/C sky130_fd_sc_hd__a21o_1
X_12625_ _16486_/C vssd1 vssd1 vccd1 vccd1 _15586_/C sky130_fd_sc_hd__buf_2
X_16393_ _16393_/A _16393_/B _16393_/C vssd1 vssd1 vccd1 vccd1 _16429_/A sky130_fd_sc_hd__nand3_1
XFILLER_106_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22835__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__A _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18132_ _18125_/X _18130_/Y _18131_/X vssd1 vssd1 vccd1 vccd1 _18132_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14834__C _14834_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15344_ _15344_/A vssd1 vssd1 vccd1 vccd1 _15344_/X sky130_fd_sc_hd__clkbuf_2
X_12556_ _12669_/A vssd1 vssd1 vccd1 vccd1 _16486_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_156_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11507_ _11502_/X _11503_/X _11504_/X _11505_/X _11779_/B vssd1 vssd1 vccd1 vccd1
+ _11507_/X sky130_fd_sc_hd__o221a_2
XANTENNA__13509__A2 _22106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18063_ _18063_/A _18063_/B vssd1 vssd1 vccd1 vccd1 _18063_/X sky130_fd_sc_hd__xor2_1
XFILLER_157_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15275_ _22879_/Q _15275_/B vssd1 vssd1 vccd1 vccd1 _22867_/D sky130_fd_sc_hd__xnor2_1
X_12487_ _16515_/A _12487_/B _12487_/C _20486_/C vssd1 vssd1 vccd1 vccd1 _12487_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_172_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12717__B1 _22821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17014_ _16990_/Y _16991_/Y _17006_/Y _17008_/Y vssd1 vssd1 vccd1 vccd1 _17025_/A
+ sky130_fd_sc_hd__o211ai_2
X_11438_ _11448_/A _11438_/B vssd1 vssd1 vccd1 vccd1 _11438_/Y sky130_fd_sc_hd__nand2_1
X_14226_ _14226_/A _15114_/D _14273_/A vssd1 vssd1 vccd1 vccd1 _14243_/A sky130_fd_sc_hd__and3_1
XANTENNA__18448__A2 _17380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13747__A _22865_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ _14157_/A vssd1 vssd1 vccd1 vccd1 _14272_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_153_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11369_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11796_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16123__A _19012_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15665__C _15665_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _22721_/Q _22720_/Q vssd1 vssd1 vccd1 vccd1 _13143_/B sky130_fd_sc_hd__nor2_2
XANTENNA__21964__A _21964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18965_ _18965_/A _18965_/B vssd1 vssd1 vccd1 vccd1 _18967_/B sky130_fd_sc_hd__nand2_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _14147_/B _14147_/C _14147_/D _14087_/Y vssd1 vssd1 vccd1 vccd1 _14167_/C
+ sky130_fd_sc_hd__a31oi_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17916_ _22903_/Q _17970_/B vssd1 vssd1 vccd1 vccd1 _18007_/C sky130_fd_sc_hd__xor2_1
XANTENNA__15962__A _17039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14485__A3 _14684_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13039_ _13039_/A _13039_/B vssd1 vssd1 vccd1 vccd1 _13040_/C sky130_fd_sc_hd__nor2_1
XFILLER_21_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18896_ _19329_/D _19329_/C _18896_/C _19587_/D vssd1 vssd1 vccd1 vccd1 _19022_/C
+ sky130_fd_sc_hd__and4_2
XANTENNA__12496__A2 _12493_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21755__A2 _14380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17847_ _17787_/B _17787_/A _17857_/B vssd1 vssd1 vccd1 vccd1 _17847_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18620__A2 _17526_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17778_ _17778_/A _17778_/B vssd1 vssd1 vccd1 vccd1 _17778_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14297__B input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19517_ _19517_/A vssd1 vssd1 vccd1 vccd1 _19981_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11456__B1 _15435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16729_ _20584_/A vssd1 vssd1 vccd1 vccd1 _20792_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12799__A3 _16498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19448_ _19301_/Y _19750_/A _19681_/B vssd1 vssd1 vccd1 vccd1 _19449_/B sky130_fd_sc_hd__a21o_1
XFILLER_34_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17592__C1 _17591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17401__B _17401_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19379_ _19379_/A _19379_/B vssd1 vssd1 vccd1 vccd1 _19379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18136__A1 _15887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11759__A1 _11703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21410_ _21410_/A _21410_/B _21410_/C vssd1 vssd1 vccd1 vccd1 _21411_/A sky130_fd_sc_hd__nand3_1
X_22390_ _22390_/A vssd1 vssd1 vccd1 vccd1 _22696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1096 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21341_ _21341_/A vssd1 vssd1 vccd1 vccd1 _21341_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20762__B _20827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21272_ _21264_/Y _21267_/X _21281_/C vssd1 vssd1 vccd1 vccd1 _21278_/A sky130_fd_sc_hd__o21ai_1
XFILLER_144_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13381__B1 _21638_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20223_ _12450_/X _15366_/A _20221_/Y _20457_/B vssd1 vssd1 vccd1 vccd1 _20224_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__20246__A2 _12735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17129__A _17234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11392__C1 _18984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15658__C1 _16361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21874__A _21874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20154_ _20154_/A _20154_/B _20197_/A _20197_/B vssd1 vssd1 vccd1 vccd1 _20158_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13133__B1 _21580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20085_ _12702_/A _20359_/C _20359_/A _20083_/X vssd1 vssd1 vccd1 vccd1 _20085_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18611__A2 _12171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14488__A _14684_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_804 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11905__A _11905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19021__C1 _17672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20987_ _20987_/A _20987_/B vssd1 vssd1 vccd1 vccd1 _21008_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__20706__B1 _20210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11998__A1 _16241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22858__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22726_ _22728_/CLK _22726_/D vssd1 vssd1 vccd1 vccd1 _22726_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__22855__D _22867_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_583 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_22 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_959 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18407__B _18407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17311__B _17311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22657_ _22657_/A vssd1 vssd1 vccd1 vccd1 _22815_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _15631_/A _15631_/B _15325_/A vssd1 vssd1 vccd1 vccd1 _16465_/A sky130_fd_sc_hd__a21oi_4
X_21608_ _21185_/X _21187_/X _21494_/B _21609_/A vssd1 vssd1 vccd1 vccd1 _21613_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ _21249_/B _13390_/B vssd1 vssd1 vccd1 vccd1 _13391_/B sky130_fd_sc_hd__xnor2_1
XFILLER_166_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22588_ _22656_/S vssd1 vssd1 vccd1 vccd1 _22597_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_139_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12341_ _12341_/A _12520_/B vssd1 vssd1 vccd1 vccd1 _12378_/A sky130_fd_sc_hd__nand2_2
XFILLER_127_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21539_ _21539_/A _21539_/B vssd1 vssd1 vccd1 vccd1 _21539_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15060_ _14818_/A _15006_/Y _15185_/B _15058_/X _15059_/Y vssd1 vssd1 vccd1 vccd1
+ _15060_/X sky130_fd_sc_hd__o311a_1
XFILLER_153_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ _12396_/C _12519_/B vssd1 vssd1 vccd1 vccd1 _12300_/B sky130_fd_sc_hd__nand2_1
XFILLER_181_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14011_ _14034_/A _14034_/B _14035_/A _14523_/A vssd1 vssd1 vccd1 vccd1 _14031_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17638__B1 _17440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13372__B1 _13202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20237__A2 _20579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17039__A _17039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13911__A2 _13814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17102__A2 _17338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12580__D1 _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17981__B _18023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16878__A _20936_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18750_ _18645_/Y _18646_/X _18748_/A vssd1 vssd1 vccd1 vccd1 _18753_/A sky130_fd_sc_hd__o21ai_1
XFILLER_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15962_ _17039_/A _20806_/C _17643_/A _17039_/D vssd1 vssd1 vccd1 vccd1 _15962_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_95_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17701_ _17701_/A _17701_/B _17701_/C vssd1 vssd1 vccd1 vccd1 _17702_/B sky130_fd_sc_hd__nand3_1
X_14913_ _14972_/A _14914_/C _14972_/B vssd1 vssd1 vccd1 vccd1 _14916_/C sky130_fd_sc_hd__o21ai_1
X_18681_ _18681_/A vssd1 vssd1 vccd1 vccd1 _18869_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15893_ _15893_/A _15901_/B _15893_/C vssd1 vssd1 vccd1 vccd1 _15900_/A sky130_fd_sc_hd__nand3_4
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15416__A2 _15919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16074__C1 _15918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17632_ _17632_/A vssd1 vssd1 vccd1 vccd1 _19774_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_84_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14844_ _14929_/A _14929_/B vssd1 vssd1 vccd1 vccd1 _14845_/C sky130_fd_sc_hd__nor2_1
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17563_ _17564_/A _17564_/B _17562_/Y _17006_/A _16124_/X vssd1 vssd1 vccd1 vccd1
+ _17574_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14775_ _14775_/A _14863_/A _14775_/C _14775_/D vssd1 vssd1 vccd1 vccd1 _14869_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_1_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ _15482_/A vssd1 vssd1 vccd1 vccd1 _16241_/A sky130_fd_sc_hd__buf_4
XFILLER_95_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19302_ _19299_/A _19299_/B _19299_/C vssd1 vssd1 vccd1 vccd1 _19302_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ _16472_/Y _16474_/Y _16513_/X vssd1 vssd1 vccd1 vccd1 _16517_/A sky130_fd_sc_hd__o21ai_1
XFILLER_56_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17502__A _17502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13726_ _13810_/A _13810_/B _13725_/Y vssd1 vssd1 vccd1 vccd1 _13727_/A sky130_fd_sc_hd__a21o_1
X_17494_ _17494_/A _17514_/A _17600_/A vssd1 vssd1 vccd1 vccd1 _17497_/B sky130_fd_sc_hd__nand3_1
XFILLER_182_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14845__B _14845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19233_ _19246_/B vssd1 vssd1 vccd1 vccd1 _19400_/B sky130_fd_sc_hd__inv_2
XFILLER_143_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16445_ _16397_/X _15630_/X _16652_/A vssd1 vssd1 vccd1 vccd1 _16445_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13657_ _13657_/A _13657_/B _13657_/C vssd1 vssd1 vccd1 vccd1 _13658_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19315__B1 _11511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14564__C _14564_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19164_ _19162_/Y _19163_/X _19185_/A _19155_/Y _19185_/C vssd1 vssd1 vccd1 vccd1
+ _19343_/A sky130_fd_sc_hd__o2111ai_4
XANTENNA__21959__A _22108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ _12606_/X _12607_/X _12450_/X vssd1 vssd1 vccd1 vccd1 _12608_/X sky130_fd_sc_hd__a21o_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _16286_/Y _16287_/Y _16288_/Y _16291_/Y vssd1 vssd1 vccd1 vccd1 _16704_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18669__A2 _18371_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13588_ _13461_/B _13521_/Y _13517_/X _13528_/X vssd1 vssd1 vccd1 vccd1 _13588_/X
+ sky130_fd_sc_hd__o211a_1
X_18115_ _18115_/A _22789_/Q _18115_/C _18115_/D vssd1 vssd1 vccd1 vccd1 _18116_/B
+ sky130_fd_sc_hd__nor4_1
XANTENNA__17877__B1 _17922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15327_ _15325_/X _15326_/X _15776_/B _15776_/A _16257_/C vssd1 vssd1 vccd1 vccd1
+ _15327_/Y sky130_fd_sc_hd__o2111ai_4
XANTENNA__20476__A2 _20579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19095_ _19095_/A _19095_/B _19095_/C vssd1 vssd1 vccd1 vccd1 _19106_/B sky130_fd_sc_hd__nand3_2
X_12539_ _12547_/A _12548_/A vssd1 vssd1 vccd1 vccd1 _20611_/B sky130_fd_sc_hd__nor2_4
XFILLER_144_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20582__B _20792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18046_ _18082_/C _18048_/A _18048_/B _18045_/Y vssd1 vssd1 vccd1 vccd1 _18046_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15258_ _15259_/A _15259_/C _15259_/B vssd1 vssd1 vccd1 vccd1 _15260_/A sky130_fd_sc_hd__o21a_1
XFILLER_144_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22622__A0 _18258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14209_ _14510_/A vssd1 vssd1 vccd1 vccd1 _14917_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15189_ _15189_/A vssd1 vssd1 vccd1 vccd1 _15238_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11913__A1 _11566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20779__A3 _17444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16301__B1 _15797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19997_ _19998_/B _19998_/A vssd1 vssd1 vccd1 vccd1 _20024_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18948_ _18778_/B _19983_/A _18626_/Y _18629_/Y _18625_/X vssd1 vssd1 vccd1 vccd1
+ _18952_/C sky130_fd_sc_hd__o32a_2
XFILLER_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18879_ _15904_/X _15905_/X _18857_/A _18858_/A vssd1 vssd1 vccd1 vccd1 _18880_/B
+ sky130_fd_sc_hd__o211a_2
X_20910_ _20514_/X _16746_/X _20854_/Y vssd1 vssd1 vccd1 vccd1 _20910_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_95_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21890_ _21896_/A vssd1 vssd1 vccd1 vccd1 _21996_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11444__B _18288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20841_ _20828_/A _20994_/B _20907_/A vssd1 vssd1 vccd1 vccd1 _20897_/A sky130_fd_sc_hd__o21ai_1
XFILLER_70_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_667 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20772_ _20772_/A _20772_/B _20772_/C _20772_/D vssd1 vssd1 vccd1 vccd1 _20773_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22511_ _22511_/A vssd1 vssd1 vccd1 vccd1 _22750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17131__B _17131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12556__A _12669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19306__B1 _19983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22442_ _22514_/A _22442_/B _22586_/C vssd1 vssd1 vccd1 vccd1 _22499_/A sky130_fd_sc_hd__and3_1
XFILLER_195_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15591__A1 _15498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18514__D1 _18876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15867__A _20678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22373_ _22373_/A vssd1 vssd1 vccd1 vccd1 _22688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21324_ _13295_/X _21329_/B _21336_/B _21336_/C _14359_/X vssd1 vssd1 vccd1 vccd1
+ _21324_/X sky130_fd_sc_hd__o311a_1
XFILLER_191_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15586__B _16771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15894__A2 _16098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22613__A0 _18128_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21255_ _21990_/B vssd1 vssd1 vccd1 vccd1 _21683_/A sky130_fd_sc_hd__buf_2
XFILLER_144_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20206_ _20463_/A _20463_/B _20357_/B _20086_/A _20101_/C vssd1 vssd1 vccd1 vccd1
+ _20206_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_81_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18293__B1 _18636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21186_ _21188_/A _21188_/B _13302_/A _14359_/X vssd1 vssd1 vccd1 vccd1 _21187_/A
+ sky130_fd_sc_hd__o31ai_2
XFILLER_131_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20137_ _12838_/B _20126_/Y _20142_/A vssd1 vssd1 vccd1 vccd1 _20137_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11338__C _15539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20068_ _20069_/A _22828_/Q vssd1 vssd1 vccd1 vccd1 _20834_/A sky130_fd_sc_hd__nor2_2
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _11868_/Y _11871_/X _11869_/X vssd1 vssd1 vccd1 vccd1 _11914_/A sky130_fd_sc_hd__a21oi_1
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22680__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18060__A3 _17839_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17025__C _17025_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _13043_/B vssd1 vssd1 vccd1 vccd1 _20183_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11841_ _11576_/B _11902_/C _11902_/B vssd1 vssd1 vccd1 vccd1 _11842_/A sky130_fd_sc_hd__a21boi_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_678 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _14560_/A vssd1 vssd1 vccd1 vccd1 _15182_/A sky130_fd_sc_hd__buf_2
X_11772_ _11772_/A vssd1 vssd1 vccd1 vccd1 _18679_/C sky130_fd_sc_hd__buf_2
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14665__B _14843_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13546_/A _13509_/X _13526_/A _13506_/C vssd1 vssd1 vccd1 vccd1 _13512_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__14909__A1 _13833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22709_ _22742_/CLK _22709_/D vssd1 vssd1 vccd1 vccd1 _22709_/Q sky130_fd_sc_hd__dfxtp_1
X_14491_ _14626_/A _14494_/B _14491_/C _14494_/D vssd1 vssd1 vccd1 vccd1 _14491_/X
+ sky130_fd_sc_hd__and4_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _17251_/A vssd1 vssd1 vccd1 vccd1 _17144_/C sky130_fd_sc_hd__buf_2
X_13442_ _13475_/C _13475_/B vssd1 vssd1 vccd1 vccd1 _13443_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16880__B _21050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13593__B1 _13126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16161_ _16154_/X _16157_/X _16159_/X _16174_/B vssd1 vssd1 vccd1 vccd1 _16161_/Y
+ sky130_fd_sc_hd__a22oi_1
X_13373_ _13373_/A _13373_/B vssd1 vssd1 vccd1 vccd1 _13426_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21498__B _21498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15112_ _15112_/A _15112_/B vssd1 vssd1 vccd1 vccd1 _15145_/A sky130_fd_sc_hd__xnor2_1
XFILLER_126_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_955 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12324_ _22703_/Q vssd1 vssd1 vccd1 vccd1 _12324_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14137__A2 _14561_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16092_ _16072_/X _16084_/Y _16086_/Y vssd1 vssd1 vccd1 vccd1 _16092_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_1018 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12913__B _20972_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22604__A0 _18115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19920_ _19881_/A _19823_/A _19875_/A vssd1 vssd1 vccd1 vccd1 _19920_/Y sky130_fd_sc_hd__a21oi_1
X_12255_ _18261_/A _18261_/B vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15043_ _14845_/B _15175_/C _15175_/D vssd1 vssd1 vccd1 vccd1 _15044_/B sky130_fd_sc_hd__o21ai_1
XFILLER_79_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13728__C _14834_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19851_ _19851_/A _19851_/B vssd1 vssd1 vccd1 vccd1 _19909_/C sky130_fd_sc_hd__nand2_1
XFILLER_123_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12186_ _12177_/B _12177_/C _12177_/A vssd1 vssd1 vccd1 vccd1 _12186_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_122_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18802_ _18613_/B _18797_/Y _19052_/A _18801_/Y vssd1 vssd1 vccd1 vccd1 _18804_/A
+ sky130_fd_sc_hd__o22ai_1
X_19782_ _19782_/A _19782_/B vssd1 vssd1 vccd1 vccd1 _19787_/B sky130_fd_sc_hd__nor2_1
X_16994_ _17087_/A _17087_/B vssd1 vssd1 vccd1 vccd1 _16994_/Y sky130_fd_sc_hd__nand2_2
XFILLER_62_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18733_ _18741_/C _18724_/A _18725_/A vssd1 vssd1 vccd1 vccd1 _18736_/A sky130_fd_sc_hd__a21bo_1
XFILLER_49_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15945_ _15945_/A _15945_/B _15945_/C vssd1 vssd1 vccd1 vccd1 _16024_/C sky130_fd_sc_hd__and3_1
XFILLER_62_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21019__A _21019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20918__B1 _17460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18664_ _19346_/A _18664_/B _19013_/C vssd1 vssd1 vccd1 vccd1 _18664_/X sky130_fd_sc_hd__and3_1
XFILLER_36_314 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15876_ _15864_/C _15864_/D _15862_/A vssd1 vssd1 vccd1 vccd1 _15876_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17615_ _17719_/A _17719_/C vssd1 vssd1 vccd1 vccd1 _17615_/X sky130_fd_sc_hd__or2_1
XFILLER_97_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14827_ _14826_/C _14916_/A _14826_/A vssd1 vssd1 vccd1 vccd1 _14828_/C sky130_fd_sc_hd__a21o_1
XFILLER_92_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18595_ _18595_/A _18595_/B _22912_/Q vssd1 vssd1 vccd1 vccd1 _18596_/B sky130_fd_sc_hd__nand3_1
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18328__A _18328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17546_ _12234_/X _12237_/X _17423_/X _17424_/X vssd1 vssd1 vccd1 vccd1 _17546_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14758_ _14758_/A _14758_/B _14758_/C vssd1 vssd1 vccd1 vccd1 _14758_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__17011__A1 _17006_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14575__B _14575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13709_ _13709_/A vssd1 vssd1 vccd1 vccd1 _14203_/B sky130_fd_sc_hd__clkbuf_2
X_17477_ _17318_/B _17318_/A _17467_/X _17466_/B vssd1 vssd1 vccd1 vccd1 _17479_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_177_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14689_ _14688_/Y _14685_/Y _14686_/X vssd1 vssd1 vccd1 vccd1 _14689_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_60_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19216_ _19507_/D _19496_/A vssd1 vssd1 vccd1 vccd1 _19216_/Y sky130_fd_sc_hd__nand2_1
X_16428_ _16431_/C vssd1 vssd1 vccd1 vccd1 _16652_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14376__A2 _14370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20593__A _20593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19147_ _19147_/A vssd1 vssd1 vccd1 vccd1 _19147_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16359_ _20854_/B vssd1 vssd1 vccd1 vccd1 _17833_/C sky130_fd_sc_hd__buf_2
XFILLER_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18511__A1 _19614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11595__C1 _18131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18511__B2 _19351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21110__A3 _21086_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19078_ _19098_/C _19097_/C vssd1 vssd1 vccd1 vccd1 _19106_/C sky130_fd_sc_hd__nand2_1
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18029_ _21086_/D _18030_/B _20012_/A _18029_/D vssd1 vssd1 vccd1 vccd1 _18029_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_160_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21040_ _21076_/C _21076_/D vssd1 vssd1 vccd1 vccd1 _21041_/B sky130_fd_sc_hd__nand2_1
XFILLER_160_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17407__A _17407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13639__B2 _21938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13654__B _21874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12847__C1 _20129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11455__A _18203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21942_ _22045_/A _22045_/B vssd1 vssd1 vccd1 vccd1 _21952_/A sky130_fd_sc_hd__or2_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21873_ _21742_/B _21939_/A _22057_/B _22173_/B _21972_/A vssd1 vssd1 vccd1 vccd1
+ _21875_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14766__A _14911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15261__B1 _15205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _20890_/A _20891_/A _20830_/B _20830_/A vssd1 vssd1 vccd1 vccd1 _20840_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_70_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11822__B1 _11762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20755_ _20658_/Y _20660_/A _20659_/Y vssd1 vssd1 vccd1 vccd1 _20755_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_168_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16761__B1 _16759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20686_ _20686_/A vssd1 vssd1 vccd1 vccd1 _20717_/A sky130_fd_sc_hd__clkbuf_2
X_22425_ _22425_/A vssd1 vssd1 vccd1 vccd1 _22712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15316__A1 _15326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22356_ _22356_/A _22356_/B _22356_/C vssd1 vssd1 vccd1 vccd1 _22358_/A sky130_fd_sc_hd__and3_1
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13327__B1 _13326_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21307_ _21307_/A _21307_/B _21307_/C vssd1 vssd1 vccd1 vccd1 _21312_/C sky130_fd_sc_hd__nand3_1
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22287_ _22684_/Q _22289_/B vssd1 vssd1 vccd1 vccd1 _22325_/A sky130_fd_sc_hd__nand2_1
XFILLER_163_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12040_ _22962_/Q vssd1 vssd1 vccd1 vccd1 _22660_/B sky130_fd_sc_hd__buf_2
XANTENNA__17069__A1 _22893_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21238_ _21237_/Y _21238_/B _21238_/C vssd1 vssd1 vccd1 vccd1 _21239_/C sky130_fd_sc_hd__nand3b_1
XFILLER_85_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17317__A _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20612__A2 _15723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21169_ _21169_/A _22852_/Q vssd1 vssd1 vccd1 vccd1 _21701_/A sky130_fd_sc_hd__and2_1
XFILLER_133_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13991_ _13877_/B _14468_/A _13986_/Y _13987_/X vssd1 vssd1 vccd1 vccd1 _13992_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_59_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _15406_/X _15404_/X _15403_/A vssd1 vssd1 vccd1 vccd1 _15731_/A sky130_fd_sc_hd__o21ai_1
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12942_ _15774_/D _12981_/B _20584_/C _12941_/X vssd1 vssd1 vccd1 vccd1 _12942_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20678__A _20678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20915__A3 _17460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _15507_/X _15601_/Y _15502_/C vssd1 vssd1 vccd1 vccd1 _15662_/C sky130_fd_sc_hd__o21ai_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _12873_/A vssd1 vssd1 vccd1 vccd1 _20169_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17400_ _17400_/A vssd1 vssd1 vccd1 vccd1 _17400_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16594__C _16594_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _13820_/X _13821_/Y _13950_/X _13823_/Y vssd1 vssd1 vccd1 vccd1 _14612_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18380_ _18520_/A _18726_/A _18520_/B vssd1 vssd1 vccd1 vccd1 _18381_/C sky130_fd_sc_hd__nand3_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _11698_/X _11700_/Y _11816_/Y _11823_/Y vssd1 vssd1 vccd1 vccd1 _12083_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15592_ _15588_/Y _16216_/A _16253_/B _15543_/Y vssd1 vssd1 vccd1 vccd1 _16287_/A
+ sky130_fd_sc_hd__a22oi_2
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12605__A2 _15799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16900__B1_N _22894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17331_ _17331_/A vssd1 vssd1 vccd1 vccd1 _17331_/Y sky130_fd_sc_hd__inv_2
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _14099_/B _14096_/C _14099_/C vssd1 vssd1 vccd1 vccd1 _14544_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__12196__A _22961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ _11755_/A _19461_/A _18303_/C vssd1 vssd1 vccd1 vccd1 _11755_/Y sky130_fd_sc_hd__nand3_1
XFILLER_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17262_ _17298_/A _17298_/B _17298_/C vssd1 vssd1 vccd1 vccd1 _17262_/X sky130_fd_sc_hd__and3_1
X_14474_ _14467_/X _14143_/X _14462_/Y _14461_/Y vssd1 vssd1 vccd1 vccd1 _14478_/B
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__16752__B1 _16599_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11686_ _11685_/X _11673_/X _11674_/A vssd1 vssd1 vccd1 vccd1 _11687_/B sky130_fd_sc_hd__a21boi_2
XFILLER_146_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19001_ _19000_/Y _18986_/Y _18991_/Y _18881_/X vssd1 vssd1 vccd1 vccd1 _19001_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_186_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16213_ _16213_/A vssd1 vssd1 vccd1 vccd1 _16213_/Y sky130_fd_sc_hd__inv_2
X_13425_ _13401_/A _13265_/A _13262_/D _13262_/A vssd1 vssd1 vccd1 vccd1 _13438_/A
+ sky130_fd_sc_hd__a22o_1
X_17193_ _17187_/X _17191_/Y _17192_/X vssd1 vssd1 vccd1 vccd1 _17193_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__19297__A2 _18023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15300__A _18107_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15307__A1 _12500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16144_ _16137_/C _16137_/A _16137_/B _16143_/Y vssd1 vssd1 vccd1 vccd1 _16145_/C
+ sky130_fd_sc_hd__a31o_1
X_13356_ _13122_/C _13122_/A _13122_/B _13141_/A _13166_/Y vssd1 vssd1 vccd1 vccd1
+ _13358_/B sky130_fd_sc_hd__a32oi_1
XFILLER_155_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ _20130_/A _12904_/A _20461_/C vssd1 vssd1 vccd1 vccd1 _12307_/Y sky130_fd_sc_hd__nand3_1
X_16075_ _11845_/X _20728_/B _15907_/Y _15993_/Y _16130_/A vssd1 vssd1 vccd1 vccd1
+ _16075_/X sky130_fd_sc_hd__o221a_1
X_13287_ _13340_/A _13286_/B _13223_/Y _13225_/X vssd1 vssd1 vccd1 vccd1 _13288_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19903_ _19901_/X _19902_/X _19846_/B _19850_/B vssd1 vssd1 vccd1 vccd1 _19905_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15026_ _15107_/C _15026_/B _15026_/C vssd1 vssd1 vccd1 vccd1 _15028_/A sky130_fd_sc_hd__and3_1
X_12238_ _12234_/X _12237_/X _18778_/A vssd1 vssd1 vccd1 vccd1 _12240_/A sky130_fd_sc_hd__a21o_1
XFILLER_111_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16807__A1 _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17227__A _17227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19834_ _19881_/A vssd1 vssd1 vccd1 vccd1 _19834_/Y sky130_fd_sc_hd__inv_2
X_12169_ _18162_/A _12175_/A _12164_/Y _12168_/X vssd1 vssd1 vccd1 vccd1 _12177_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__16131__A _16131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19765_ _19813_/A _19813_/B _19764_/Y vssd1 vssd1 vccd1 vccd1 _19765_/Y sky130_fd_sc_hd__a21oi_1
X_16977_ _15545_/X _15723_/X _16941_/X _16944_/Y _16934_/A vssd1 vssd1 vccd1 vccd1
+ _17158_/B sky130_fd_sc_hd__o221ai_4
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15491__B1 _15586_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 wb_adr_i[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_18716_ _18716_/A _19358_/C _19358_/D vssd1 vssd1 vccd1 vccd1 _18862_/B sky130_fd_sc_hd__and3_1
X_15928_ _15886_/Y _15917_/X _15927_/Y vssd1 vssd1 vccd1 vccd1 _15945_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__18984__C _19480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19696_ _19697_/D _19697_/B _19899_/A _17388_/X vssd1 vssd1 vccd1 vccd1 _19698_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18647_ _11819_/A _12010_/A _18536_/Y vssd1 vssd1 vccd1 vccd1 _18657_/A sky130_fd_sc_hd__o21ai_1
XFILLER_37_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15859_ _15859_/A _15859_/B _15859_/C _15859_/D vssd1 vssd1 vccd1 vccd1 _15861_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14046__A1 _14561_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18578_ _18578_/A _18578_/B _18578_/C vssd1 vssd1 vccd1 vccd1 _18774_/C sky130_fd_sc_hd__nand3_1
XANTENNA__15794__A1 _15918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22919__CLK _22922_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17529_ _17531_/D _17678_/A _15840_/X _17439_/X vssd1 vssd1 vccd1 vccd1 _17529_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20540_ _20843_/A _15890_/X _20393_/A vssd1 vssd1 vccd1 vccd1 _20540_/X sky130_fd_sc_hd__o21a_1
XANTENNA__22953__D _22953_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20471_ _20471_/A _20471_/B _20471_/C vssd1 vssd1 vccd1 vccd1 _20471_/Y sky130_fd_sc_hd__nand3_1
X_22210_ _22094_/A _22096_/X _22209_/Y _22290_/C vssd1 vssd1 vccd1 vccd1 _22211_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_195_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22141_ _22075_/X _22074_/Y _22138_/A _22138_/B _22079_/B vssd1 vssd1 vccd1 vccd1
+ _22159_/B sky130_fd_sc_hd__o2111ai_4
XANTENNA__19617__A _19772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22072_ _22072_/A _22072_/B vssd1 vssd1 vccd1 vccd1 _22073_/B sky130_fd_sc_hd__nand2_1
XANTENNA__19336__B _19619_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21023_ _21023_/A _21023_/B vssd1 vssd1 vccd1 vccd1 _21027_/A sky130_fd_sc_hd__xor2_1
XFILLER_101_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19460__A2 _15808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14809__B1 _14503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21925_ _22678_/Q _21925_/B vssd1 vssd1 vccd1 vccd1 _21925_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15785__A1 _11295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21856_ _21220_/X _21853_/X _21852_/Y _21850_/Y vssd1 vssd1 vccd1 vccd1 _21857_/C
+ sky130_fd_sc_hd__o211ai_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14993__C1 _14942_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20807_ _20178_/A _15935_/A _20806_/Y vssd1 vssd1 vccd1 vccd1 _20884_/B sky130_fd_sc_hd__o21a_1
X_21787_ _21846_/A _21846_/D vssd1 vssd1 vccd1 vccd1 _21787_/Y sky130_fd_sc_hd__nand2_1
XFILLER_169_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15537__A1 _14430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ _11333_/X _18367_/C _16058_/C _11521_/X vssd1 vssd1 vccd1 vccd1 _11644_/A
+ sky130_fd_sc_hd__a31o_2
XANTENNA__22863__D _22863_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20738_ _20738_/A _20738_/B _20738_/C vssd1 vssd1 vccd1 vccd1 _20738_/X sky130_fd_sc_hd__and3_1
Xclkbuf_4_2_0_bq_clk_i clkbuf_4_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _22933_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20664__C _20827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11471_ _11418_/A _11608_/A _11471_/C vssd1 vssd1 vccd1 vccd1 _11587_/A sky130_fd_sc_hd__nand3b_2
X_20669_ _20559_/A _20667_/Y _20770_/A _20666_/X vssd1 vssd1 vccd1 vccd1 _20670_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_167_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13210_ _13210_/A _13210_/B _13210_/C vssd1 vssd1 vccd1 vccd1 _13215_/A sky130_fd_sc_hd__and3_1
XFILLER_136_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22408_ _22408_/A vssd1 vssd1 vccd1 vccd1 _22704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ _14489_/C vssd1 vssd1 vccd1 vccd1 _14595_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11574__A2 _18629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13141_ _13141_/A vssd1 vssd1 vccd1 vccd1 _13286_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1059 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22339_ _22686_/Q _22347_/A vssd1 vssd1 vccd1 vccd1 _22346_/A sky130_fd_sc_hd__xor2_1
XFILLER_125_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13072_ _13145_/A vssd1 vssd1 vccd1 vccd1 _13097_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15774__B _15774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input56_A wb_dat_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16900_ _16899_/B _16899_/C _22894_/Q vssd1 vssd1 vccd1 vccd1 _17070_/A sky130_fd_sc_hd__a21bo_1
X_12023_ _11809_/A _11809_/B _11810_/C vssd1 vssd1 vccd1 vccd1 _12024_/B sky130_fd_sc_hd__o21ai_1
XFILLER_3_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17880_ _17880_/A vssd1 vssd1 vccd1 vccd1 _21044_/B sky130_fd_sc_hd__buf_2
XANTENNA__15493__C _16489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16831_ _16831_/A _16831_/B _16831_/C vssd1 vssd1 vccd1 vccd1 _16831_/X sky130_fd_sc_hd__and3_1
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19550_ _19454_/X _19455_/X _19545_/Y _19549_/Y vssd1 vssd1 vccd1 vccd1 _19555_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_111_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15790__A _20359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16762_ _16762_/A _16946_/A vssd1 vssd1 vccd1 vccd1 _16766_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19203__A2 _18814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13974_ _13974_/A vssd1 vssd1 vccd1 vccd1 _14963_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16017__A2 _13022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18501_ _11783_/A _18500_/Y _18099_/A vssd1 vssd1 vccd1 vccd1 _18698_/B sky130_fd_sc_hd__o21ai_4
X_15713_ _15713_/A vssd1 vssd1 vccd1 vccd1 _15775_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__21010__A2 _21048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19481_ _19481_/A vssd1 vssd1 vccd1 vccd1 _20012_/C sky130_fd_sc_hd__clkbuf_2
X_12925_ _12700_/Y _12705_/X _12950_/C vssd1 vssd1 vccd1 vccd1 _12926_/C sky130_fd_sc_hd__o21a_1
X_16693_ _16438_/A _16424_/A _16424_/B _16424_/C vssd1 vssd1 vccd1 vccd1 _16693_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_19_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18432_ _18432_/A _18432_/B _18432_/C vssd1 vssd1 vccd1 vccd1 _18434_/A sky130_fd_sc_hd__nand3_1
X_15644_ _15621_/X _15630_/X _15660_/C _15660_/A vssd1 vssd1 vccd1 vccd1 _15644_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _12856_/A _12856_/B _12856_/C vssd1 vssd1 vccd1 vccd1 _12857_/A sky130_fd_sc_hd__nand3_1
XFILLER_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12638__B _20853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _18363_/A _18363_/B vssd1 vssd1 vccd1 vccd1 _18471_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11591_/B _11591_/C _11591_/A vssd1 vssd1 vccd1 vccd1 _11807_/Y sky130_fd_sc_hd__a21oi_1
X_15575_ _18848_/D vssd1 vssd1 vccd1 vccd1 _19012_/D sky130_fd_sc_hd__clkbuf_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _12671_/A _12497_/A _12786_/Y vssd1 vssd1 vccd1 vccd1 _12788_/C sky130_fd_sc_hd__o21ai_2
X_17314_ _17313_/A _19482_/A _15887_/X _17007_/A vssd1 vssd1 vccd1 vccd1 _17520_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _13948_/X _13949_/X _14669_/A vssd1 vssd1 vccd1 vccd1 _14530_/A sky130_fd_sc_hd__a21o_1
X_18294_ _11818_/A _17635_/A _18200_/Y _18199_/Y vssd1 vssd1 vccd1 vccd1 _18294_/X
+ sky130_fd_sc_hd__o22a_1
X_11738_ _11738_/A vssd1 vssd1 vccd1 vccd1 _11738_/X sky130_fd_sc_hd__clkbuf_4
X_17245_ _17138_/X _17142_/X _17149_/B _17145_/Y vssd1 vssd1 vccd1 vccd1 _17255_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_159_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14457_ _14863_/C _22876_/Q vssd1 vssd1 vccd1 vccd1 _15205_/B sky130_fd_sc_hd__xor2_2
X_11669_ _15484_/A _11560_/C _11667_/Y _11668_/Y vssd1 vssd1 vccd1 vccd1 _11734_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__12654__A _16067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13408_ _21442_/A vssd1 vssd1 vccd1 vccd1 _21665_/D sky130_fd_sc_hd__clkbuf_2
X_17176_ _17173_/C _17173_/D _17175_/Y vssd1 vssd1 vccd1 vccd1 _17177_/C sky130_fd_sc_hd__a21o_1
XFILLER_162_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14388_ _22768_/Q _14330_/X _14379_/X _22736_/Q _14387_/X vssd1 vssd1 vccd1 vccd1
+ _14388_/X sky130_fd_sc_hd__a221o_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12373__B _20605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12762__A1 _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16127_ _16126_/Y _16122_/Y _12765_/X _16015_/X vssd1 vssd1 vccd1 vccd1 _16143_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_13339_ _13315_/X _13354_/B _13338_/Y vssd1 vssd1 vccd1 vccd1 _13339_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_116_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19690__A2 _19839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17883__C _21044_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16058_ _20249_/C _19000_/A _16058_/C _16100_/A vssd1 vssd1 vccd1 vccd1 _16080_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19156__B _19156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15009_ _14503_/X _14854_/X _15005_/Y _15007_/Y _15008_/X vssd1 vssd1 vccd1 vccd1
+ _15080_/A sky130_fd_sc_hd__o311a_1
XFILLER_69_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17453__A1 _17304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19817_ _19817_/A _19817_/B _19817_/C vssd1 vssd1 vccd1 vccd1 _19818_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11717__B _22658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19748_ _19658_/B _19658_/A _19814_/C _19670_/A vssd1 vssd1 vccd1 vccd1 _19760_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_84_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19679_ _19757_/A _19757_/B vssd1 vssd1 vccd1 vccd1 _22899_/D sky130_fd_sc_hd__xor2_1
XFILLER_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11733__A _15557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19900__A _19900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21710_ _21709_/X _21573_/B _21570_/A vssd1 vssd1 vccd1 vccd1 _21711_/B sky130_fd_sc_hd__o21a_1
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22690_ _22690_/CLK _22690_/D vssd1 vssd1 vccd1 vccd1 _22690_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21641_ _21641_/A vssd1 vssd1 vccd1 vccd1 _21654_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22891__CLK _22952_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21572_ _22674_/Q _21433_/A _21571_/Y vssd1 vssd1 vccd1 vccd1 _21573_/B sky130_fd_sc_hd__o21a_1
XFILLER_177_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20523_ _20403_/C _20403_/B _20403_/A vssd1 vssd1 vccd1 vccd1 _20526_/A sky130_fd_sc_hd__a21boi_1
XFILLER_193_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20454_ _20449_/Y _20454_/B _20454_/C vssd1 vssd1 vccd1 vccd1 _20532_/B sky130_fd_sc_hd__nand3b_1
XFILLER_137_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20781__A _20781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20385_ _20397_/A _20398_/A vssd1 vssd1 vccd1 vccd1 _20386_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22124_ _22128_/A _22219_/A _22128_/C vssd1 vssd1 vccd1 vccd1 _22124_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_134_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22055_ _21579_/A _21169_/A _21580_/B vssd1 vssd1 vccd1 vccd1 _22055_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13826__C _13826_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18610__A1_N _11877_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21006_ _21006_/A _21006_/B vssd1 vssd1 vccd1 vccd1 _21067_/D sky130_fd_sc_hd__nand2_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19984__A3 _20012_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16798__A3 _20255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22858__D _22858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12808__A2 _15335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22957_ _22964_/CLK _22957_/D vssd1 vssd1 vccd1 vccd1 _22957_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12710_ _12737_/A _12737_/B _12709_/Y vssd1 vssd1 vccd1 vccd1 _12710_/Y sky130_fd_sc_hd__a21oi_2
X_21908_ _22008_/A _22007_/A _21908_/C vssd1 vssd1 vccd1 vccd1 _21908_/X sky130_fd_sc_hd__and3_2
XFILLER_83_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13690_ _22752_/Q vssd1 vssd1 vccd1 vccd1 _13707_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16955__B1 _16947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22888_ _22915_/CLK input71/X vssd1 vssd1 vccd1 vccd1 _22888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11362__B _22786_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12641_ _12668_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _12745_/C sky130_fd_sc_hd__nand2_1
X_21839_ _21781_/C _21781_/A _21781_/B _21799_/B vssd1 vssd1 vccd1 vccd1 _21899_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_93_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18157__C1 _19168_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19354__D1 _18197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20675__B _20675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15360_ _12288_/A _15362_/D _15369_/C _15370_/A vssd1 vssd1 vccd1 vccd1 _20341_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__20503__A1 _20359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ _12785_/B vssd1 vssd1 vccd1 vccd1 _16947_/A sky130_fd_sc_hd__buf_2
XFILLER_196_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14311_ _22586_/D _22514_/A _22586_/B vssd1 vssd1 vccd1 vccd1 _14410_/A sky130_fd_sc_hd__and3_1
X_11523_ _11285_/A _11285_/B _11295_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11578_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15291_ _22884_/Q _15288_/A _15288_/C vssd1 vssd1 vccd1 vccd1 _15292_/B sky130_fd_sc_hd__o21ai_1
XFILLER_184_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17030_ _17036_/A _17036_/B _17031_/C vssd1 vssd1 vccd1 vccd1 _17033_/A sky130_fd_sc_hd__a21o_1
XFILLER_144_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14242_ _14243_/A _14243_/B _14246_/A _14253_/A vssd1 vssd1 vccd1 vccd1 _14245_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_183_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11454_ _11454_/A vssd1 vssd1 vccd1 vccd1 _18203_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14173_ _14054_/Y _14055_/X _14089_/Y _14167_/X vssd1 vssd1 vccd1 vccd1 _14175_/B
+ sky130_fd_sc_hd__o22ai_1
X_11385_ _11273_/X _11421_/A _11385_/C vssd1 vssd1 vccd1 vccd1 _11386_/A sky130_fd_sc_hd__and3b_1
XFILLER_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19672__A2 _19294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13124_ _13577_/A _21341_/A _13105_/A _13300_/A vssd1 vssd1 vccd1 vccd1 _13322_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_194_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18981_ _19694_/D vssd1 vssd1 vccd1 vccd1 _19772_/B sky130_fd_sc_hd__buf_2
XFILLER_124_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11818__A _11818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17932_ _17932_/A _17932_/B vssd1 vssd1 vccd1 vccd1 _17932_/Y sky130_fd_sc_hd__xnor2_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _13055_/A vssd1 vssd1 vccd1 vccd1 _13057_/C sky130_fd_sc_hd__inv_2
XANTENNA__13736__C _13736_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12640__C _12742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ _12006_/A _12006_/B vssd1 vssd1 vccd1 vccd1 _12006_/Y sky130_fd_sc_hd__nand2_2
XFILLER_61_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17863_ _17800_/Y _18048_/C _17910_/B _17862_/Y vssd1 vssd1 vccd1 vccd1 _17863_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_39_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19602_ _19602_/A _19602_/B _19602_/C _19769_/B vssd1 vssd1 vccd1 vccd1 _19602_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16814_ _16479_/X _16513_/X _16474_/Y vssd1 vssd1 vccd1 vccd1 _16822_/A sky130_fd_sc_hd__a21oi_2
XFILLER_38_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17794_ _17866_/A _17794_/B vssd1 vssd1 vccd1 vccd1 _17795_/C sky130_fd_sc_hd__or2_1
XFILLER_4_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19188__B2 _19015_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19533_ _19379_/B _19369_/Y _19363_/Y _19356_/X vssd1 vssd1 vccd1 vccd1 _19538_/C
+ sky130_fd_sc_hd__o2bb2a_2
X_16745_ _16745_/A vssd1 vssd1 vccd1 vccd1 _17091_/A sky130_fd_sc_hd__clkbuf_2
X_13957_ _13957_/A _13957_/B _13957_/C vssd1 vssd1 vccd1 vccd1 _14034_/B sky130_fd_sc_hd__nand3_1
XFILLER_98_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19464_ _19464_/A vssd1 vssd1 vccd1 vccd1 _19839_/D sky130_fd_sc_hd__buf_2
X_12908_ _15558_/C vssd1 vssd1 vccd1 vccd1 _15988_/B sky130_fd_sc_hd__buf_2
X_16676_ _16702_/B _16663_/Y _16675_/Y vssd1 vssd1 vccd1 vccd1 _16700_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__15749__A1 _15479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13888_ _13807_/A _14118_/B _13984_/C _13808_/Y vssd1 vssd1 vccd1 vccd1 _13888_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_50_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18415_ _18415_/A _18415_/B _18415_/C vssd1 vssd1 vccd1 vccd1 _18416_/A sky130_fd_sc_hd__nand3_1
X_15627_ _20461_/B vssd1 vssd1 vccd1 vccd1 _20471_/B sky130_fd_sc_hd__clkbuf_2
X_19395_ _19344_/Y _19338_/X _19390_/Y _19389_/X _19458_/A vssd1 vssd1 vccd1 vccd1
+ _19399_/A sky130_fd_sc_hd__o221ai_1
XFILLER_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12839_ _16708_/A vssd1 vssd1 vccd1 vccd1 _16300_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18346_ _18355_/A vssd1 vssd1 vccd1 vccd1 _18726_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15558_ _18107_/B _18107_/C _15558_/C _20133_/B vssd1 vssd1 vccd1 vccd1 _15558_/Y
+ sky130_fd_sc_hd__nand4_4
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19360__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14509_ _13793_/Y _14869_/B _13815_/X _14503_/A vssd1 vssd1 vccd1 vccd1 _14629_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_159_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18277_ _18277_/A _18277_/B vssd1 vssd1 vccd1 vccd1 _18411_/A sky130_fd_sc_hd__nand2_1
XFILLER_175_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15489_ _15489_/A vssd1 vssd1 vccd1 vccd1 _16786_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_684 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17228_ _17370_/A _17370_/B vssd1 vssd1 vccd1 vccd1 _17228_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput30 wb_adr_i[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
Xinput41 wb_dat_i[15] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput52 wb_dat_i[25] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput63 wb_dat_i[6] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17159_ _16978_/B _17158_/Y _16978_/A vssd1 vssd1 vccd1 vccd1 _17181_/B sky130_fd_sc_hd__a21boi_1
Xinput74 x[3] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17674__A1 _19619_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20170_ _20170_/A _20170_/B _20170_/C vssd1 vssd1 vccd1 vccd1 _20181_/B sky130_fd_sc_hd__nand3_2
XANTENNA__17674__B2 _17431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19317__D _19317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12499__B1 _20255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11447__B _15435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21222__A2 _21220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19614__B _19614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15437__B1 _12211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22040__B _22106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22811_ _22813_/CLK _22811_/D vssd1 vssd1 vccd1 vccd1 _22811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17729__A2 _11672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12559__A _12769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11463__A _15888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19630__A _19630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22742_ _22742_/CLK _22742_/D vssd1 vssd1 vccd1 vccd1 _22742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20733__A1 _20928_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20733__B2 _20734_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16401__A2 _16400_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22673_ _22944_/CLK _22673_/D vssd1 vssd1 vccd1 vccd1 _22673_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18246__A _18246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21624_ _21624_/A _21624_/B vssd1 vssd1 vccd1 vccd1 _21624_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18154__A2 _12158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12974__A1 _20792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__B2 _13016_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12294__A _12294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21555_ _21553_/B _21553_/C _21553_/D _21553_/A vssd1 vssd1 vccd1 vccd1 _21838_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20506_ _20503_/Y _20505_/Y _20502_/X vssd1 vssd1 vccd1 vccd1 _20506_/Y sky130_fd_sc_hd__a21oi_1
X_21486_ _21486_/A vssd1 vssd1 vccd1 vccd1 _21874_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15101__C _15205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11529__A2 _15797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20437_ _20437_/A _20554_/A _20554_/D _20764_/A vssd1 vssd1 vccd1 vccd1 _20439_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12726__B2 _12716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16468__A2 _16842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20368_ _20368_/A vssd1 vssd1 vccd1 vccd1 _20511_/A sky130_fd_sc_hd__buf_2
XFILLER_134_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22107_ _22221_/A _22221_/B _22221_/C vssd1 vssd1 vccd1 vccd1 _22179_/A sky130_fd_sc_hd__nand3_2
XFILLER_121_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20299_ _20165_/Y _20175_/Y _20181_/B vssd1 vssd1 vccd1 vccd1 _20300_/C sky130_fd_sc_hd__a21boi_1
X_22038_ _22182_/B _22037_/A _22037_/B _22037_/C vssd1 vssd1 vccd1 vccd1 _22038_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18090__A1 _18116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ _15050_/C _15050_/A vssd1 vssd1 vccd1 vccd1 _14997_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15979__B2 _15978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17648__A2_N _19689_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ _13826_/C _13826_/A _13849_/C vssd1 vssd1 vccd1 vccd1 _13814_/A sky130_fd_sc_hd__nand3b_4
XFILLER_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16586__D _16879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ _14791_/A _14791_/B _22765_/Q vssd1 vssd1 vccd1 vccd1 _14792_/B sky130_fd_sc_hd__nand3_1
XANTENNA_input19_A wb_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16530_ _16530_/A _16530_/B _16530_/C _16530_/D vssd1 vssd1 vccd1 vccd1 _16530_/X
+ sky130_fd_sc_hd__and4_1
X_13742_ _13897_/A _13833_/B _13821_/A _13833_/C vssd1 vssd1 vccd1 vccd1 _13745_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16461_ _20086_/A vssd1 vssd1 vccd1 vccd1 _20608_/A sky130_fd_sc_hd__buf_4
X_13673_ _13647_/Y _13671_/Y _13672_/Y vssd1 vssd1 vccd1 vccd1 _13674_/C sky130_fd_sc_hd__o21ai_1
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18200_ _18200_/A _19351_/C _18453_/C vssd1 vssd1 vccd1 vccd1 _18200_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__18156__A _18156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15412_ _15412_/A vssd1 vssd1 vccd1 vccd1 _15919_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19180_ _19014_/X _19015_/Y _19017_/Y _19026_/B vssd1 vssd1 vccd1 vccd1 _19182_/C
+ sky130_fd_sc_hd__a2bb2o_2
X_12624_ _12624_/A vssd1 vssd1 vccd1 vccd1 _12745_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16392_ _15763_/Y _15683_/Y _15681_/D vssd1 vssd1 vccd1 vccd1 _16393_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__12414__B1 _12413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18131_ _18328_/A _18131_/B _18131_/C vssd1 vssd1 vccd1 vccd1 _18131_/X sky130_fd_sc_hd__and3_1
XFILLER_106_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15343_ _15343_/A vssd1 vssd1 vccd1 vccd1 _15343_/X sky130_fd_sc_hd__buf_2
XFILLER_40_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16156__A1 _15936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12555_ _12515_/A _12565_/A _12567_/A _12523_/A _22824_/Q vssd1 vssd1 vccd1 vccd1
+ _12557_/B sky130_fd_sc_hd__a32o_1
XFILLER_157_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18062_ _18036_/B _18061_/Y _18062_/C _18062_/D vssd1 vssd1 vccd1 vccd1 _18063_/B
+ sky130_fd_sc_hd__and4bb_1
X_11506_ _11506_/A vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__buf_2
XFILLER_184_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15274_ _22877_/Q _22878_/Q _15271_/B vssd1 vssd1 vccd1 vccd1 _15275_/B sky130_fd_sc_hd__o21ai_1
XFILLER_172_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12486_ _12683_/A vssd1 vssd1 vccd1 vccd1 _20486_/C sky130_fd_sc_hd__buf_2
X_17013_ _17009_/X _17011_/Y _17025_/C vssd1 vssd1 vccd1 vccd1 _17019_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__12717__A1 _15325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14225_ _15006_/B vssd1 vssd1 vccd1 vccd1 _15114_/D sky130_fd_sc_hd__buf_2
X_11437_ _22957_/Q vssd1 vssd1 vccd1 vccd1 _11438_/B sky130_fd_sc_hd__buf_4
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14156_ _14148_/Y _14149_/X _14147_/A _14147_/B vssd1 vssd1 vccd1 vccd1 _14163_/B
+ sky130_fd_sc_hd__o211ai_1
X_11368_ _15932_/A _18795_/A _11333_/X _11319_/Y vssd1 vssd1 vccd1 vccd1 _11477_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_112_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _22723_/Q _22722_/Q vssd1 vssd1 vccd1 vccd1 _13143_/A sky130_fd_sc_hd__nor2_2
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ _19137_/A _19138_/B _19138_/C _18964_/D vssd1 vssd1 vccd1 vccd1 _18965_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14085_/Y _14086_/X _14075_/Y _14076_/Y vssd1 vssd1 vccd1 vccd1 _14087_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_140_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11299_ _11420_/B vssd1 vssd1 vccd1 vccd1 _11299_/X sky130_fd_sc_hd__clkbuf_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _17915_/A _17915_/B vssd1 vssd1 vccd1 vccd1 _17970_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13038_ _13038_/A _13038_/B _13038_/C _13038_/D vssd1 vssd1 vccd1 vccd1 _13039_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__15962__B _20806_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18895_ _11636_/X _18889_/X _18890_/X _19695_/A _15888_/X vssd1 vssd1 vccd1 vccd1
+ _18895_/X sky130_fd_sc_hd__o32a_1
XFILLER_67_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17235__A _18200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17846_ _17860_/B vssd1 vssd1 vccd1 vccd1 _17857_/B sky130_fd_sc_hd__inv_2
XFILLER_14_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13175__B1_N _13465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17777_ _17785_/B _17954_/A _17777_/C vssd1 vssd1 vccd1 vccd1 _17778_/B sky130_fd_sc_hd__and3b_1
X_14989_ _14989_/A _14989_/B vssd1 vssd1 vccd1 vccd1 _22678_/D sky130_fd_sc_hd__nor2_1
XANTENNA__13445__A2 _13465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19516_ _19521_/D vssd1 vssd1 vccd1 vccd1 _19516_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11456__A1 _11727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16728_ _16325_/A _16325_/B _15932_/X _16727_/X vssd1 vssd1 vccd1 vccd1 _16732_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19447_ _19447_/A _19681_/B vssd1 vssd1 vccd1 vccd1 _19449_/A sky130_fd_sc_hd__nand2_1
X_16659_ _16659_/A _16659_/B _16659_/C vssd1 vssd1 vccd1 vccd1 _16673_/A sky130_fd_sc_hd__nand3_2
XFILLER_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12405__B1 _12687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19378_ _19356_/X _19363_/Y _19369_/Y _19374_/A _19374_/B vssd1 vssd1 vccd1 vccd1
+ _19378_/Y sky130_fd_sc_hd__o2111ai_4
XANTENNA__17401__C _17401_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12826__B _16322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18329_ _18322_/Y _18327_/Y _18529_/B vssd1 vssd1 vccd1 vccd1 _18354_/A sky130_fd_sc_hd__o21ai_2
XFILLER_31_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21340_ _21615_/A _21498_/D _21741_/B _21454_/A vssd1 vssd1 vccd1 vccd1 _21344_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_30_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20762__C _20827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21271_ _13419_/A _13416_/B _21270_/X vssd1 vssd1 vccd1 vccd1 _21281_/C sky130_fd_sc_hd__o21ai_1
XFILLER_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13381__A1 _21498_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20222_ _20222_/A vssd1 vssd1 vccd1 vccd1 _20457_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__13381__B2 _21741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18844__B1 _18862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15658__B1 _16062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__B1 _18984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20153_ _20143_/Y _20144_/Y _20125_/A vssd1 vssd1 vccd1 vccd1 _20197_/B sky130_fd_sc_hd__o21bai_1
XFILLER_170_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20084_ _12734_/X _16708_/X _20219_/A _20083_/X vssd1 vssd1 vccd1 vccd1 _20084_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_170_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11608__D _18115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16083__B1 _12765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_816 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_592 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19021__B1 _19194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20706__A1 _17423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20986_ _20986_/A _20985_/Y vssd1 vssd1 vccd1 vccd1 _20987_/B sky130_fd_sc_hd__or2b_1
XANTENNA__19572__A1 _22917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11998__A2 _11988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22725_ _22725_/CLK _22725_/D vssd1 vssd1 vccd1 vccd1 _22725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_595 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22656_ _22815_/Q input59/X _22656_/S vssd1 vssd1 vccd1 vccd1 _22657_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14936__A2 _14861_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17311__C _17311_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19324__A1 _12111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16208__B _16402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21607_ _21607_/A vssd1 vssd1 vccd1 vccd1 _21607_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21131__A1 _22942_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22587_ _22643_/A vssd1 vssd1 vccd1 vccd1 _22656_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12340_ _12340_/A _12822_/A _12822_/B _12340_/D vssd1 vssd1 vccd1 vccd1 _12341_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_138_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21538_ _21538_/A _21538_/B vssd1 vssd1 vccd1 vccd1 _21538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12271_ _12369_/A vssd1 vssd1 vccd1 vccd1 _12519_/B sky130_fd_sc_hd__buf_2
X_21469_ _13112_/Y _21469_/B _21583_/B _21583_/C vssd1 vssd1 vccd1 vccd1 _21578_/A
+ sky130_fd_sc_hd__nand4b_1
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13372__A1 _21185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14010_ _14033_/A _14033_/B _14033_/C vssd1 vssd1 vccd1 vccd1 _14523_/A sky130_fd_sc_hd__nand3_2
XANTENNA__17638__A1 _12234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21434__A2 _22673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17039__B _17840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12580__C1 _20101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17981__C _19983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15961_ _17645_/D vssd1 vssd1 vccd1 vccd1 _17643_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21198__A1 _13662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14679__A _14868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17700_ _17701_/A _17701_/B _17701_/C vssd1 vssd1 vccd1 vccd1 _17702_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13583__A _21195_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14912_ _14912_/A _14912_/B vssd1 vssd1 vccd1 vccd1 _14972_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11686__A1 _11685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15892_ _12772_/A _12774_/A _11504_/X _11505_/X _11506_/A vssd1 vssd1 vccd1 vccd1
+ _15900_/B sky130_fd_sc_hd__o221ai_4
X_18680_ _12154_/Y _18857_/A _18858_/A _18680_/D vssd1 vssd1 vccd1 vccd1 _18681_/A
+ sky130_fd_sc_hd__nand4b_2
XFILLER_75_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17631_ _17631_/A vssd1 vssd1 vccd1 vccd1 _17632_/A sky130_fd_sc_hd__buf_2
XANTENNA__15416__A3 _15350_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14843_ _14843_/A _14843_/B _14843_/C vssd1 vssd1 vccd1 vccd1 _14929_/A sky130_fd_sc_hd__nand3_1
XFILLER_76_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17562_ _17442_/A _16737_/X _16016_/X _16746_/X vssd1 vssd1 vccd1 vccd1 _17562_/Y
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__12096__D1 _11583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ _14775_/D _14571_/X _14869_/C _14791_/A _14791_/B vssd1 vssd1 vccd1 vccd1
+ _14859_/A sky130_fd_sc_hd__o2111ai_4
X_11986_ _11986_/A vssd1 vssd1 vccd1 vccd1 _11986_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15006__C _15006_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19301_ _19301_/A _19301_/B _19301_/C _19301_/D vssd1 vssd1 vccd1 vccd1 _19301_/Y
+ sky130_fd_sc_hd__nand4_1
X_16513_ _16513_/A vssd1 vssd1 vccd1 vccd1 _16513_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13725_ _13725_/A _13733_/B vssd1 vssd1 vccd1 vccd1 _13725_/Y sky130_fd_sc_hd__nand2_4
X_17493_ _17493_/A vssd1 vssd1 vccd1 vccd1 _17600_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15514__A1_N _15397_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16444_ _16444_/A vssd1 vssd1 vccd1 vccd1 _16444_/Y sky130_fd_sc_hd__inv_2
X_19232_ _19074_/B _19074_/C _19074_/D _19231_/X vssd1 vssd1 vccd1 vccd1 _19246_/B
+ sky130_fd_sc_hd__a31oi_4
X_13656_ _13657_/A _13657_/B _13657_/C vssd1 vssd1 vccd1 vccd1 _13658_/A sky130_fd_sc_hd__a21o_1
XFILLER_143_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22952__CLK _22952_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19163_ _11636_/X _19517_/A _18493_/A _15888_/X vssd1 vssd1 vccd1 vccd1 _19163_/X
+ sky130_fd_sc_hd__o22a_1
X_12607_ _12607_/A vssd1 vssd1 vccd1 vccd1 _12607_/X sky130_fd_sc_hd__clkbuf_2
X_16375_ _16366_/Y _16370_/Y _16374_/Y vssd1 vssd1 vccd1 vccd1 _16636_/A sky130_fd_sc_hd__a21oi_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13587_ _21445_/C _21489_/A _13586_/Y _13528_/X vssd1 vssd1 vccd1 vccd1 _13587_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18114_ _18279_/A _18278_/A _18184_/B vssd1 vssd1 vccd1 vccd1 _18114_/X sky130_fd_sc_hd__and3_1
XFILLER_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ _15326_/A vssd1 vssd1 vccd1 vccd1 _15326_/X sky130_fd_sc_hd__buf_4
XFILLER_184_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19094_ _19004_/Y _19010_/X _19028_/X _19032_/Y vssd1 vssd1 vccd1 vccd1 _19095_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__20476__A3 _12680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12538_ _22824_/Q vssd1 vssd1 vccd1 vccd1 _12548_/A sky130_fd_sc_hd__inv_2
XFILLER_9_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18045_ _18045_/A _18045_/B vssd1 vssd1 vccd1 vccd1 _18045_/Y sky130_fd_sc_hd__nand2_1
X_15257_ _15257_/A _15266_/B vssd1 vssd1 vccd1 vccd1 _15259_/B sky130_fd_sc_hd__xor2_1
XFILLER_172_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12662__A _12913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12469_ _12469_/A vssd1 vssd1 vccd1 vccd1 _12543_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14208_ _14259_/A _14259_/B _14261_/C _14207_/Y vssd1 vssd1 vccd1 vccd1 _14267_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22622__A1 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15188_ _15188_/A _15188_/B _15240_/C _15212_/A vssd1 vssd1 vccd1 vccd1 _15189_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_153_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_bq_clk_i clkbuf_3_7_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _22952_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11913__A2 _15936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14139_ _14154_/B _14154_/C vssd1 vssd1 vccd1 vccd1 _14239_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19996_ _19952_/B _19991_/B _19955_/B _19955_/A vssd1 vssd1 vccd1 vccd1 _19998_/A
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__11709__C _16257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16301__B2 _17443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16852__A2 _16853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18947_ _18952_/A _18952_/B _18946_/X vssd1 vssd1 vccd1 vccd1 _18951_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21189__A1 _21473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18878_ _18492_/A _18875_/Y _18881_/A vssd1 vssd1 vccd1 vccd1 _18880_/A sky130_fd_sc_hd__o21ai_1
XFILLER_95_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17829_ _17755_/A _17755_/B _17746_/X _17753_/Y vssd1 vssd1 vccd1 vccd1 _17831_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14076__C1 _14270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20840_ _20840_/A _20840_/B vssd1 vssd1 vccd1 vccd1 _20994_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11444__C _16711_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17014__C1 _17008_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21215__A _21724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20771_ _20772_/B _20772_/C _20772_/D _20772_/A vssd1 vssd1 vccd1 vccd1 _20773_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17565__B1 _16276_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12837__A _20130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15213__A _15213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22510_ _22750_/Q input58/X _22512_/S vssd1 vssd1 vccd1 vccd1 _22511_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19306__A1 _11345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19306__B2 _18371_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22441_ input68/X input67/X input34/X vssd1 vssd1 vccd1 vccd1 _22586_/C sky130_fd_sc_hd__and3_1
XFILLER_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22372_ _12876_/X input35/X _22380_/S vssd1 vssd1 vccd1 vccd1 _22373_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21323_ _21466_/A _21482_/A vssd1 vssd1 vccd1 vccd1 _21323_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15375__A2_N _15665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15586__C _15586_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21254_ _21990_/B _21299_/B _21260_/B vssd1 vssd1 vccd1 vccd1 _21254_/X sky130_fd_sc_hd__and3_1
XANTENNA__22613__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18293__A1 _16940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20205_ _20107_/A _20107_/B _20107_/C _20119_/C _20119_/D vssd1 vssd1 vccd1 vccd1
+ _20205_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_143_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21185_ _21185_/A vssd1 vssd1 vccd1 vccd1 _21185_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11619__C _18115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20136_ _12838_/B _20126_/Y _20132_/X _20142_/B _20142_/A vssd1 vssd1 vccd1 vccd1
+ _20155_/C sky130_fd_sc_hd__o2111ai_4
XANTENNA__14499__A _14611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_930 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11916__A _18459_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20067_ _22930_/Q vssd1 vssd1 vccd1 vccd1 _20191_/A sky130_fd_sc_hd__inv_2
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22825__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16056__B1 _15972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11840_ _11840_/A vssd1 vssd1 vccd1 vccd1 _11902_/B sky130_fd_sc_hd__clkbuf_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _18319_/B vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__buf_4
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ _20969_/A vssd1 vssd1 vccd1 vccd1 _20969_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11651__A _11942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ _13237_/X _13601_/A _13506_/C _13526_/A _13509_/X vssd1 vssd1 vccd1 vccd1
+ _13552_/A sky130_fd_sc_hd__o221a_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18137__C _18876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22708_ _22804_/CLK _22708_/D vssd1 vssd1 vccd1 vccd1 _22708_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14909__A2 _13736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14490_ _14857_/A _14494_/D _14626_/A _14494_/B vssd1 vssd1 vccd1 vccd1 _14490_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13441_ _13546_/A _13546_/B vssd1 vssd1 vccd1 vccd1 _13501_/A sky130_fd_sc_hd__xor2_1
X_22639_ _22807_/Q input50/X _22641_/S vssd1 vssd1 vccd1 vccd1 _22640_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0_0_bq_clk_i_A clkbuf_3_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18505__C1 _18698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16880__C _17039_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16160_ _16160_/A _16997_/C _16160_/C _16166_/B vssd1 vssd1 vccd1 vccd1 _16174_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_142_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13372_ _21185_/A _13067_/A _13202_/A vssd1 vssd1 vccd1 vccd1 _13373_/B sky130_fd_sc_hd__o21ai_2
XFILLER_182_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15111_ _15111_/A _15111_/B vssd1 vssd1 vccd1 vccd1 _15112_/B sky130_fd_sc_hd__nor2_1
XFILLER_155_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12323_ _12307_/Y _12314_/Y _12322_/X vssd1 vssd1 vccd1 vccd1 _12323_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16091_ _15936_/X _20728_/B _15988_/Y _16011_/B vssd1 vssd1 vccd1 vccd1 _16190_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__12482__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15042_ _15175_/D _15176_/A _15175_/C vssd1 vssd1 vccd1 vccd1 _15044_/A sky130_fd_sc_hd__or3_1
X_12254_ _12249_/A _18241_/B _12251_/A vssd1 vssd1 vccd1 vccd1 _18261_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22604__A1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19850_ _19850_/A _19850_/B _19850_/C vssd1 vssd1 vccd1 vccd1 _19851_/B sky130_fd_sc_hd__nand3_2
XANTENNA__18284__A1 _12204_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12185_ _12181_/B _12181_/C _12181_/A vssd1 vssd1 vccd1 vccd1 _12185_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16295__B1 _12094_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18801_ _12170_/X _12171_/X _12202_/A _12202_/B vssd1 vssd1 vccd1 vccd1 _18801_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_19781_ _19781_/A _19781_/B vssd1 vssd1 vccd1 vccd1 _19784_/A sky130_fd_sc_hd__nand2_1
XFILLER_150_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16993_ _11904_/X _11905_/X _20854_/A _20854_/B vssd1 vssd1 vccd1 vccd1 _17087_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_27_1150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18732_ _18729_/Y _18730_/Y _18731_/X vssd1 vssd1 vccd1 vccd1 _18732_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_62_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15944_ _15944_/A _15944_/B _15944_/C vssd1 vssd1 vccd1 vccd1 _15945_/A sky130_fd_sc_hd__nand3_1
XANTENNA__21019__B _21019_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15875_ _15875_/A _15875_/B vssd1 vssd1 vccd1 vccd1 _15875_/Y sky130_fd_sc_hd__nand2_1
X_18663_ _18663_/A vssd1 vssd1 vccd1 vccd1 _19346_/A sky130_fd_sc_hd__buf_2
XFILLER_36_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17614_ _17608_/X _17610_/Y _17722_/A vssd1 vssd1 vccd1 vccd1 _17720_/A sky130_fd_sc_hd__a21boi_1
X_14826_ _14826_/A _14916_/A _14826_/C vssd1 vssd1 vccd1 vccd1 _14828_/B sky130_fd_sc_hd__nand3_1
XFILLER_92_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12608__B1 _12450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18594_ _18595_/A _18595_/B _22912_/Q vssd1 vssd1 vccd1 vccd1 _18970_/A sky130_fd_sc_hd__a21o_1
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _17529_/X _17531_/X _17541_/Y _17544_/Y vssd1 vssd1 vccd1 vccd1 _17552_/A
+ sky130_fd_sc_hd__o211ai_1
X_14757_ _14752_/X _14757_/B vssd1 vssd1 vccd1 vccd1 _14761_/A sky130_fd_sc_hd__and2b_1
XANTENNA__17547__B1 _17546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ _11969_/A _12126_/A vssd1 vssd1 vccd1 vccd1 _12137_/A sky130_fd_sc_hd__nand2_2
XANTENNA__16129__A _16129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11561__A _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17011__A2 _17008_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ _14258_/B _14258_/D vssd1 vssd1 vccd1 vccd1 _13709_/A sky130_fd_sc_hd__nor2_1
X_17476_ _17301_/A _17301_/B _17301_/C _17486_/C vssd1 vssd1 vccd1 vccd1 _17476_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_149_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14688_ _14688_/A _14785_/B _14693_/B _14693_/A vssd1 vssd1 vccd1 vccd1 _14688_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_32_554 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19215_ _19215_/A vssd1 vssd1 vccd1 vccd1 _19215_/X sky130_fd_sc_hd__clkbuf_2
X_16427_ _16209_/A _16402_/B _16403_/A vssd1 vssd1 vccd1 vccd1 _16432_/A sky130_fd_sc_hd__a21boi_1
X_13639_ _13664_/B _22062_/A _13664_/D _21938_/B vssd1 vssd1 vccd1 vccd1 _13640_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19146_ _22914_/Q _18967_/B _19290_/A _19142_/B _19143_/Y vssd1 vssd1 vccd1 vccd1
+ _19290_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_157_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16358_ _20471_/B vssd1 vssd1 vccd1 vccd1 _20854_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_145_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11595__B1 _18131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15309_ _15309_/A _15309_/B vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16522__A1 _16248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19077_ _18825_/A _18825_/B _18824_/X vssd1 vssd1 vccd1 vccd1 _19097_/C sky130_fd_sc_hd__a21o_1
X_16289_ _16595_/A _16596_/A _16595_/B vssd1 vssd1 vccd1 vccd1 _16289_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_161_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18028_ _18028_/A vssd1 vssd1 vccd1 vccd1 _18029_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16799__A _17379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13887__A2 _14013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__A1 _11899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22848__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19979_ _19891_/Y _19974_/Y _19978_/Y vssd1 vssd1 vccd1 vccd1 _20057_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__17407__B _18303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13639__A2 _22062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22359__B1 _22352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14112__A _14112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12847__B1 _20250_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19775__B2 _19839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21941_ _22182_/A _22062_/A _22182_/C vssd1 vssd1 vccd1 vccd1 _22045_/B sky130_fd_sc_hd__nand3_1
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17423__A _17423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21872_ _21872_/A vssd1 vssd1 vccd1 vccd1 _22173_/B sky130_fd_sc_hd__buf_2
XFILLER_131_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15261__A1 _15230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20790__C1 _17462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14766__B _15082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ _20890_/B _20890_/C vssd1 vssd1 vccd1 vccd1 _20830_/B sky130_fd_sc_hd__nand2_1
XFILLER_78_1070 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20137__A2 _20126_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16039__A _16039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12567__A _12567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11822__A1 _18778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20754_ _20754_/A _20754_/B _20754_/C vssd1 vssd1 vccd1 vccd1 _20759_/B sky130_fd_sc_hd__nand3_4
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16761__A1 _16225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20685_ _20685_/A vssd1 vssd1 vccd1 vccd1 _21009_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22424_ _22712_/Q input51/X _22424_/S vssd1 vssd1 vccd1 vccd1 _22425_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_570 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12783__C1 _15696_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15316__A2 _15325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22355_ _22355_/A vssd1 vssd1 vccd1 vccd1 _22356_/C sky130_fd_sc_hd__inv_2
XFILLER_137_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16205__C _16402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21306_ _21312_/A vssd1 vssd1 vccd1 vccd1 _21738_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22286_ _22286_/A vssd1 vssd1 vccd1 vccd1 _22289_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21237_ _21237_/A _21237_/B vssd1 vssd1 vccd1 vccd1 _21237_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_116_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16277__B1 _16276_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17317__B _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21168_ _21169_/A _22852_/Q vssd1 vssd1 vccd1 vccd1 _21700_/A sky130_fd_sc_hd__nor2_1
XFILLER_49_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15118__A _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20119_ _20119_/A _20119_/B _20119_/C _20119_/D vssd1 vssd1 vccd1 vccd1 _20121_/B
+ sky130_fd_sc_hd__nand4_2
X_13990_ _14013_/A _14013_/B _14786_/B vssd1 vssd1 vccd1 vccd1 _14468_/A sky130_fd_sc_hd__nand3_2
X_21099_ _21115_/A vssd1 vssd1 vccd1 vccd1 _21138_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ _16489_/A _15696_/D _12973_/A _13016_/C vssd1 vssd1 vccd1 vccd1 _12941_/X
+ sky130_fd_sc_hd__and4_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20678__B _20678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _15660_/A _15660_/B _15660_/C vssd1 vssd1 vccd1 vccd1 _15662_/B sky130_fd_sc_hd__nand3_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _12872_/A _12872_/B _12872_/C vssd1 vssd1 vccd1 vccd1 _12873_/A sky130_fd_sc_hd__nand3_1
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19518__A1 _17083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14611_/A _14611_/B _14611_/C _14611_/D vssd1 vssd1 vccd1 vccd1 _14636_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _11811_/Y _11815_/Y _11817_/Y _11822_/X vssd1 vssd1 vccd1 vccd1 _11823_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_57_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15591_ _15498_/B _15589_/X _16265_/B vssd1 vssd1 vccd1 vccd1 _16216_/A sky130_fd_sc_hd__a21o_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17529__B1 _15840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12605__A3 _20463_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17330_ _17485_/A _17330_/B _17485_/B vssd1 vssd1 vccd1 vccd1 _17330_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__11381__A _11633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14524_/Y _14535_/X _14536_/Y vssd1 vssd1 vccd1 vccd1 _14544_/B sky130_fd_sc_hd__o21ai_2
X_11754_ _17280_/A vssd1 vssd1 vccd1 vccd1 _19461_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11813__A1 _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20694__A _20694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12196__B _22962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _17268_/B vssd1 vssd1 vccd1 vccd1 _17298_/C sky130_fd_sc_hd__clkbuf_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14473_ _13987_/X _13984_/Y _14470_/X vssd1 vssd1 vccd1 vccd1 _14478_/A sky130_fd_sc_hd__a21oi_1
X_11685_ _18203_/A _18203_/B _15580_/A _16276_/A vssd1 vssd1 vccd1 vccd1 _11685_/X
+ sky130_fd_sc_hd__or4_4
X_16212_ _16422_/A _16204_/Y _16211_/Y vssd1 vssd1 vccd1 vccd1 _16212_/Y sky130_fd_sc_hd__a21oi_1
X_19000_ _19000_/A _19161_/A _19000_/C _19614_/C vssd1 vssd1 vccd1 vccd1 _19000_/Y
+ sky130_fd_sc_hd__nand4_4
X_13424_ _13424_/A vssd1 vssd1 vccd1 vccd1 _13546_/A sky130_fd_sc_hd__clkbuf_2
X_17192_ _17200_/B _17200_/C _17200_/A vssd1 vssd1 vccd1 vccd1 _17192_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16143_ _16143_/A _16143_/B _16143_/C vssd1 vssd1 vccd1 vccd1 _16143_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__15300__B _18107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13355_ _13349_/X _13351_/Y _13354_/Y vssd1 vssd1 vccd1 vccd1 _13358_/A sky130_fd_sc_hd__o21ai_1
XFILLER_155_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15307__A2 _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13318__A1 _13633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ _12348_/A vssd1 vssd1 vccd1 vccd1 _20461_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_154_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16074_ _12294_/A _12294_/B _16130_/A _16051_/C _15918_/X vssd1 vssd1 vccd1 vccd1
+ _16074_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_142_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13286_ _13340_/A _13286_/B _13286_/C _13286_/D vssd1 vssd1 vccd1 vccd1 _13288_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_170_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22589__A0 _18953_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19902_ _17873_/A _19981_/A _17876_/A _19987_/C vssd1 vssd1 vccd1 vccd1 _19902_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15025_ _15023_/Y _14951_/A _15024_/Y vssd1 vssd1 vccd1 vccd1 _15026_/B sky130_fd_sc_hd__a21boi_1
X_12237_ _15531_/A vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_107_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12940__A _20463_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19833_ _19833_/A vssd1 vssd1 vccd1 vccd1 _19881_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16807__A2 _15631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12168_ _11500_/Y _15887_/A _12167_/X _12163_/X _12156_/X vssd1 vssd1 vccd1 vccd1
+ _12168_/X sky130_fd_sc_hd__o311a_2
XFILLER_96_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19206__B1 _19211_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19764_ _19814_/A _19764_/B _19764_/C vssd1 vssd1 vccd1 vccd1 _19764_/Y sky130_fd_sc_hd__nand3b_1
X_16976_ _16976_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _17158_/A sky130_fd_sc_hd__nand2_1
X_12099_ _12117_/A _12096_/Y _12098_/Y vssd1 vssd1 vccd1 vccd1 _12099_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15491__A1 _12209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18715_ _18715_/A _18722_/D vssd1 vssd1 vccd1 vccd1 _18721_/A sky130_fd_sc_hd__nand2_1
X_15927_ _15967_/A _15967_/B _15967_/C vssd1 vssd1 vccd1 vccd1 _15927_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__18984__D _19481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 wb_adr_i[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_19695_ _19695_/A vssd1 vssd1 vccd1 vccd1 _19899_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13771__A _22872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18646_ _18646_/A _18646_/B _18646_/C vssd1 vssd1 vccd1 vccd1 _18646_/X sky130_fd_sc_hd__and3_1
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15858_ _15854_/A _15854_/B _15864_/B _15756_/X vssd1 vssd1 vccd1 vccd1 _15861_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__19509__A1 _19652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14809_ _14808_/B _14808_/C _14503_/A _14562_/X vssd1 vssd1 vccd1 vccd1 _14809_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18577_ _18576_/Y _18411_/B _18219_/B _18417_/C vssd1 vssd1 vccd1 vccd1 _18578_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15794__A2 _15792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15789_ _12413_/X _12576_/X _16058_/C _16192_/B _15960_/A vssd1 vssd1 vccd1 vccd1
+ _15834_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_33_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17528_ _17531_/B vssd1 vssd1 vccd1 vccd1 _17678_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17459_ _17479_/A _17479_/B vssd1 vssd1 vccd1 vccd1 _17470_/A sky130_fd_sc_hd__nand2_1
XFILLER_193_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20470_ _20495_/B _20495_/A _20468_/X _20469_/X vssd1 vssd1 vccd1 vccd1 _20470_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_119_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19129_ _19129_/A _19129_/B _19129_/C vssd1 vssd1 vccd1 vccd1 _19130_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13624__D_N _21866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17153__D1 _19504_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22140_ _22140_/A _22140_/B vssd1 vssd1 vccd1 vccd1 _22164_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21866__C _21866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22071_ _22131_/A _22196_/B _22132_/B _22135_/A vssd1 vssd1 vccd1 vccd1 _22073_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__16322__A _16322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18799__A2 _17388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21022_ _20980_/A _20980_/B _20985_/C vssd1 vssd1 vccd1 vccd1 _21023_/B sky130_fd_sc_hd__o21ai_2
XFILLER_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16976__B _16976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21924_ _21931_/A _21924_/B vssd1 vssd1 vccd1 vccd1 _21925_/B sky130_fd_sc_hd__xor2_1
XFILLER_55_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13245__B1 _21584_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21855_ _21850_/Y _21852_/Y _21854_/X vssd1 vssd1 vccd1 vccd1 _21857_/B sky130_fd_sc_hd__a21o_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15785__A2 _11295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _20806_/A _20806_/B _20806_/C vssd1 vssd1 vccd1 vccd1 _20806_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__14993__B1 _14942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21786_ _21846_/B _21846_/C vssd1 vssd1 vccd1 vccd1 _21786_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20737_ _20737_/A _20737_/B _20737_/C _20737_/D vssd1 vssd1 vccd1 vccd1 _20748_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_11_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11470_ _11587_/C vssd1 vssd1 vccd1 vccd1 _18093_/A sky130_fd_sc_hd__buf_2
XFILLER_13_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20668_ _20565_/Y _20566_/Y _20770_/A _20666_/X _20667_/Y vssd1 vssd1 vccd1 vccd1
+ _20670_/A sky130_fd_sc_hd__o221a_1
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22407_ _22704_/Q input42/X _22413_/S vssd1 vssd1 vccd1 vccd1 _22408_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_67 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20599_ _20599_/A _20599_/B vssd1 vssd1 vccd1 vccd1 _20599_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13140_ _13322_/B _13128_/X _13136_/Y _13139_/Y vssd1 vssd1 vccd1 vccd1 _13141_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_137_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22338_ _22338_/A _22338_/B vssd1 vssd1 vccd1 vccd1 _22347_/A sky130_fd_sc_hd__xnor2_1
XFILLER_164_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13071_ _22842_/Q vssd1 vssd1 vccd1 vccd1 _13519_/B sky130_fd_sc_hd__buf_2
XFILLER_2_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22269_ _22221_/C _22221_/A _22221_/B _22308_/B _22308_/C vssd1 vssd1 vccd1 vccd1
+ _22309_/A sky130_fd_sc_hd__a311o_1
XANTENNA__16232__A _16770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15774__C _15774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ _11972_/Y _11976_/Y _12006_/A _12006_/B _11986_/X vssd1 vssd1 vccd1 vccd1
+ _12025_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_78_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input49_A wb_dat_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16830_ _16828_/A _16828_/B _16831_/C vssd1 vssd1 vccd1 vccd1 _16830_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16761_ _16225_/A _16227_/A _16759_/A _17251_/A vssd1 vssd1 vccd1 vccd1 _16946_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_150_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13973_ _13973_/A _13973_/B vssd1 vssd1 vccd1 vccd1 _14475_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18500_ _18677_/A _18678_/C _18500_/C _18677_/C vssd1 vssd1 vccd1 vccd1 _18500_/Y
+ sky130_fd_sc_hd__nand4_4
X_15712_ _11462_/A _12727_/A _15406_/A vssd1 vssd1 vccd1 vccd1 _15713_/A sky130_fd_sc_hd__o21ai_1
X_12924_ _12611_/Y _12588_/Y _12608_/X vssd1 vssd1 vccd1 vccd1 _12926_/B sky130_fd_sc_hd__a21o_1
X_16692_ _16424_/B _16424_/C _16691_/Y vssd1 vssd1 vccd1 vccd1 _16692_/X sky130_fd_sc_hd__a21o_1
X_19480_ _19480_/A vssd1 vssd1 vccd1 vccd1 _20012_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21010__A3 _21048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18431_ _18601_/B _18601_/A _18430_/A _18600_/A vssd1 vssd1 vccd1 vccd1 _18432_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15643_ _15636_/Y _15640_/Y _15642_/X vssd1 vssd1 vccd1 vccd1 _15660_/A sky130_fd_sc_hd__a21o_1
X_12855_ _12855_/A _12855_/B _20120_/A _12859_/A vssd1 vssd1 vccd1 vccd1 _12856_/C
+ sky130_fd_sc_hd__nand4_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11806_ _11809_/A _11809_/B _11814_/A vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__12638__C _20972_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15574_ _17436_/A _16191_/A _15574_/C vssd1 vssd1 vccd1 vccd1 _15574_/X sky130_fd_sc_hd__and3_1
X_18362_ _18365_/A _18995_/A _18154_/X vssd1 vssd1 vccd1 vccd1 _18363_/B sky130_fd_sc_hd__o21ai_1
XFILLER_61_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12786_ _15559_/C _15559_/D _20130_/C vssd1 vssd1 vccd1 vccd1 _12786_/Y sky130_fd_sc_hd__nand3_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _17313_/A _17313_/B _19482_/A _17313_/D vssd1 vssd1 vccd1 vccd1 _17523_/A
+ sky130_fd_sc_hd__nand4_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _22874_/Q vssd1 vssd1 vccd1 vccd1 _14669_/A sky130_fd_sc_hd__inv_2
X_11737_ _11737_/A vssd1 vssd1 vccd1 vccd1 _11737_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ _16940_/X _19043_/A _18636_/A _12216_/X vssd1 vssd1 vccd1 vccd1 _18293_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14456_ _11667_/Y _22658_/A _14448_/A vssd1 vssd1 vccd1 vccd1 _22671_/D sky130_fd_sc_hd__a21oi_1
X_17244_ _17269_/B vssd1 vssd1 vccd1 vccd1 _17298_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11668_ _11668_/A _12210_/A vssd1 vssd1 vccd1 vccd1 _11668_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13407_ _22850_/Q vssd1 vssd1 vccd1 vccd1 _21442_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17175_ _17323_/A _17127_/A _17174_/Y vssd1 vssd1 vccd1 vccd1 _17175_/Y sky130_fd_sc_hd__a21oi_1
X_14387_ _22800_/Q _14381_/X _14382_/X _14331_/X _22704_/Q vssd1 vssd1 vccd1 vccd1
+ _14387_/X sky130_fd_sc_hd__a32o_1
X_11599_ _15932_/A _11598_/X _11793_/A _11528_/Y _11589_/X vssd1 vssd1 vccd1 vccd1
+ _11600_/C sky130_fd_sc_hd__o221ai_1
XFILLER_143_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16126_ _16126_/A _16126_/B _16126_/C vssd1 vssd1 vccd1 vccd1 _16126_/Y sky130_fd_sc_hd__nand3_1
X_13338_ _21234_/A _13338_/B vssd1 vssd1 vccd1 vccd1 _13338_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12762__A2 _12761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16057_ _11912_/A _15890_/A _15993_/Y vssd1 vssd1 vccd1 vccd1 _16080_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12670__A _12758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ _13272_/A _13272_/B _21632_/A _13572_/B _13268_/X vssd1 vssd1 vccd1 vccd1
+ _13269_/X sky130_fd_sc_hd__o2111a_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15008_ _15107_/A _15107_/B _15008_/C vssd1 vssd1 vccd1 vccd1 _15008_/X sky130_fd_sc_hd__and3_1
XFILLER_29_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19816_ _19658_/A _19658_/B _19747_/A _19746_/Y vssd1 vssd1 vccd1 vccd1 _19817_/C
+ sky130_fd_sc_hd__o31a_1
XANTENNA__15981__A _18512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16661__B1 _17502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19747_ _19747_/A _19746_/Y vssd1 vssd1 vccd1 vccd1 _19814_/C sky130_fd_sc_hd__or2b_1
XFILLER_38_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16959_ _16959_/A _16959_/B vssd1 vssd1 vccd1 vccd1 _16959_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19678_ _19452_/B _19574_/A _19574_/B _19452_/A _19677_/Y vssd1 vssd1 vccd1 vccd1
+ _19757_/B sky130_fd_sc_hd__a41oi_4
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18629_ _18629_/A _18629_/B vssd1 vssd1 vccd1 vccd1 _18629_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15205__B _15205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13778__A1 _13948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21640_ _21640_/A _21640_/B _21640_/C _21640_/D vssd1 vssd1 vccd1 vccd1 _21641_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_178_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21571_ _22674_/Q _21433_/A _21434_/Y _21294_/C vssd1 vssd1 vccd1 vccd1 _21571_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20522_ _20522_/A _20522_/B _20522_/C vssd1 vssd1 vccd1 vccd1 _20529_/A sky130_fd_sc_hd__nand3_1
XFILLER_193_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18469__A1 _18770_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20453_ _20723_/A _20734_/A _20335_/B _20335_/C _20447_/Y vssd1 vssd1 vccd1 vccd1
+ _20454_/C sky130_fd_sc_hd__a221o_2
XFILLER_107_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18532__A _18665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20781__B _20781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20276__A1 _12500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20384_ _20403_/A _20376_/A _20337_/A vssd1 vssd1 vccd1 vccd1 _20388_/A sky130_fd_sc_hd__a21o_1
XFILLER_161_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22123_ _22051_/Y _22054_/Y _22060_/X vssd1 vssd1 vccd1 vccd1 _22128_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__17148__A _20129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22054_ _22100_/C _22099_/B _22099_/A vssd1 vssd1 vccd1 vccd1 _22054_/Y sky130_fd_sc_hd__nand3_1
XFILLER_173_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15891__A _15891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21005_ _21004_/A _21004_/B _21076_/B vssd1 vssd1 vccd1 vccd1 _21041_/A sky130_fd_sc_hd__o21a_1
XANTENNA__18641__A1 _18619_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22956_ _22959_/CLK _22956_/D vssd1 vssd1 vccd1 vccd1 _22956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_700 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21907_ _22007_/B vssd1 vssd1 vccd1 vccd1 _21908_/C sky130_fd_sc_hd__inv_2
XFILLER_16_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22887_ _22952_/CLK input70/X vssd1 vssd1 vccd1 vccd1 _22887_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__16955__A1 _16225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _12640_/A _12640_/B _12742_/A vssd1 vssd1 vccd1 vccd1 _12668_/B sky130_fd_sc_hd__nand3_1
XFILLER_169_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21838_ _21838_/A _21838_/B vssd1 vssd1 vccd1 vccd1 _21917_/A sky130_fd_sc_hd__nor2_2
XANTENNA__19354__C1 _19496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12441__A1 _15558_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ _12571_/A _12571_/B vssd1 vssd1 vccd1 vccd1 _12785_/B sky130_fd_sc_hd__nand2_1
X_21769_ _21769_/A _21769_/B vssd1 vssd1 vccd1 vccd1 _21769_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12441__B2 _20456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16227__A _16227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _14310_/A vssd1 vssd1 vccd1 vccd1 _22586_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_196_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _11333_/A _18445_/C _15624_/A _11521_/X vssd1 vssd1 vccd1 vccd1 _11536_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_62_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15290_ _15290_/A _15290_/B vssd1 vssd1 vccd1 vccd1 _22872_/D sky130_fd_sc_hd__nor2_1
XFILLER_157_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20972__A _20972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ _14155_/B _14237_/X _14239_/Y _14240_/X vssd1 vssd1 vccd1 vccd1 _14253_/A
+ sky130_fd_sc_hd__o211ai_4
X_11453_ _11565_/A _11444_/Y _11452_/X vssd1 vssd1 vccd1 vccd1 _11894_/A sky130_fd_sc_hd__a21o_1
XFILLER_11_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14172_ _14172_/A _14172_/B _14172_/C vssd1 vssd1 vccd1 vccd1 _14285_/A sky130_fd_sc_hd__nand3_1
X_11384_ _11384_/A vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_192_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13586__A _13630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13123_ _13176_/A vssd1 vssd1 vccd1 vccd1 _13577_/A sky130_fd_sc_hd__buf_2
XFILLER_98_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18980_ _18980_/A _19771_/A _18980_/C vssd1 vssd1 vccd1 vccd1 _18980_/X sky130_fd_sc_hd__and3_1
XFILLER_125_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _17833_/X _19896_/B _19842_/D _17930_/X vssd1 vssd1 vccd1 vccd1 _17932_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _22726_/Q vssd1 vssd1 vccd1 vccd1 _13055_/A sky130_fd_sc_hd__buf_2
XFILLER_3_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22909__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12005_ _12018_/A _11511_/A _11425_/Y _18508_/A _12001_/Y vssd1 vssd1 vccd1 vccd1
+ _12006_/B sky130_fd_sc_hd__o221ai_4
XANTENNA__18632__A1 _12204_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17862_ _22902_/Q vssd1 vssd1 vccd1 vccd1 _17862_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16643__B1 _16351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19601_ _19477_/X _19475_/Y _19479_/C vssd1 vssd1 vccd1 vccd1 _19605_/B sky130_fd_sc_hd__o21ai_2
XFILLER_121_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16813_ _16831_/A vssd1 vssd1 vccd1 vccd1 _16828_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17793_ _22901_/Q _17793_/B _17793_/C vssd1 vssd1 vccd1 vccd1 _17794_/B sky130_fd_sc_hd__nor3_1
XFILLER_4_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21519__A1 _21376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19532_ _19532_/A vssd1 vssd1 vccd1 vccd1 _19538_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15306__A _16256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16744_ _16742_/Y _16743_/X _16732_/Y vssd1 vssd1 vccd1 vccd1 _16749_/B sky130_fd_sc_hd__o21ai_1
X_13956_ _13957_/B _13957_/C _13957_/A vssd1 vssd1 vccd1 vccd1 _14034_/A sky130_fd_sc_hd__a21o_1
XFILLER_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19463_ _19318_/Y _19625_/A _19461_/X _19462_/Y vssd1 vssd1 vccd1 vccd1 _19476_/C
+ sky130_fd_sc_hd__o211ai_4
X_12907_ _16129_/C _16078_/B _15804_/C _20355_/D vssd1 vssd1 vccd1 vccd1 _12958_/B
+ sky130_fd_sc_hd__nand4_2
X_16675_ _16675_/A _22893_/Q _16675_/C vssd1 vssd1 vccd1 vccd1 _16675_/Y sky130_fd_sc_hd__nand3_1
X_13887_ _14118_/B _14013_/A _14013_/B _13877_/B _13877_/A vssd1 vssd1 vccd1 vccd1
+ _13887_/X sky130_fd_sc_hd__a32o_1
XFILLER_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18414_ _18308_/Y _18309_/X _18406_/Y _18409_/Y vssd1 vssd1 vccd1 vccd1 _18415_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15626_ _20471_/A vssd1 vssd1 vccd1 vccd1 _16563_/A sky130_fd_sc_hd__clkbuf_2
X_12838_ _12838_/A _12838_/B vssd1 vssd1 vccd1 vccd1 _12855_/A sky130_fd_sc_hd__nand2_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ _19394_/A _19394_/B _19394_/C vssd1 vssd1 vccd1 vccd1 _19407_/A sky130_fd_sc_hd__nand3_1
XFILLER_62_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18345_ _18345_/A _18345_/B _18345_/C vssd1 vssd1 vccd1 vccd1 _18355_/A sky130_fd_sc_hd__nand3_1
X_15557_ _15557_/A _15559_/B _15558_/C _20133_/B vssd1 vssd1 vccd1 vccd1 _15557_/Y
+ sky130_fd_sc_hd__nand4_4
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _12769_/A _12769_/B vssd1 vssd1 vccd1 vccd1 _12769_/Y sky130_fd_sc_hd__nand2_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19360__A2 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14508_ _14699_/B vssd1 vssd1 vccd1 vccd1 _14869_/B sky130_fd_sc_hd__buf_2
XFILLER_174_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15488_ _16217_/A _16218_/A vssd1 vssd1 vccd1 vccd1 _15489_/A sky130_fd_sc_hd__nand2_2
X_18276_ _18276_/A _18276_/B vssd1 vssd1 vccd1 vccd1 _18277_/B sky130_fd_sc_hd__nand2_1
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14185__A1 _13930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17227_ _17227_/A vssd1 vssd1 vccd1 vccd1 _17227_/X sky130_fd_sc_hd__buf_2
Xinput20 wb_adr_i[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
X_14439_ _14439_/A _22967_/Q _16242_/B _14439_/D vssd1 vssd1 vccd1 vccd1 _14440_/A
+ sky130_fd_sc_hd__and4_1
Xinput31 wb_adr_i[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput42 wb_dat_i[16] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__20258__A1 _12671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput53 wb_dat_i[26] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput64 wb_dat_i[7] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_4
X_17158_ _17158_/A _17158_/B vssd1 vssd1 vccd1 vccd1 _17158_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput75 x[4] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1014 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16109_ _12500_/X _12501_/X _16613_/C _16166_/A _16107_/X vssd1 vssd1 vccd1 vccd1
+ _16166_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_6_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17674__A2 _21083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17089_ _17081_/Y _17082_/X _17086_/Y _17088_/X vssd1 vssd1 vccd1 vccd1 _17310_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_115_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12499__B2 _15455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15437__A1 _15482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19614__C _19614_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21218__A _21638_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22810_ _22810_/CLK _22810_/D vssd1 vssd1 vccd1 vccd1 _22810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_700 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12120__B1 _12115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17729__A3 _11666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22741_ _22742_/CLK _22741_/D vssd1 vssd1 vccd1 vccd1 _22741_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__20194__B1 _12754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20733__A2 _16129_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19337__A2_N _19512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17431__A _19615_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22672_ _22943_/CLK _22672_/D vssd1 vssd1 vccd1 vccd1 _22672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18246__B _18246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21623_ _21620_/X _21622_/X _21645_/A _21763_/A vssd1 vssd1 vccd1 vccd1 _21624_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_34_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12423__A1 _15326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12974__A2 _16067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21554_ _21560_/A _21576_/A _21695_/A _21556_/A vssd1 vssd1 vccd1 vccd1 _21566_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_166_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12294__B _12294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20505_ _15631_/X _12378_/B _20611_/B _16450_/B _15911_/A vssd1 vssd1 vccd1 vccd1
+ _20505_/Y sky130_fd_sc_hd__o2111ai_4
XANTENNA_clkbuf_3_5_0_bq_clk_i_A clkbuf_3_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19358__A _19358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16597__A1_N _16599_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21485_ _21485_/A vssd1 vssd1 vccd1 vccd1 _21485_/X sky130_fd_sc_hd__buf_2
XFILLER_107_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20436_ _20553_/A _20553_/B _20309_/A vssd1 vssd1 vccd1 vccd1 _20437_/A sky130_fd_sc_hd__a21o_1
XFILLER_146_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20367_ _20363_/Y _20365_/Y _20366_/Y vssd1 vssd1 vccd1 vccd1 _20367_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_161_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22106_ _22106_/A vssd1 vssd1 vccd1 vccd1 _22221_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_161_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20298_ _20298_/A _20298_/B _20319_/B vssd1 vssd1 vccd1 vccd1 _20300_/B sky130_fd_sc_hd__nand3_1
XFILLER_103_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22037_ _22037_/A _22037_/B _22037_/C _22182_/B vssd1 vssd1 vccd1 vccd1 _22037_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_88_652 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_847 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20032__A _22926_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13810_ _13810_/A _13810_/B _13810_/C vssd1 vssd1 vccd1 vccd1 _13826_/A sky130_fd_sc_hd__nand3_4
XFILLER_21_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14790_ _14366_/X _14863_/B _14869_/B _14775_/D vssd1 vssd1 vccd1 vccd1 _14792_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__13572__C _21866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1038 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22174__A1 _22231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13741_ _13963_/D vssd1 vssd1 vccd1 vccd1 _13833_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22939_ _22943_/CLK _22939_/D vssd1 vssd1 vccd1 vccd1 _22939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17341__A _17341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16460_ _11935_/B _15341_/X _16451_/A vssd1 vssd1 vccd1 vccd1 _16463_/B sky130_fd_sc_hd__o21ai_1
X_13672_ _13672_/A _13672_/B _13672_/C vssd1 vssd1 vccd1 vccd1 _13672_/Y sky130_fd_sc_hd__nand3_1
X_15411_ _15411_/A vssd1 vssd1 vccd1 vccd1 _15703_/B sky130_fd_sc_hd__buf_2
X_12623_ _12455_/Y _12620_/Y _12621_/Y _12622_/Y vssd1 vssd1 vccd1 vccd1 _12624_/A
+ sky130_fd_sc_hd__o211ai_2
X_16391_ _16391_/A _16391_/B _16391_/C vssd1 vssd1 vccd1 vccd1 _16393_/B sky130_fd_sc_hd__nand3_1
XFILLER_31_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12485__A _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20488__A1 _12721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15342_ _15891_/A _15341_/X _15336_/Y vssd1 vssd1 vccd1 vccd1 _15342_/Y sky130_fd_sc_hd__o21ai_1
X_18130_ _18133_/A _19587_/D _18130_/C vssd1 vssd1 vccd1 vccd1 _18130_/Y sky130_fd_sc_hd__nand3b_1
X_12554_ _12771_/A _12773_/A _12515_/A _20128_/A _12970_/A vssd1 vssd1 vccd1 vccd1
+ _12557_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_106_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16156__A2 _20429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11505_ _11505_/A vssd1 vssd1 vccd1 vccd1 _11505_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18061_ _18061_/A _18061_/B vssd1 vssd1 vccd1 vccd1 _18061_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15273_ _15273_/A _15273_/B vssd1 vssd1 vccd1 vccd1 _22866_/D sky130_fd_sc_hd__nand2_1
XFILLER_145_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ _17141_/A vssd1 vssd1 vccd1 vccd1 _16515_/A sky130_fd_sc_hd__buf_2
XFILLER_156_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17012_ _16732_/A _16732_/B _16723_/X _16743_/X vssd1 vssd1 vccd1 vccd1 _17025_/C
+ sky130_fd_sc_hd__a31o_2
X_14224_ _14506_/B vssd1 vssd1 vccd1 vccd1 _15006_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12717__A2 _15326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11436_ _11436_/A _11713_/B vssd1 vssd1 vccd1 vccd1 _11448_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14155_ _14238_/B _14155_/B vssd1 vssd1 vccd1 vccd1 _14163_/A sky130_fd_sc_hd__nand2_1
X_11367_ _12018_/A vssd1 vssd1 vccd1 vccd1 _18795_/A sky130_fd_sc_hd__buf_2
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13106_ _21315_/B vssd1 vssd1 vccd1 vccd1 _21750_/C sky130_fd_sc_hd__buf_2
XFILLER_140_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18963_ _19293_/A _19294_/A _18783_/A _18958_/A vssd1 vssd1 vccd1 vccd1 _18964_/D
+ sky130_fd_sc_hd__o211ai_1
X_14086_ _14510_/A _14126_/B _14868_/C _14191_/A _14270_/A vssd1 vssd1 vccd1 vccd1
+ _14086_/X sky130_fd_sc_hd__a32o_1
XFILLER_98_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _22786_/Q vssd1 vssd1 vccd1 vccd1 _11420_/B sky130_fd_sc_hd__inv_2
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17914_ _17914_/A _17960_/A vssd1 vssd1 vccd1 vccd1 _17915_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18605__A1 _18432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _13037_/A _13037_/B vssd1 vssd1 vccd1 vccd1 _13038_/D sky130_fd_sc_hd__nand2_1
XFILLER_152_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15962__C _17643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18894_ _18901_/A _18897_/A _18891_/X _18893_/X vssd1 vssd1 vccd1 vccd1 _18899_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_65_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22881__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17845_ _17869_/A _17845_/B vssd1 vssd1 vccd1 vccd1 _17860_/B sky130_fd_sc_hd__xnor2_4
XFILLER_113_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17235__B _19351_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19015__D1 _19490_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17776_ _17776_/A vssd1 vssd1 vccd1 vccd1 _17954_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14988_ _15046_/A _14987_/C _15046_/B vssd1 vssd1 vccd1 vccd1 _14989_/B sky130_fd_sc_hd__a21oi_1
X_19515_ _19511_/B _19580_/A _19511_/A vssd1 vssd1 vccd1 vccd1 _19521_/C sky130_fd_sc_hd__a21o_1
X_16727_ _11295_/A _11295_/B _16582_/A _16584_/A vssd1 vssd1 vccd1 vccd1 _16727_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13939_ _14465_/B vssd1 vssd1 vccd1 vccd1 _14771_/A sky130_fd_sc_hd__buf_2
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13850__B1 _13896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17041__B1 _17040_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17251__A _17251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19446_ _19446_/A _19561_/B vssd1 vssd1 vccd1 vccd1 _19681_/B sky130_fd_sc_hd__nand2_2
X_16658_ _16206_/X _15879_/A _16406_/A _16433_/Y vssd1 vssd1 vccd1 vccd1 _16659_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15609_ _20461_/B vssd1 vssd1 vccd1 vccd1 _20463_/B sky130_fd_sc_hd__buf_2
X_19377_ _19179_/A _19179_/B _19179_/C _19182_/C vssd1 vssd1 vccd1 vccd1 _19377_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_72_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16589_ _16595_/B _16588_/Y _16595_/A vssd1 vssd1 vccd1 vccd1 _16594_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12395__A _12467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17401__D _17401_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18136__A3 _19464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18328_ _18328_/A _18328_/B _18328_/C vssd1 vssd1 vccd1 vccd1 _18529_/B sky130_fd_sc_hd__and3_1
XFILLER_188_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18541__B1 _18534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18259_ _18259_/A _18259_/B vssd1 vssd1 vccd1 vccd1 _18590_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12169__B1 _12164_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21270_ _21270_/A _21841_/A _21270_/C _21299_/B vssd1 vssd1 vccd1 vccd1 _21270_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_118_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20221_ _20355_/A _20477_/A _20456_/C _20463_/C vssd1 vssd1 vccd1 vccd1 _20221_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_190_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18844__A1 _19470_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20100__B1 _12988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18810__A _18810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17129__C _20323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__A1 _11502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14115__A _14165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15658__A1 _15616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20152_ _20143_/A _20143_/B _20125_/A _20155_/A vssd1 vssd1 vccd1 vccd1 _20197_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17426__A _17426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ _20219_/B vssd1 vssd1 vccd1 vccd1 _20083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16083__A1 _11561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11474__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20985_ _20985_/A _20985_/B _20985_/C vssd1 vssd1 vccd1 vccd1 _20985_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__20706__A2 _17424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22724_ _22725_/CLK _22724_/D vssd1 vssd1 vccd1 vccd1 _22724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18780__B1 _18779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22655_ _22655_/A vssd1 vssd1 vccd1 vccd1 _22814_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16791__C1 _19358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19324__A2 _19464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21606_ _21606_/A vssd1 vssd1 vccd1 vccd1 _21606_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22586_ _22514_/A _22586_/B _22586_/C _22586_/D vssd1 vssd1 vccd1 vccd1 _22643_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_159_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_903 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21537_ _21537_/A vssd1 vssd1 vccd1 vccd1 _21537_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15897__A1 _15891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12270_ _22703_/Q vssd1 vssd1 vccd1 vccd1 _12369_/A sky130_fd_sc_hd__clkbuf_2
X_21468_ _22730_/Q _22731_/Q _22732_/Q vssd1 vssd1 vccd1 vccd1 _21583_/C sky130_fd_sc_hd__nor3_1
XFILLER_182_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11907__B1 _18953_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17638__A2 _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20419_ _20281_/A _20281_/B _20429_/C vssd1 vssd1 vccd1 vccd1 _20420_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__19493__D1 _19351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17039__C _17039_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21399_ _21399_/A _21399_/B _21399_/C _22851_/Q vssd1 vssd1 vccd1 vccd1 _21547_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_4_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_991 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12580__B1 _17532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1075 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17981__D _17981_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15960_ _15960_/A vssd1 vssd1 vccd1 vccd1 _17645_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_89_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_A wb_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14911_ _14911_/A _14963_/C _14911_/C vssd1 vssd1 vccd1 vccd1 _14912_/B sky130_fd_sc_hd__and3_1
X_15891_ _15891_/A vssd1 vssd1 vccd1 vccd1 _16098_/A sky130_fd_sc_hd__buf_4
XANTENNA__11686__A2 _11673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16074__A1 _12294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17630_ _19772_/C vssd1 vssd1 vccd1 vccd1 _19844_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_124_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17810__A2 _20972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14842_ _14842_/A _14842_/B vssd1 vssd1 vccd1 vccd1 _14845_/A sky130_fd_sc_hd__xnor2_4
XFILLER_76_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20697__A _20697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17561_ _16579_/X _16580_/X _19013_/C _21011_/A vssd1 vssd1 vccd1 vccd1 _17564_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_90_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11985_ _12137_/B _11981_/X _11982_/Y _11984_/Y vssd1 vssd1 vccd1 vccd1 _11986_/A
+ sky130_fd_sc_hd__o211ai_1
X_14773_ _14362_/X _13973_/B _13907_/X _13970_/X _14593_/B vssd1 vssd1 vccd1 vccd1
+ _14791_/A sky130_fd_sc_hd__o41ai_4
X_19300_ _19131_/B _19131_/A _19147_/X _19299_/Y _19274_/Y vssd1 vssd1 vccd1 vccd1
+ _19301_/C sky130_fd_sc_hd__o2111ai_1
X_16512_ _16512_/A _16512_/B vssd1 vssd1 vccd1 vccd1 _16512_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13724_ _22753_/Q vssd1 vssd1 vccd1 vccd1 _13810_/B sky130_fd_sc_hd__clkinv_2
XFILLER_56_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17492_ _17514_/A _17493_/A _17494_/A vssd1 vssd1 vccd1 vccd1 _17497_/A sky130_fd_sc_hd__a21o_1
XFILLER_140_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19231_ _19231_/A _19231_/B _19231_/C vssd1 vssd1 vccd1 vccd1 _19231_/X sky130_fd_sc_hd__and3_1
X_16443_ _16422_/A _16204_/Y _16442_/Y vssd1 vssd1 vccd1 vccd1 _17078_/A sky130_fd_sc_hd__a21oi_2
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13655_ _13658_/C _13655_/B _13655_/C vssd1 vssd1 vccd1 vccd1 _13660_/A sky130_fd_sc_hd__nand3b_1
XFILLER_158_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19162_ _15936_/A _19517_/A _19792_/A _16554_/C _19156_/B vssd1 vssd1 vccd1 vccd1
+ _19162_/Y sky130_fd_sc_hd__o2111ai_4
X_12606_ _12606_/A vssd1 vssd1 vccd1 vccd1 _12606_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16374_ _15510_/B _15672_/Y _16373_/Y vssd1 vssd1 vccd1 vccd1 _16374_/Y sky130_fd_sc_hd__o21ai_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13586_ _13630_/A _21805_/B _13664_/A _21878_/C vssd1 vssd1 vccd1 vccd1 _13586_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18113_ _18279_/A _18278_/A _18184_/B vssd1 vssd1 vccd1 vccd1 _18113_/Y sky130_fd_sc_hd__a21oi_1
X_15325_ _15325_/A vssd1 vssd1 vccd1 vccd1 _15325_/X sky130_fd_sc_hd__buf_4
X_12537_ _22823_/Q vssd1 vssd1 vccd1 vccd1 _12547_/A sky130_fd_sc_hd__inv_2
XFILLER_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17877__A2 _21048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19093_ _18908_/C _19091_/X _18871_/Y _19092_/Y vssd1 vssd1 vccd1 vccd1 _19095_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_76_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14861__C _14861_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18044_ _18044_/A vssd1 vssd1 vccd1 vccd1 _18082_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15256_ _15242_/A _15241_/A _15241_/B _15243_/B _15243_/A vssd1 vssd1 vccd1 vccd1
+ _15266_/B sky130_fd_sc_hd__a32oi_4
XFILLER_32_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ _20210_/A _12988_/C vssd1 vssd1 vccd1 vccd1 _12469_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14207_ _14203_/X _14185_/X _14206_/Y vssd1 vssd1 vccd1 vccd1 _14207_/Y sky130_fd_sc_hd__o21ai_1
X_11419_ _11378_/X _12148_/B _11420_/D _11394_/A _11430_/C vssd1 vssd1 vccd1 vccd1
+ _12170_/A sky130_fd_sc_hd__a311oi_4
X_15187_ _15186_/B _15186_/C _15182_/A _14942_/B vssd1 vssd1 vccd1 vccd1 _15187_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_12399_ _12598_/A vssd1 vssd1 vccd1 vccd1 _12844_/A sky130_fd_sc_hd__buf_2
XANTENNA__18630__A _19507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16837__B1 _16836_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ _14134_/Y _14135_/X _14491_/C _14111_/X _14191_/B vssd1 vssd1 vccd1 vccd1
+ _14154_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_154_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19995_ _19995_/A _19995_/B vssd1 vssd1 vccd1 vccd1 _19998_/B sky130_fd_sc_hd__xor2_1
XFILLER_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17246__A _17246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18946_ _18953_/A _20012_/A _18953_/C _18627_/Y vssd1 vssd1 vccd1 vccd1 _18946_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_101_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14069_ _14069_/A _14200_/A _14069_/C vssd1 vssd1 vccd1 vccd1 _14085_/A sky130_fd_sc_hd__nand3_4
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18877_ _18877_/A _18983_/A vssd1 vssd1 vccd1 vccd1 _18881_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17828_ _17890_/A _17827_/C _17827_/A vssd1 vssd1 vccd1 vccd1 _17831_/C sky130_fd_sc_hd__a21o_1
XANTENNA__19461__A _19461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14076__B1 _14721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17759_ _17760_/B _17760_/C _17760_/A vssd1 vssd1 vccd1 vccd1 _17761_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11444__D _15912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13823__B1 _13799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17014__B1 _17006_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21215__B _21609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20770_ _20770_/A vssd1 vssd1 vccd1 vccd1 _20772_/A sky130_fd_sc_hd__inv_2
XFILLER_74_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17565__A1 _17427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12837__B _20130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19429_ _19271_/Y _19268_/Y _19130_/B _19147_/X _19274_/Y vssd1 vssd1 vccd1 vccd1
+ _19429_/Y sky130_fd_sc_hd__o2111ai_2
XFILLER_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19306__A2 _11351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_566 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22440_ _22440_/A vssd1 vssd1 vccd1 vccd1 _22719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18514__B1 _15893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22371_ _22439_/S vssd1 vssd1 vccd1 vccd1 _22380_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__13949__A _13949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16325__A _16325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21322_ _21197_/Y _21591_/B _21615_/A _21202_/Y vssd1 vssd1 vccd1 vccd1 _21332_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__20872__A1 _17816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19636__A _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21253_ _21251_/X _21299_/A vssd1 vssd1 vccd1 vccd1 _21260_/B sky130_fd_sc_hd__and2b_1
XFILLER_150_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11365__A1 _18116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20204_ _20084_/Y _20085_/X _20088_/X _20093_/Y vssd1 vssd1 vccd1 vccd1 _20204_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18293__A2 _19043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21184_ _13050_/X _21183_/X _13316_/X _13317_/X vssd1 vssd1 vccd1 vccd1 _21184_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22062__A _22062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20135_ _12786_/Y _20133_/Y _20134_/X _20131_/Y vssd1 vssd1 vccd1 vccd1 _20142_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_942 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20066_ _13041_/Y _20064_/Y _20065_/Y _22929_/Q vssd1 vssd1 vccd1 vccd1 _20192_/A
+ sky130_fd_sc_hd__a211oi_4
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11783_/A vssd1 vssd1 vccd1 vccd1 _11770_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ _20844_/A _17928_/D _20923_/B _20936_/D vssd1 vssd1 vccd1 vccd1 _20969_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22707_ _22802_/CLK _22707_/D vssd1 vssd1 vccd1 vccd1 _22707_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20899_ _20961_/A _20961_/B _22937_/Q vssd1 vssd1 vccd1 vccd1 _20901_/A sky130_fd_sc_hd__a21oi_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ _13440_/A _13440_/B vssd1 vssd1 vccd1 vccd1 _13546_/B sky130_fd_sc_hd__nand2_1
XFILLER_139_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22638_ _22638_/A vssd1 vssd1 vccd1 vccd1 _22806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16880__D _17039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14790__A1 _14366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13371_ _13257_/B _13234_/A _13234_/B _21584_/C _13202_/Y vssd1 vssd1 vccd1 vccd1
+ _13373_/A sky130_fd_sc_hd__o311ai_4
XANTENNA__13859__A _22858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22569_ _22776_/Q input51/X _22569_/S vssd1 vssd1 vccd1 vccd1 _22570_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21498__D _21498_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15110_ _15108_/Y _15074_/C _15149_/A _15152_/A vssd1 vssd1 vccd1 vccd1 _15111_/B
+ sky130_fd_sc_hd__o211a_1
X_12322_ _16267_/A _16266_/A _12596_/A _16268_/A vssd1 vssd1 vccd1 vccd1 _12322_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16090_ _16090_/A _16090_/B vssd1 vssd1 vccd1 vccd1 _16090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input79_A x[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15041_ _15046_/A _15046_/B vssd1 vssd1 vccd1 vccd1 _15175_/C sky130_fd_sc_hd__nor2_1
XFILLER_119_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12253_ _18272_/A _18272_/C vssd1 vssd1 vccd1 vccd1 _18241_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21812__B1 _21806_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18284__A2 _17388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12184_ _12184_/A vssd1 vssd1 vccd1 vccd1 _12184_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18800_ _15530_/X _15531_/X _11598_/X vssd1 vssd1 vccd1 vccd1 _19052_/A sky130_fd_sc_hd__a21oi_2
X_19780_ _19848_/B _19783_/B vssd1 vssd1 vccd1 vccd1 _19781_/A sky130_fd_sc_hd__nand2_1
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16992_ _11504_/X _11505_/X _11779_/B _16563_/B _16563_/A vssd1 vssd1 vccd1 vccd1
+ _16998_/A sky130_fd_sc_hd__o2111ai_2
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ _18741_/C _18741_/D _18725_/A vssd1 vssd1 vccd1 vccd1 _18731_/X sky130_fd_sc_hd__a21o_1
XFILLER_122_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15943_ _15784_/Y _15803_/Y _15828_/X _15826_/Y vssd1 vssd1 vccd1 vccd1 _15944_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20918__A2 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18662_ _18662_/A vssd1 vssd1 vccd1 vccd1 _18827_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15874_ _15883_/A _15874_/B vssd1 vssd1 vccd1 vccd1 _15875_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12003__A _12003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14058__B1 _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18992__B1 _18986_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17613_ _17611_/X _17713_/A _17612_/Y vssd1 vssd1 vccd1 vccd1 _17722_/A sky130_fd_sc_hd__o21ai_1
XFILLER_97_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14825_ _14825_/A _14902_/B _14825_/C vssd1 vssd1 vccd1 vccd1 _14826_/C sky130_fd_sc_hd__nand3_1
XANTENNA__12608__A1 _12606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18593_ _19293_/A _19294_/A _18430_/A _18592_/Y _18960_/C vssd1 vssd1 vccd1 vccd1
+ _18595_/B sky130_fd_sc_hd__o221ai_2
XANTENNA__21328__C1 _14380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12938__A _12938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _17536_/X _17544_/B _17544_/C vssd1 vssd1 vccd1 vccd1 _17544_/Y sky130_fd_sc_hd__nand3b_2
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14756_ _14756_/A _14756_/B _14756_/C vssd1 vssd1 vccd1 vccd1 _14757_/B sky130_fd_sc_hd__nand3_1
X_11968_ _11974_/A _11968_/B _11974_/C vssd1 vssd1 vccd1 vccd1 _12126_/A sky130_fd_sc_hd__nand3_1
XANTENNA__16129__B _20390_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11292__B1 _22968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ _13707_/A _13707_/B _13845_/B vssd1 vssd1 vccd1 vccd1 _14258_/D sky130_fd_sc_hd__and3_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17475_ _17475_/A _17475_/B _17475_/C vssd1 vssd1 vccd1 vccd1 _17475_/X sky130_fd_sc_hd__and3_1
XANTENNA__16755__C1 _16853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14687_ _14998_/A _14467_/X _14793_/A _14685_/Y _14686_/X vssd1 vssd1 vccd1 vccd1
+ _14687_/X sky130_fd_sc_hd__o311a_1
X_11899_ _11899_/A _11899_/B _11902_/B _11902_/C vssd1 vssd1 vccd1 vccd1 _11900_/B
+ sky130_fd_sc_hd__nand4_1
X_19214_ _19062_/B _19055_/Y _19051_/X _19059_/Y vssd1 vssd1 vccd1 vccd1 _19227_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16426_ _16664_/A vssd1 vssd1 vccd1 vccd1 _16426_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13638_ _21866_/C vssd1 vssd1 vccd1 vccd1 _22062_/A sky130_fd_sc_hd__buf_2
XFILLER_158_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20593__C _20593_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19145_ _19145_/A _19145_/B vssd1 vssd1 vccd1 vccd1 _22895_/D sky130_fd_sc_hd__xor2_1
XFILLER_192_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16357_ _20854_/A vssd1 vssd1 vccd1 vccd1 _17833_/B sky130_fd_sc_hd__buf_2
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13569_ _21621_/C vssd1 vssd1 vccd1 vccd1 _21944_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11595__A1 _15904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15308_ _15308_/A vssd1 vssd1 vccd1 vccd1 _15309_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19076_ _19104_/A _19096_/A vssd1 vssd1 vccd1 vccd1 _19098_/C sky130_fd_sc_hd__nand2_1
XFILLER_157_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16288_ _16288_/A _16540_/A _16288_/C vssd1 vssd1 vccd1 vccd1 _16288_/Y sky130_fd_sc_hd__nand3_1
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18027_ _19418_/C vssd1 vssd1 vccd1 vccd1 _20012_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11289__A _22968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15239_ _15240_/D _15240_/B _14990_/X _15217_/B vssd1 vssd1 vccd1 vccd1 _15241_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14533__B2 _14273_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13887__A3 _14013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11898__A2 _11899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19978_ _19975_/Y _19974_/B _19976_/Y _19977_/X vssd1 vssd1 vccd1 vccd1 _19978_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_119_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17407__C _18303_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18929_ _18929_/A _18929_/B vssd1 vssd1 vccd1 vccd1 _18977_/B sky130_fd_sc_hd__nand2_2
XFILLER_80_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22610__A _22656_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21940_ _21940_/A vssd1 vssd1 vccd1 vccd1 _22045_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21871_ _21871_/A vssd1 vssd1 vccd1 vccd1 _21939_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__20790__B1 _20793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20130__A _20130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15261__A2 _15247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14766__C _14911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20822_ _20822_/A _20822_/B _20822_/C vssd1 vssd1 vccd1 vccd1 _20890_/C sky130_fd_sc_hd__nand3_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1030 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20753_ _20539_/Y _20543_/Y _20652_/Y _20660_/A _20546_/Y vssd1 vssd1 vccd1 vccd1
+ _20754_/C sky130_fd_sc_hd__o2111a_1
XANTENNA__11822__A2 _11736_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20684_ _20717_/B _20686_/A vssd1 vssd1 vccd1 vccd1 _20718_/A sky130_fd_sc_hd__nor2_1
XANTENNA__16761__A2 _16227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22423_ _22423_/A vssd1 vssd1 vccd1 vccd1 _22711_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12232__C1 _11721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12583__A _12583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12783__B1 _20502_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__B2 _18156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22354_ _22354_/A _22354_/B _22687_/Q vssd1 vssd1 vccd1 vccd1 _22355_/A sky130_fd_sc_hd__nor3b_1
XFILLER_40_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21305_ _21307_/A _21307_/C _21307_/B vssd1 vssd1 vccd1 vccd1 _21312_/A sky130_fd_sc_hd__a21o_1
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22285_ _22285_/A _22285_/B vssd1 vssd1 vccd1 vccd1 _22286_/A sky130_fd_sc_hd__or2_1
XFILLER_191_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21236_ _21234_/X _21235_/Y _13315_/X vssd1 vssd1 vccd1 vccd1 _21239_/B sky130_fd_sc_hd__o21ai_1
XFILLER_116_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16277__A1 _16179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16277__B2 _16177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21167_ _21167_/A _21167_/B vssd1 vssd1 vccd1 vccd1 _22928_/D sky130_fd_sc_hd__nand2_2
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13845__C _13896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_78 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20118_ _20118_/A _20118_/B vssd1 vssd1 vccd1 vccd1 _20121_/A sky130_fd_sc_hd__nand2_1
XFILLER_77_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22942__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21098_ _21097_/Y _21068_/A _21094_/Y vssd1 vssd1 vccd1 vccd1 _21115_/A sky130_fd_sc_hd__o21bai_1
XFILLER_105_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19766__A2 _19842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20049_ _20049_/A _20049_/B _20049_/C vssd1 vssd1 vccd1 vccd1 _20051_/A sky130_fd_sc_hd__and3_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12940_ _20463_/C vssd1 vssd1 vccd1 vccd1 _13016_/C sky130_fd_sc_hd__buf_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_934 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20678__C _20917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12871_ _12862_/A _12857_/A _12864_/B vssd1 vssd1 vccd1 vccd1 _12872_/C sky130_fd_sc_hd__a21o_1
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12758__A _12758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19518__A2 _18980_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11662__A _18648_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14610_ _14600_/Y _14602_/Y _14712_/A _14712_/B vssd1 vssd1 vccd1 vccd1 _14611_/D
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _18778_/A _11736_/Y _11821_/X _11762_/B _11932_/A vssd1 vssd1 vccd1 vccd1
+ _11822_/X sky130_fd_sc_hd__o311a_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _16940_/A _12727_/A _15439_/A _15524_/X vssd1 vssd1 vccd1 vccd1 _16265_/B
+ sky130_fd_sc_hd__o22ai_4
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _16447_/A vssd1 vssd1 vccd1 vccd1 _17280_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _14524_/Y _14541_/B _14541_/C _14541_/D vssd1 vssd1 vccd1 vccd1 _14544_/A
+ sky130_fd_sc_hd__nand4b_2
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11813__A2 _11809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18445__A _18445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20694__B _20793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_847 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17260_/A _17260_/B _17260_/C vssd1 vssd1 vccd1 vccd1 _17268_/B sky130_fd_sc_hd__nand3_1
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ _12117_/A vssd1 vssd1 vccd1 vccd1 _16276_/A sky130_fd_sc_hd__clkbuf_2
X_14472_ _14472_/A _14472_/B _14472_/C vssd1 vssd1 vccd1 vccd1 _14500_/A sky130_fd_sc_hd__nand3_2
XFILLER_42_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16752__A2 _16598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16211_ _16206_/X _15879_/X _16210_/Y vssd1 vssd1 vccd1 vccd1 _16211_/Y sky130_fd_sc_hd__o21ai_1
X_13423_ _13423_/A _21259_/B _13487_/A _21259_/C vssd1 vssd1 vccd1 vccd1 _13424_/A
+ sky130_fd_sc_hd__or4_1
X_17191_ _17019_/A _17019_/B _17190_/Y _16989_/C vssd1 vssd1 vccd1 vccd1 _17191_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_139_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12493__A _12493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16142_ _16132_/Y _16137_/Y _16140_/Y _16141_/X vssd1 vssd1 vccd1 vccd1 _16145_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_13354_ _13354_/A _13354_/B vssd1 vssd1 vccd1 vccd1 _13354_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15300__C _15901_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12305_ _22820_/Q vssd1 vssd1 vccd1 vccd1 _12348_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16073_ _16050_/Y _16051_/X _16047_/A _16047_/B vssd1 vssd1 vccd1 vccd1 _16073_/Y
+ sky130_fd_sc_hd__o211ai_4
X_13285_ _13475_/C _13475_/A _13475_/B vssd1 vssd1 vccd1 vccd1 _13288_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__22589__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_596 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19901_ _19901_/A _19901_/B _19901_/C _19901_/D vssd1 vssd1 vccd1 vccd1 _19901_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_154_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _15445_/B vssd1 vssd1 vccd1 vccd1 _15531_/A sky130_fd_sc_hd__buf_2
X_15024_ _15213_/A _14562_/X _15023_/B vssd1 vssd1 vccd1 vccd1 _15024_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_142_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17508__B _22898_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19832_ _19832_/A vssd1 vssd1 vccd1 vccd1 _22901_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15309__A _15309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ _18855_/A vssd1 vssd1 vccd1 vccd1 _12167_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19763_ _19764_/C _19746_/Y _19747_/A vssd1 vssd1 vccd1 vccd1 _19763_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__19206__A1 _19211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16975_ _16941_/X _16944_/Y _16934_/A vssd1 vssd1 vccd1 vccd1 _16976_/A sky130_fd_sc_hd__o21ai_1
XFILLER_111_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12098_ _11366_/A _11819_/A _12097_/Y vssd1 vssd1 vccd1 vccd1 _12098_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_65_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15491__A2 _12211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18714_ _18491_/A _18518_/A _18916_/B vssd1 vssd1 vccd1 vccd1 _18723_/A sky130_fd_sc_hd__a21oi_1
X_15926_ _15793_/Y _15794_/X _15915_/A _15915_/B vssd1 vssd1 vccd1 vccd1 _15967_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_65_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19694_ _19694_/A _19694_/B _19771_/A _19694_/D vssd1 vssd1 vccd1 vccd1 _19697_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11501__A1 _11381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 wb_adr_i[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21564__A2 _21285_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18645_ _18646_/A _18646_/B _18646_/C vssd1 vssd1 vccd1 vccd1 _18645_/Y sky130_fd_sc_hd__a21oi_2
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _15883_/A _15874_/B _15856_/Y vssd1 vssd1 vccd1 vccd1 _15952_/A sky130_fd_sc_hd__a21oi_2
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11572__A _18303_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14808_ _14808_/A _14808_/B _14808_/C _14808_/D vssd1 vssd1 vccd1 vccd1 _14808_/Y
+ sky130_fd_sc_hd__nand4_1
X_18576_ _18409_/Y _18443_/Y _18406_/Y _18277_/B _18277_/A vssd1 vssd1 vccd1 vccd1
+ _18576_/Y sky130_fd_sc_hd__a32oi_4
XANTENNA__14451__B1 _14448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _15788_/A vssd1 vssd1 vccd1 vccd1 _15921_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16991__A2 _16822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15794__A3 _15792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12387__B _12387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17527_ _15940_/A _17526_/X _17443_/A _17636_/A vssd1 vssd1 vccd1 vccd1 _17531_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14739_ _14733_/A _14733_/B _14737_/A _14737_/B vssd1 vssd1 vccd1 vccd1 _14740_/D
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16728__C1 _16727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17458_ _17458_/A _17458_/B _17458_/C vssd1 vssd1 vccd1 vccd1 _17479_/B sky130_fd_sc_hd__nand3_2
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16409_ _16418_/A _16418_/B _16038_/B _15964_/Y vssd1 vssd1 vccd1 vccd1 _16421_/D
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_20_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17389_ _15941_/A _17388_/X _17235_/Y _17386_/X _17383_/Y vssd1 vssd1 vccd1 vccd1
+ _17550_/B sky130_fd_sc_hd__o311a_1
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19128_ _19113_/X _18812_/Y _18830_/B _19121_/B _19122_/Y vssd1 vssd1 vccd1 vccd1
+ _19129_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_195_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19693__A1 _12207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17153__C1 _16937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19059_ _17381_/A _17380_/A _18665_/A _19351_/B vssd1 vssd1 vccd1 vccd1 _19059_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_195_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22070_ _22075_/A _22075_/B _22079_/B _22079_/C vssd1 vssd1 vccd1 vccd1 _22163_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_195_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20125__A _20125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16322__B _16322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19336__D _19771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21252__A1 _21399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21021_ _21021_/A _21021_/B vssd1 vssd1 vccd1 vccd1 _21023_/A sky130_fd_sc_hd__xor2_1
XFILLER_113_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17434__A _17434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_614 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21923_ _21700_/X _21701_/X _21931_/B vssd1 vssd1 vccd1 vccd1 _21924_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12578__A _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21854_ _21338_/A _21338_/B _21853_/X vssd1 vssd1 vccd1 vccd1 _21854_/X sky130_fd_sc_hd__a21o_2
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20805_ _20717_/B _20717_/A _20683_/B vssd1 vssd1 vccd1 vccd1 _20806_/A sky130_fd_sc_hd__o21ai_1
X_21785_ _21784_/X _21624_/B _21624_/A _21779_/X vssd1 vssd1 vccd1 vccd1 _21785_/Y
+ sky130_fd_sc_hd__a31oi_2
X_20736_ _20631_/B _20631_/C _20631_/A _20735_/Y vssd1 vssd1 vccd1 vccd1 _20737_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17392__C1 _17532_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15401__B _20502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20667_ _22933_/Q _20566_/A _20566_/B _20563_/B _20563_/A vssd1 vssd1 vccd1 vccd1
+ _20667_/Y sky130_fd_sc_hd__o311ai_4
XFILLER_104_1120 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13202__A _13202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22406_ _22406_/A vssd1 vssd1 vccd1 vccd1 _22703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20598_ _20697_/A _17111_/A _20587_/B _20581_/A _20495_/B vssd1 vssd1 vccd1 vccd1
+ _20598_/X sky130_fd_sc_hd__o311a_1
XFILLER_167_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22337_ _22341_/C _22341_/A _22341_/B vssd1 vssd1 vccd1 vccd1 _22338_/B sky130_fd_sc_hd__a21o_1
XFILLER_124_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16513__A _16513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ _13073_/A _13243_/A _13301_/A vssd1 vssd1 vccd1 vccd1 _21213_/A sky130_fd_sc_hd__a21o_1
X_22268_ _22308_/A _22308_/B _22308_/C vssd1 vssd1 vccd1 vccd1 _22272_/C sky130_fd_sc_hd__o21ai_1
XFILLER_3_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16232__B _16771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15774__D _15774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12021_ _12017_/X _12019_/X _12020_/Y vssd1 vssd1 vccd1 vccd1 _12025_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11657__A _15539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21219_ _21237_/B _21944_/A _21219_/C vssd1 vssd1 vccd1 vccd1 _21219_/X sky130_fd_sc_hd__and3_1
X_22199_ _22162_/Y _22166_/Y _22198_/Y vssd1 vssd1 vccd1 vccd1 _22202_/A sky130_fd_sc_hd__a21oi_1
XFILLER_116_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20689__B _20793_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16760_ _16956_/A vssd1 vssd1 vccd1 vccd1 _16760_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13972_ _14583_/B vssd1 vssd1 vccd1 vccd1 _13973_/B sky130_fd_sc_hd__buf_2
XFILLER_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14681__B1 _14998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15711_ _15711_/A vssd1 vssd1 vccd1 vccd1 _16554_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_19_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12923_ _13022_/C _12922_/X _12592_/A _12592_/B _12588_/Y vssd1 vssd1 vccd1 vccd1
+ _12926_/A sky130_fd_sc_hd__o221ai_1
X_16691_ _16669_/A _16670_/A _16695_/C _16695_/D vssd1 vssd1 vccd1 vccd1 _16691_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_46_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18430_ _18430_/A _18601_/A _18601_/B _18600_/A vssd1 vssd1 vccd1 vccd1 _18432_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_34_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15642_ _15336_/Y _16720_/C _16809_/B _15343_/X vssd1 vssd1 vccd1 vccd1 _15642_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_34_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12854_ _12432_/A _12432_/B _12358_/X vssd1 vssd1 vccd1 vccd1 _12856_/B sky130_fd_sc_hd__a21oi_1
XFILLER_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22396__S _22402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _18367_/A _18367_/B _18360_/X vssd1 vssd1 vccd1 vccd1 _18471_/B sky130_fd_sc_hd__a21o_1
XANTENNA__15799__A _15799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11805_ _12024_/A _11810_/C vssd1 vssd1 vccd1 vccd1 _11814_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12638__D _16498_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _16937_/B vssd1 vssd1 vccd1 vccd1 _16191_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12000__B _12154_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _20611_/B _12785_/B _15559_/D _15559_/C vssd1 vssd1 vccd1 vccd1 _12788_/B
+ sky130_fd_sc_hd__nand4_4
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11798__A1 _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17312_ _17312_/A vssd1 vssd1 vccd1 vccd1 _19482_/A sky130_fd_sc_hd__clkbuf_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22838__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14524_ _14540_/A _14540_/C _14540_/B vssd1 vssd1 vccd1 vccd1 _14524_/Y sky130_fd_sc_hd__a21oi_4
X_18292_ _18292_/A vssd1 vssd1 vccd1 vccd1 _18636_/A sky130_fd_sc_hd__clkbuf_4
X_11736_ _11502_/A _11503_/A _18093_/C _18093_/D vssd1 vssd1 vccd1 vccd1 _11736_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_109_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17243_ _17236_/X _17239_/Y _17242_/Y vssd1 vssd1 vccd1 vccd1 _17269_/B sky130_fd_sc_hd__o21ai_1
XFILLER_70_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14455_ _22658_/A _15435_/C _14448_/A vssd1 vssd1 vccd1 vccd1 _22670_/D sky130_fd_sc_hd__a21o_1
XFILLER_147_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11667_ _15435_/D vssd1 vssd1 vccd1 vccd1 _11667_/Y sky130_fd_sc_hd__inv_2
XFILLER_168_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13406_ _13262_/D _13438_/B _13413_/A _13413_/B vssd1 vssd1 vccd1 vccd1 _13406_/Y
+ sky130_fd_sc_hd__a22oi_1
X_17174_ _17323_/A _17122_/Y _17123_/X vssd1 vssd1 vccd1 vccd1 _17174_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11598_ _18156_/A vssd1 vssd1 vccd1 vccd1 _11598_/X sky130_fd_sc_hd__clkbuf_4
X_14386_ _20069_/A _14370_/X _14379_/X _21169_/A _14385_/X vssd1 vssd1 vccd1 vccd1
+ _14386_/X sky130_fd_sc_hd__a221o_1
X_16125_ _16119_/Y _16120_/Y _16122_/Y _16124_/X _12876_/X vssd1 vssd1 vccd1 vccd1
+ _16143_/A sky130_fd_sc_hd__o2111ai_2
XFILLER_170_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13337_ _13337_/A _13337_/B _13337_/C vssd1 vssd1 vccd1 vccd1 _13338_/B sky130_fd_sc_hd__and3_1
XFILLER_155_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12951__A _16947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16056_ _15997_/X _16053_/X _15972_/X _16110_/B _16055_/Y vssd1 vssd1 vccd1 vccd1
+ _16056_/Y sky130_fd_sc_hd__o2111ai_4
X_13268_ _21398_/B _21448_/B _21398_/A _21629_/B _13370_/A vssd1 vssd1 vccd1 vccd1
+ _13268_/X sky130_fd_sc_hd__a32o_1
XFILLER_68_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15007_ _14818_/A _14854_/X _15006_/Y vssd1 vssd1 vccd1 vccd1 _15007_/Y sky130_fd_sc_hd__o21ai_1
X_12219_ _12219_/A _12219_/B vssd1 vssd1 vccd1 vccd1 _12220_/B sky130_fd_sc_hd__nand2_1
X_13199_ _13199_/A _13199_/B vssd1 vssd1 vccd1 vccd1 _13210_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20588__A3 _20584_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19815_ _19815_/A _19815_/B vssd1 vssd1 vccd1 vccd1 _19817_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19746_ _19746_/A _19808_/B _19746_/C vssd1 vssd1 vccd1 vccd1 _19746_/Y sky130_fd_sc_hd__nand3_1
X_16958_ _20129_/B _17405_/A _17406_/A vssd1 vssd1 vccd1 vccd1 _16959_/B sky130_fd_sc_hd__and3_1
XFILLER_2_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14672__B1 _14670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_580 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15909_ _15909_/A _16192_/B _20502_/A _15988_/A vssd1 vssd1 vccd1 vccd1 _15978_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19677_ _19449_/Y _19574_/B _19676_/Y vssd1 vssd1 vccd1 vccd1 _19677_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16889_ _17076_/A _16889_/B _16889_/C vssd1 vssd1 vccd1 vccd1 _16892_/B sky130_fd_sc_hd__nand3_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17610__B1 _22899_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18628_ _18625_/X _18627_/Y _18629_/A _18830_/D vssd1 vssd1 vccd1 vccd1 _18633_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15205__C _15205_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18559_ _18559_/A _18559_/B vssd1 vssd1 vccd1 vccd1 _18561_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13778__A2 _13949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13632__D1 _21399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_650 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19902__A2 _19981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21570_ _21570_/A _21570_/B vssd1 vssd1 vccd1 vccd1 _21573_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17913__A1 _17226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20521_ _20337_/A _20376_/A _20367_/Y _20362_/Y vssd1 vssd1 vccd1 vccd1 _20522_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_162_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14118__A _14765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13022__A _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20452_ _20452_/A _20452_/B _20452_/C vssd1 vssd1 vccd1 vccd1 _20454_/B sky130_fd_sc_hd__and3_1
XFILLER_134_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20781__C _20972_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20276__A2 _12501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20383_ _20363_/Y _20365_/Y _20366_/Y _20382_/X vssd1 vssd1 vccd1 vccd1 _20403_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_174_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22122_ _22190_/B _22223_/A _22122_/C _22190_/A vssd1 vssd1 vccd1 vccd1 _22219_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18626__C1 _17401_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22053_ _22045_/Y _22048_/Y _22044_/X _22039_/Y vssd1 vssd1 vccd1 vccd1 _22099_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_142_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21004_ _21004_/A _21004_/B vssd1 vssd1 vccd1 vccd1 _22919_/D sky130_fd_sc_hd__xor2_2
XFILLER_101_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16101__B1 _11541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18641__A2 _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22955_ _22959_/CLK _22955_/D vssd1 vssd1 vccd1 vccd1 _22955_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20736__B1 _20735_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21906_ _21906_/A vssd1 vssd1 vccd1 vccd1 _22007_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_189_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15115__C _15115_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22886_ _22952_/CLK input80/X vssd1 vssd1 vccd1 vccd1 _22886_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16955__A2 _16227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21837_ _21837_/A _21837_/B _21837_/C _21837_/D vssd1 vssd1 vccd1 vccd1 _21838_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18157__A1 _11904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19354__B1 _19496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22229__B _22229_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12570_ _12335_/A _12403_/A _12493_/A vssd1 vssd1 vccd1 vccd1 _12571_/B sky130_fd_sc_hd__o21ai_4
XFILLER_11_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21768_ _21767_/X _21606_/X _21607_/X _21742_/A _21730_/A vssd1 vssd1 vccd1 vccd1
+ _21769_/B sky130_fd_sc_hd__o221ai_1
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12441__A2 _20130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20503__A3 _20359_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11521_ _11936_/A _18875_/C _11936_/C _18875_/D vssd1 vssd1 vccd1 vccd1 _11521_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14718__A1 _15114_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20719_ _20711_/Y _20712_/Y _20718_/X vssd1 vssd1 vccd1 vccd1 _20721_/B sky130_fd_sc_hd__o21ai_1
XFILLER_184_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21699_ _21930_/A _21834_/A _21815_/B _21702_/B vssd1 vssd1 vccd1 vccd1 _21704_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_196_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20972__B _20972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12729__B1 _12583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11452_ _11459_/A _11459_/B _11778_/A _11778_/B _11454_/A vssd1 vssd1 vccd1 vccd1
+ _11452_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14240_ _14198_/B _14198_/C _14198_/D _14234_/Y vssd1 vssd1 vccd1 vccd1 _14240_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22110__C1 _22173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14171_ _14054_/Y _14055_/X _14169_/X _14090_/Y _14170_/X vssd1 vssd1 vccd1 vccd1
+ _14172_/C sky130_fd_sc_hd__o221ai_1
XFILLER_164_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11383_ _11450_/A _11772_/A _11273_/X vssd1 vssd1 vccd1 vccd1 _11384_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__12771__A _12771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13122_ _13122_/A _13122_/B _13122_/C vssd1 vssd1 vccd1 vccd1 _13340_/A sky130_fd_sc_hd__nand3_4
XANTENNA_input61_A wb_dat_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13586__B _21805_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_875 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17930_ _19839_/C _17880_/A _17928_/D _17927_/A vssd1 vssd1 vccd1 vccd1 _17930_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _13158_/A _22723_/Q vssd1 vssd1 vccd1 vccd1 _13067_/B sky130_fd_sc_hd__nor2_1
XFILLER_124_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12004_ _12017_/A _12004_/B vssd1 vssd1 vccd1 vccd1 _12006_/A sky130_fd_sc_hd__nand2_1
X_17861_ _17861_/A _17861_/B vssd1 vssd1 vccd1 vccd1 _17910_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18632__A2 _17400_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17074__A _22896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19600_ _19607_/A _19607_/B _19608_/A vssd1 vssd1 vccd1 vccd1 _19605_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__16643__A1 _16613_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16812_ _16812_/A _16812_/B _16812_/C vssd1 vssd1 vccd1 vccd1 _16831_/A sky130_fd_sc_hd__nand3_2
XFILLER_94_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17792_ _17793_/B _17793_/C _22901_/Q vssd1 vssd1 vccd1 vccd1 _17866_/A sky130_fd_sc_hd__o21a_2
XFILLER_120_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19531_ _19458_/A _19458_/B _19398_/C _19530_/X vssd1 vssd1 vccd1 vccd1 _19540_/A
+ sky130_fd_sc_hd__a31oi_2
X_16743_ _16743_/A _16743_/B _16743_/C vssd1 vssd1 vccd1 vccd1 _16743_/X sky130_fd_sc_hd__and3_1
XFILLER_4_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15306__B _16256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13955_ _13951_/X _13926_/Y _14026_/C vssd1 vssd1 vccd1 vccd1 _13957_/A sky130_fd_sc_hd__o21ai_4
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1011 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12906_ _15901_/C vssd1 vssd1 vccd1 vccd1 _15804_/C sky130_fd_sc_hd__buf_2
X_19462_ _12111_/X _19160_/A _19323_/X vssd1 vssd1 vccd1 vccd1 _19462_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_34_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16674_ _17226_/A _17227_/A _16672_/X _16673_/Y _16665_/X vssd1 vssd1 vccd1 vccd1
+ _16675_/C sky130_fd_sc_hd__o221ai_1
XFILLER_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _13920_/A _13920_/B vssd1 vssd1 vccd1 vccd1 _13886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18413_ _18212_/A _18182_/A _18191_/A vssd1 vssd1 vccd1 vccd1 _18415_/B sky130_fd_sc_hd__a21bo_1
XFILLER_146_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15625_ _20461_/A vssd1 vssd1 vccd1 vccd1 _20471_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19393_ _19389_/X _19390_/Y _19398_/A vssd1 vssd1 vccd1 vccd1 _19394_/C sky130_fd_sc_hd__o21ai_1
XFILLER_36_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12837_ _20130_/A _20130_/B _22822_/Q vssd1 vssd1 vccd1 vccd1 _12838_/B sky130_fd_sc_hd__and3_1
XFILLER_146_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19345__B1 _17393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11850__A _18303_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _18337_/X _18343_/X _18340_/Y _19587_/D _15624_/A vssd1 vssd1 vccd1 vccd1
+ _18345_/C sky130_fd_sc_hd__o2111ai_4
X_15556_ _15838_/A _12716_/A _15498_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _15565_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_15_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _16067_/D vssd1 vssd1 vccd1 vccd1 _13024_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14507_ _13950_/X _13924_/A _14506_/Y vssd1 vssd1 vccd1 vccd1 _14512_/B sky130_fd_sc_hd__o21ai_1
X_11719_ _12046_/A vssd1 vssd1 vccd1 vccd1 _16226_/C sky130_fd_sc_hd__clkbuf_4
X_18275_ _18275_/A _18275_/B vssd1 vssd1 vccd1 vccd1 _18275_/X sky130_fd_sc_hd__and2_1
XANTENNA__15906__B1 _20502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11640__B1 _11626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15041__B _15046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15487_ _15539_/A _14439_/A _12046_/A _16226_/A vssd1 vssd1 vccd1 vccd1 _16218_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_187_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12699_ _20466_/B vssd1 vssd1 vccd1 vccd1 _20579_/C sky130_fd_sc_hd__buf_2
X_17226_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17226_/X sky130_fd_sc_hd__buf_2
XFILLER_159_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14438_ _14438_/A _16241_/D vssd1 vssd1 vccd1 vccd1 _14439_/D sky130_fd_sc_hd__nor2_1
Xinput10 wb_adr_i[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__14185__A2 _13930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput21 wb_adr_i[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_1
Xinput32 wb_adr_i[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput43 wb_dat_i[17] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput54 wb_dat_i[27] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__20258__A2 _12735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17157_ _17270_/A _17270_/B _17180_/B _17180_/C vssd1 vssd1 vccd1 vccd1 _17181_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput65 wb_dat_i[8] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_4
X_14369_ _22701_/Q vssd1 vssd1 vccd1 vccd1 _14369_/X sky130_fd_sc_hd__clkbuf_4
Xinput76 x[5] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16108_ _16586_/B _15899_/B _20134_/B _16166_/A _16107_/X vssd1 vssd1 vccd1 vccd1
+ _16160_/A sky130_fd_sc_hd__a32o_1
X_17088_ _16994_/Y _17431_/C _16997_/C _17087_/Y vssd1 vssd1 vccd1 vccd1 _17088_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17674__A3 _21083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18871__A2 _19091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11297__A _18691_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19464__A _19464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16039_ _16039_/A vssd1 vssd1 vccd1 vccd1 _16040_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_143_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13448__A1 _13050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19729_ _19735_/A vssd1 vssd1 vccd1 vccd1 _19731_/A sky130_fd_sc_hd__inv_2
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19584__B1 _17647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12120__B2 _12119_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22740_ _22751_/CLK _22740_/D vssd1 vssd1 vccd1 vccd1 _22740_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16398__B1 _16397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19630__C _19630_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20733__A3 _16078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22671_ _22949_/CLK _22671_/D vssd1 vssd1 vccd1 vccd1 _22671_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16328__A _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__A _11762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21622_ _13326_/Y _21958_/A _21742_/A _21614_/A _21766_/B vssd1 vssd1 vccd1 vccd1
+ _21622_/X sky130_fd_sc_hd__o311a_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13081__C1 _13304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__A2 _15325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21553_ _21553_/A _21553_/B _21553_/C _21553_/D vssd1 vssd1 vccd1 vccd1 _21556_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_193_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20504_ _15723_/A _20123_/X _15341_/X _20502_/X _20503_/Y vssd1 vssd1 vccd1 vccd1
+ _20504_/X sky130_fd_sc_hd__o311a_1
XFILLER_138_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21484_ _21466_/X _21467_/Y _21504_/B _21504_/C vssd1 vssd1 vccd1 vccd1 _21485_/A
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__19358__B _19358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13687__A _22672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20435_ _20554_/A _20554_/D _21066_/A _20434_/Y vssd1 vssd1 vccd1 vccd1 _20439_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_146_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16063__A _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20366_ _20366_/A _20366_/B _20366_/C vssd1 vssd1 vccd1 vccd1 _20366_/Y sky130_fd_sc_hd__nand3_1
XFILLER_134_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22105_ _22105_/A vssd1 vssd1 vccd1 vccd1 _22105_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20297_ _20298_/A _20298_/B _20319_/B vssd1 vssd1 vccd1 vccd1 _20300_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20406__C1 _20405_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22036_ _22036_/A _22036_/B _22036_/C vssd1 vssd1 vccd1 vccd1 _22064_/B sky130_fd_sc_hd__nand3_1
XFILLER_88_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11935__A _18292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22683__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13439__A1 _13434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13572__D _21938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18718__A _19176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22174__A2 _22173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13740_ _22758_/Q vssd1 vssd1 vccd1 vccd1 _13821_/A sky130_fd_sc_hd__inv_2
XANTENNA__22885__D input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22938_ _22948_/CLK _22938_/D vssd1 vssd1 vccd1 vccd1 _22938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16928__A2 _15940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17050__B2 _16644_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13671_ _13671_/A _13671_/B vssd1 vssd1 vccd1 vccd1 _13671_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22869_ _22916_/CLK _22869_/D vssd1 vssd1 vccd1 vccd1 _22869_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19327__B1 _12114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11670__A _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15410_ _11911_/A _15412_/A _15637_/A _12009_/A vssd1 vssd1 vccd1 vccd1 _15411_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_25_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14684__C _14684_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12622_ _12613_/Y _12602_/Y _12601_/Y _12584_/Y vssd1 vssd1 vccd1 vccd1 _12622_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_16390_ _16636_/B vssd1 vssd1 vccd1 vccd1 _16391_/C sky130_fd_sc_hd__inv_2
XFILLER_19_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20488__A2 _15939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15341_ _15409_/A vssd1 vssd1 vccd1 vccd1 _15341_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_145_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12553_ _12553_/A vssd1 vssd1 vccd1 vccd1 _12672_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_157_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18453__A _19199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18060_ _18029_/D _17839_/B _17839_/C _18023_/X _21081_/B vssd1 vssd1 vccd1 vccd1
+ _18063_/A sky130_fd_sc_hd__a311o_1
X_11504_ _11504_/A vssd1 vssd1 vccd1 vccd1 _11504_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15272_ _15279_/A _15271_/B _22878_/Q vssd1 vssd1 vccd1 vccd1 _15273_/B sky130_fd_sc_hd__a21bo_1
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12484_ _20250_/C _15774_/C _12792_/A _12487_/C vssd1 vssd1 vccd1 vccd1 _12484_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_185_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17011_ _17006_/Y _17008_/Y _17010_/X vssd1 vssd1 vccd1 vccd1 _17011_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14223_ _14195_/D _14222_/Y _14195_/A vssd1 vssd1 vccd1 vccd1 _14226_/A sky130_fd_sc_hd__a21boi_1
XFILLER_125_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11435_ _11675_/A _11325_/A _11311_/Y _11407_/B vssd1 vssd1 vccd1 vccd1 _11435_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21988__A2 _21522_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15116__A1 _15188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__B2 _11924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11366_ _11366_/A vssd1 vssd1 vccd1 vccd1 _12018_/A sky130_fd_sc_hd__buf_2
X_14154_ _14238_/A _14154_/B _14154_/C vssd1 vssd1 vccd1 vccd1 _14155_/B sky130_fd_sc_hd__nand3_1
XFILLER_98_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13105_ _13105_/A _13105_/B vssd1 vssd1 vccd1 vccd1 _13105_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14324__C1 _14323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16864__B2 _16740_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18962_ _18589_/A _18590_/A _18960_/C _18960_/B vssd1 vssd1 vccd1 vccd1 _19137_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_11297_ _18691_/C vssd1 vssd1 vccd1 vccd1 _18985_/C sky130_fd_sc_hd__buf_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _14085_/A _14085_/B vssd1 vssd1 vccd1 vccd1 _14085_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__12006__A _12006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17913_ _17226_/X _17227_/X _17849_/Y _17800_/Y vssd1 vssd1 vccd1 vccd1 _17960_/A
+ sky130_fd_sc_hd__o22ai_4
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _13036_/A _13036_/B vssd1 vssd1 vccd1 vccd1 _13038_/C sky130_fd_sc_hd__xor2_1
XFILLER_140_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18893_ _17083_/A _18856_/A _19771_/A _17313_/D vssd1 vssd1 vccd1 vccd1 _18893_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15962__D _17039_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11845__A _15792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17844_ _17785_/A _17785_/B _17954_/A vssd1 vssd1 vccd1 vccd1 _17845_/B sky130_fd_sc_hd__o21a_1
XANTENNA__16616__B2 _16310_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17235__C _20870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19015__C1 _19490_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17775_ _17855_/A _17855_/B _17778_/A vssd1 vssd1 vccd1 vccd1 _17775_/X sky130_fd_sc_hd__or3_2
XFILLER_19_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14987_ _15046_/A _15046_/B _14987_/C vssd1 vssd1 vccd1 vccd1 _14989_/A sky130_fd_sc_hd__and3_1
XFILLER_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19514_ _19356_/X _19363_/Y _19369_/Y _19379_/B vssd1 vssd1 vccd1 vccd1 _19514_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__17532__A _17532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16726_ _16724_/X _16725_/Y _16743_/C _16743_/A vssd1 vssd1 vccd1 vccd1 _16726_/Y
+ sky130_fd_sc_hd__o211ai_4
X_13938_ _14465_/A vssd1 vssd1 vccd1 vccd1 _14770_/A sky130_fd_sc_hd__buf_2
XFILLER_62_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_222 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19445_ _19440_/X _19447_/A _22917_/Q vssd1 vssd1 vccd1 vccd1 _19445_/Y sky130_fd_sc_hd__o21bai_1
X_16657_ _16657_/A _16657_/B _16657_/C vssd1 vssd1 vccd1 vccd1 _16659_/B sky130_fd_sc_hd__nand3_4
X_13869_ _22759_/Q _13869_/B _13869_/C vssd1 vssd1 vccd1 vccd1 _13875_/A sky130_fd_sc_hd__nand3b_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15608_ _15608_/A _22700_/Q _15608_/C vssd1 vssd1 vccd1 vccd1 _20461_/B sky130_fd_sc_hd__nand3_2
XFILLER_72_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19376_ _19376_/A _19376_/B _19376_/C vssd1 vssd1 vccd1 vccd1 _19457_/A sky130_fd_sc_hd__nand3_2
XFILLER_195_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19869__A1 _19836_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16588_ _16265_/A _16265_/B _16263_/C _16263_/D vssd1 vssd1 vccd1 vccd1 _16588_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_72_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18327_ _18495_/A _18495_/B _18326_/Y vssd1 vssd1 vccd1 vccd1 _18327_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15539_ _15539_/A vssd1 vssd1 vccd1 vccd1 _18258_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__15987__A _16261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _18258_/A _18258_/B vssd1 vssd1 vccd1 vccd1 _18589_/A sky130_fd_sc_hd__nor2_1
XFILLER_163_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17209_ _17513_/C vssd1 vssd1 vccd1 vccd1 _17210_/B sky130_fd_sc_hd__inv_2
XANTENNA__12169__B2 _12168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18189_ _18163_/Y _18404_/A _18113_/Y _18114_/X vssd1 vssd1 vccd1 vccd1 _18189_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__20636__C1 _20737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20220_ _20093_/B _20219_/Y _20090_/Y vssd1 vssd1 vccd1 vccd1 _20224_/B sky130_fd_sc_hd__o21ai_4
XFILLER_162_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18844__A2 _19161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18810__B _19507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15658__A2 _16397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__A2 _11503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19194__A _19194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20151_ _12864_/B _12862_/B _12851_/Y _12843_/X vssd1 vssd1 vccd1 vccd1 _20158_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_170_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16611__A _16611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14866__B1 _14861_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20082_ _20089_/A _20089_/B _20338_/C vssd1 vssd1 vccd1 vccd1 _20219_/B sky130_fd_sc_hd__nand3_2
XANTENNA__17426__B _20854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20133__A _20133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14131__A _14686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16083__A2 _11563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19557__B1 _19211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17442__A _17442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14492__A1_N _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19021__A2 _19015_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ _20985_/B _20985_/C _20985_/A vssd1 vssd1 vccd1 vccd1 _20986_/A sky130_fd_sc_hd__a21oi_1
XFILLER_150_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14785__B _14785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22723_ _22725_/CLK _22723_/D vssd1 vssd1 vccd1 vccd1 _22723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16058__A _20249_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15043__B1 _15175_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22654_ _22814_/Q input58/X _22656_/S vssd1 vssd1 vccd1 vccd1 _22655_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16791__B1 _19358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21605_ _21645_/B vssd1 vssd1 vccd1 vccd1 _21763_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__21667__A1 _21269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22585_ _22585_/A vssd1 vssd1 vccd1 vccd1 _22783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21536_ _21404_/A _21404_/B _21403_/A _21401_/Y vssd1 vssd1 vccd1 vccd1 _21536_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_193_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15897__A2 _15504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21467_ _21467_/A _21467_/B vssd1 vssd1 vccd1 vccd1 _21467_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11907__A1 _11904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20418_ _20420_/A _20545_/A _20414_/X _20429_/C vssd1 vssd1 vccd1 vccd1 _20423_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19493__C1 _19490_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21398_ _21398_/A _21398_/B _21445_/A _21665_/D vssd1 vssd1 vccd1 vccd1 _21399_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17039__D _17039_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12580__A1 _12576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20349_ _20349_/A vssd1 vssd1 vccd1 vccd1 _20366_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1087 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22019_ _22016_/X _22017_/X _22018_/Y vssd1 vssd1 vccd1 vccd1 _22021_/A sky130_fd_sc_hd__a21o_1
X_14910_ _14906_/X _14816_/B _14909_/Y vssd1 vssd1 vccd1 vccd1 _14912_/A sky130_fd_sc_hd__a21boi_1
XFILLER_49_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15890_ _15890_/A vssd1 vssd1 vccd1 vccd1 _15890_/X sky130_fd_sc_hd__buf_2
XFILLER_75_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14041__A _14220_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16074__A2 _12294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input24_A wb_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ _14756_/B _14839_/Y _14840_/Y vssd1 vssd1 vccd1 vccd1 _14842_/B sky130_fd_sc_hd__o21ai_2
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17560_ _18659_/D vssd1 vssd1 vccd1 vccd1 _19013_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__12096__B1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14772_ _22766_/Q vssd1 vssd1 vccd1 vccd1 _14869_/C sky130_fd_sc_hd__inv_2
X_11984_ _11984_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _11984_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13832__A1 _13737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16511_ _15997_/C _16491_/B _16964_/A _15810_/C _16231_/X vssd1 vssd1 vccd1 vccd1
+ _16512_/B sky130_fd_sc_hd__o2111a_1
XFILLER_186_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13723_ _22754_/Q _22752_/Q vssd1 vssd1 vccd1 vccd1 _13810_/A sky130_fd_sc_hd__nor2_2
X_17491_ _17491_/A _17491_/B _17491_/C vssd1 vssd1 vccd1 vccd1 _17493_/A sky130_fd_sc_hd__nand3_1
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11843__B1 _11899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19230_ _19400_/A _19244_/A vssd1 vssd1 vccd1 vccd1 _19246_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16442_ _16206_/X _15879_/X _16432_/Y _16433_/Y _16210_/Y vssd1 vssd1 vccd1 vccd1
+ _16442_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_108_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13654_ _13657_/B _21874_/A _13657_/A _13664_/D vssd1 vssd1 vccd1 vccd1 _13655_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19161_ _19161_/A vssd1 vssd1 vccd1 vccd1 _19792_/A sky130_fd_sc_hd__buf_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _15799_/A _15799_/B _20463_/C _12938_/A _20456_/C vssd1 vssd1 vccd1 vccd1
+ _12605_/Y sky130_fd_sc_hd__a32oi_4
X_16373_ _16371_/Y _16372_/X _15678_/A _15678_/C vssd1 vssd1 vccd1 vccd1 _16373_/Y
+ sky130_fd_sc_hd__o211ai_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13104__B _21595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13585_ _21195_/B vssd1 vssd1 vccd1 vccd1 _21878_/C sky130_fd_sc_hd__buf_2
XFILLER_185_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _18278_/B vssd1 vssd1 vccd1 vccd1 _18184_/B sky130_fd_sc_hd__clkbuf_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _15324_/A vssd1 vssd1 vccd1 vccd1 _15426_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19092_ _18907_/A _18907_/B _18907_/C vssd1 vssd1 vccd1 vccd1 _19092_/Y sky130_fd_sc_hd__a21oi_1
X_12536_ _20134_/A _15776_/D _12515_/A _16759_/A _20128_/A vssd1 vssd1 vccd1 vccd1
+ _12536_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_129_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17877__A3 _21048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18043_ _18042_/Y _18048_/A _18040_/A vssd1 vssd1 vccd1 vccd1 _18049_/B sky130_fd_sc_hd__a21oi_2
XFILLER_145_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15255_ _14990_/X _15217_/B _15253_/Y _15266_/A vssd1 vssd1 vccd1 vccd1 _15257_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_173_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12467_ _12467_/A _15466_/C _22821_/Q vssd1 vssd1 vccd1 vccd1 _12988_/C sky130_fd_sc_hd__nand3_2
XFILLER_138_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14206_ _14143_/X _14057_/A _14203_/X _14205_/Y vssd1 vssd1 vccd1 vccd1 _14206_/Y
+ sky130_fd_sc_hd__o22ai_2
X_11418_ _11418_/A vssd1 vssd1 vccd1 vccd1 _11430_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_193_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15186_ _15186_/A _15186_/B _15186_/C _15186_/D vssd1 vssd1 vccd1 vccd1 _15186_/X
+ sky130_fd_sc_hd__and4_1
X_12398_ _15466_/B _15466_/C vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__nand2_2
XFILLER_125_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14137_ _13923_/X _14561_/C _14231_/C vssd1 vssd1 vccd1 vccd1 _14154_/B sky130_fd_sc_hd__o21ai_1
X_11349_ _18115_/C vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__clkbuf_4
X_19994_ _19994_/A _19994_/B vssd1 vssd1 vccd1 vccd1 _19995_/B sky130_fd_sc_hd__nand2_1
XFILLER_152_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16431__A _16431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17246__B _17532_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18945_ _18945_/A _18945_/B _18945_/C vssd1 vssd1 vccd1 vccd1 _18952_/B sky130_fd_sc_hd__nand3_1
X_14068_ _14510_/A _14126_/B _14868_/C vssd1 vssd1 vccd1 vccd1 _14068_/X sky130_fd_sc_hd__and3_1
XANTENNA__11575__A _11899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ _15577_/D _12711_/X _13017_/X _12989_/B _13016_/X vssd1 vssd1 vccd1 vccd1
+ _13019_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_79_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18876_ _18876_/A _18876_/B _18876_/C vssd1 vssd1 vccd1 vccd1 _18983_/A sky130_fd_sc_hd__nand3_1
XANTENNA__11294__B _11404_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17827_ _17827_/A _17890_/A _17827_/C vssd1 vssd1 vccd1 vccd1 _17890_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19461__B _19461_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13790__A _22874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17758_ _17662_/B _17662_/A _17660_/B vssd1 vssd1 vccd1 vccd1 _17760_/A sky130_fd_sc_hd__o21ai_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16709_ _11904_/A _11905_/A _16715_/A _20098_/D vssd1 vssd1 vccd1 vccd1 _16709_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_81_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17689_ _17626_/X _17627_/X _17697_/B _17690_/A vssd1 vssd1 vccd1 vccd1 _17693_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21215__C _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19428_ _19428_/A _19561_/A vssd1 vssd1 vccd1 vccd1 _19663_/A sky130_fd_sc_hd__nand2_1
XFILLER_168_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19306__A3 _19983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19359_ _19359_/A vssd1 vssd1 vccd1 vccd1 _19359_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18514__A1 _16241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15328__A1 _12090_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22370_ _22426_/A vssd1 vssd1 vccd1 vccd1 _22439_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__16325__B _16325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21321_ _21321_/A vssd1 vssd1 vccd1 vccd1 _21386_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20872__A2 _20806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21252_ _21399_/A _21442_/A _21251_/B _21251_/A vssd1 vssd1 vccd1 vccd1 _21299_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20203_ _20116_/A _20197_/Y _20202_/Y vssd1 vssd1 vccd1 vccd1 _20268_/A sky130_fd_sc_hd__a21oi_1
XFILLER_190_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21183_ _21220_/A vssd1 vssd1 vccd1 vccd1 _21183_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20134_ _20134_/A _20134_/B _20134_/C vssd1 vssd1 vccd1 vccd1 _20134_/X sky130_fd_sc_hd__and3_1
XFILLER_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19652__A _19652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20065_ _20064_/Y _20304_/A _13041_/Y vssd1 vssd1 vccd1 vccd1 _20065_/Y sky130_fd_sc_hd__a21oi_4
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17789__C1 _17959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16056__A2 _16053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12078__B1 _11909_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ _20923_/B _20936_/D _20966_/X vssd1 vssd1 vccd1 vccd1 _20967_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22706_ _22738_/CLK _22706_/D vssd1 vssd1 vccd1 vccd1 _22706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20898_ _20834_/X _20835_/X _20994_/A _20994_/B _20906_/C vssd1 vssd1 vccd1 vccd1
+ _20961_/B sky130_fd_sc_hd__o221ai_4
XANTENNA__13578__B1 _13662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21422__A _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22637_ _22806_/Q input49/X _22641_/S vssd1 vssd1 vccd1 vccd1 _22638_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22871__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _13370_/A vssd1 vssd1 vccd1 vccd1 _13650_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13453__A2_N _21750_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22568_ _22568_/A vssd1 vssd1 vccd1 vccd1 _22775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ _16319_/A _12402_/A _12319_/Y _12320_/Y vssd1 vssd1 vccd1 vccd1 _16268_/A
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__20642__A2_N _20737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21519_ _21376_/X _13343_/X _13366_/Y _21179_/B vssd1 vssd1 vccd1 vccd1 _21519_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_182_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22499_ _22499_/A vssd1 vssd1 vccd1 vccd1 _22508_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_108_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15040_ _15040_/A _15040_/B vssd1 vssd1 vccd1 vccd1 _15175_/D sky130_fd_sc_hd__xor2_4
XFILLER_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12252_ _11834_/Y _11832_/Y _18239_/B vssd1 vssd1 vccd1 vccd1 _18272_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__19466__C1 _19694_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12183_ _18208_/A _12123_/B _12123_/C vssd1 vssd1 vccd1 vccd1 _12183_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_122_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13594__B _21750_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16991_ _16822_/A _16822_/B _16822_/C _16831_/C vssd1 vssd1 vccd1 vccd1 _16991_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_68_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11395__A _11395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18730_ _18527_/B _18527_/C _18527_/A _18555_/B vssd1 vssd1 vccd1 vccd1 _18730_/Y
+ sky130_fd_sc_hd__a31oi_2
X_15942_ _15918_/X _15941_/X _15725_/Y _15935_/X vssd1 vssd1 vccd1 vccd1 _15942_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18661_ _18661_/A _18661_/B _18661_/C vssd1 vssd1 vccd1 vccd1 _18662_/A sky130_fd_sc_hd__nand3_1
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15873_ _15758_/A _15758_/B _15758_/C _15862_/Y vssd1 vssd1 vccd1 vccd1 _15873_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_23_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14058__B2 _14057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17612_ _17713_/A _17611_/X _22899_/Q vssd1 vssd1 vccd1 vccd1 _17612_/Y sky130_fd_sc_hd__a21boi_1
X_14824_ _14825_/C _14902_/B _14825_/A vssd1 vssd1 vccd1 vccd1 _14916_/A sky130_fd_sc_hd__a21o_1
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18592_ _18437_/Y _18586_/B _18591_/X vssd1 vssd1 vccd1 vccd1 _18592_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12608__A2 _12607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ _17252_/Y _17535_/A _17408_/B _17394_/Y vssd1 vssd1 vccd1 vccd1 _17544_/C
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__21879__A1 _21383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _14836_/A _14749_/B _14751_/B vssd1 vssd1 vccd1 vccd1 _14756_/C sky130_fd_sc_hd__a21o_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _11799_/A _11799_/B _11799_/C _11965_/X _11966_/X vssd1 vssd1 vccd1 vccd1
+ _11967_/Y sky130_fd_sc_hd__a32oi_2
XFILLER_189_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11292__A1 _22954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16129__C _16129_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ _22767_/Q vssd1 vssd1 vccd1 vccd1 _13845_/B sky130_fd_sc_hd__buf_2
X_17474_ _17474_/A _17474_/B _17474_/C vssd1 vssd1 vccd1 vccd1 _17490_/A sky130_fd_sc_hd__nand3_1
X_14686_ _14785_/A _14686_/B _14786_/C vssd1 vssd1 vccd1 vccd1 _14686_/X sky130_fd_sc_hd__and3_1
XFILLER_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11898_ _11899_/A _11899_/B _11902_/B _11902_/C vssd1 vssd1 vccd1 vccd1 _11900_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16425_ _16686_/A _16686_/B _16424_/Y vssd1 vssd1 vccd1 vccd1 _16664_/A sky130_fd_sc_hd__a21oi_1
X_19213_ _19195_/Y _19218_/B _19200_/B vssd1 vssd1 vccd1 vccd1 _19213_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_177_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13637_ _13666_/A _13666_/B _13666_/C vssd1 vssd1 vccd1 vccd1 _13637_/Y sky130_fd_sc_hd__nand3_1
XFILLER_158_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21676__A_N _21680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19144_ _22914_/Q _18967_/B _19143_/Y vssd1 vssd1 vccd1 vccd1 _19145_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__15330__A _20130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16356_ _20471_/A vssd1 vssd1 vccd1 vccd1 _20854_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__20593__D _20593_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13568_ _21741_/B _21250_/C _21250_/A _21498_/D _13572_/B vssd1 vssd1 vccd1 vccd1
+ _13573_/A sky130_fd_sc_hd__a32o_1
XFILLER_173_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15307_ _12500_/A _12501_/A _15557_/A _11734_/A vssd1 vssd1 vccd1 vccd1 _15308_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_121_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11595__A2 _15905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19075_ _19148_/A _19148_/B _19148_/C vssd1 vssd1 vccd1 vccd1 _19096_/A sky130_fd_sc_hd__nand3_1
X_12519_ _12549_/A _12519_/B _12669_/A vssd1 vssd1 vccd1 vccd1 _12522_/A sky130_fd_sc_hd__nand3b_4
XFILLER_185_594 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16287_ _16287_/A _16287_/B vssd1 vssd1 vccd1 vccd1 _16287_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13499_ _13493_/A _21280_/A _13493_/B vssd1 vssd1 vccd1 vccd1 _13499_/X sky130_fd_sc_hd__a21o_1
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18026_ _19945_/B vssd1 vssd1 vccd1 vccd1 _19418_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15238_ _15238_/A _15238_/B vssd1 vssd1 vccd1 vccd1 _15240_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _15169_/A _15169_/B _15181_/B vssd1 vssd1 vccd1 vccd1 _15171_/A sky130_fd_sc_hd__or3_1
XFILLER_158_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19977_ _19977_/A _19977_/B _22924_/Q vssd1 vssd1 vccd1 vccd1 _19977_/X sky130_fd_sc_hd__and3_1
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18928_ _18748_/B _18737_/X _18732_/Y _18725_/X vssd1 vssd1 vccd1 vccd1 _18932_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_80_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19224__A2 _19023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12847__A2 _20358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18859_ _19480_/A _19481_/A vssd1 vssd1 vccd1 vccd1 _19313_/A sky130_fd_sc_hd__nand2_4
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21870_ _21767_/X _21970_/A _21880_/A vssd1 vssd1 vccd1 vccd1 _21875_/A sky130_fd_sc_hd__o21ai_1
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20790__A1 _16579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20130__B _20130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20821_ _20822_/A _20822_/B _20822_/C vssd1 vssd1 vccd1 vccd1 _20890_/B sky130_fd_sc_hd__a21o_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22894__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1042 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20752_ _20758_/B vssd1 vssd1 vccd1 vccd1 _20830_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11822__A3 _11821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22338__A _22338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20683_ _20683_/A _20683_/B vssd1 vssd1 vccd1 vccd1 _20686_/A sky130_fd_sc_hd__nand2_1
XFILLER_149_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22057__B _22057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22422_ _22711_/Q input50/X _22424_/S vssd1 vssd1 vccd1 vccd1 _22423_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12583__B _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22353_ _22354_/A _22354_/B _22687_/Q vssd1 vssd1 vccd1 vccd1 _22356_/B sky130_fd_sc_hd__o21bai_1
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20845__A2 _15919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21304_ _13112_/Y _21469_/B _21583_/B _21304_/D vssd1 vssd1 vccd1 vccd1 _21307_/A
+ sky130_fd_sc_hd__nand4b_2
X_22284_ _22300_/B _22300_/A _22284_/C vssd1 vssd1 vccd1 vccd1 _22285_/B sky130_fd_sc_hd__and3_1
XFILLER_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21235_ _13314_/B _13314_/C _13314_/A vssd1 vssd1 vccd1 vccd1 _21235_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13695__A _22872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16277__A2 _17434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21166_ _21162_/A _21162_/B _21164_/Y _21165_/Y vssd1 vssd1 vccd1 vccd1 _21167_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_120_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20117_ _20119_/A _20119_/B vssd1 vssd1 vccd1 vccd1 _20118_/A sky130_fd_sc_hd__nand2_1
X_21097_ _21097_/A vssd1 vssd1 vccd1 vccd1 _21097_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20048_ _20059_/A _20059_/B _22927_/Q vssd1 vssd1 vccd1 vccd1 _20049_/C sky130_fd_sc_hd__o21ai_1
XFILLER_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_902 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _12843_/X _12851_/Y _12862_/B _12864_/B vssd1 vssd1 vccd1 vccd1 _12872_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_171_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19518__A3 _19981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _16014_/A vssd1 vssd1 vccd1 vccd1 _11821_/X sky130_fd_sc_hd__buf_4
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21999_ _21996_/A _21996_/B _21997_/Y _21998_/X vssd1 vssd1 vccd1 vccd1 _21999_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20975__B _20975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17630__A _19772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14540_/A _14540_/B _14540_/C vssd1 vssd1 vccd1 vccd1 _14541_/D sky130_fd_sc_hd__nand3_1
XFILLER_121_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11752_ _11708_/Y _11935_/C _11751_/X vssd1 vssd1 vccd1 vccd1 _11752_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18445__B _18797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _13987_/X _13984_/Y _14470_/X vssd1 vssd1 vccd1 vccd1 _14472_/C sky130_fd_sc_hd__a21o_1
XFILLER_42_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11683_ _11702_/A vssd1 vssd1 vccd1 vccd1 _12117_/A sky130_fd_sc_hd__buf_2
XANTENNA__12774__A _12774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16246__A _19197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16210_ _16210_/A _16210_/B _16210_/C _16210_/D vssd1 vssd1 vccd1 vccd1 _16210_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_81_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13422_ _13623_/A _22041_/B vssd1 vssd1 vccd1 vccd1 _13487_/A sky130_fd_sc_hd__nand2_1
X_17190_ _17188_/Y _16982_/A _17189_/Y _16845_/A vssd1 vssd1 vccd1 vccd1 _17190_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_167_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _16119_/Y _16120_/Y _15812_/D _16122_/Y vssd1 vssd1 vccd1 vccd1 _16141_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13353_ _13340_/Y _13341_/X _13352_/Y vssd1 vssd1 vccd1 vccd1 _13353_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_167_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18461__A _18464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12304_ _12387_/B _12824_/A _16328_/A _12273_/B vssd1 vssd1 vccd1 vccd1 _12904_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__15712__A1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16072_ _16126_/A _16126_/B _16126_/C vssd1 vssd1 vccd1 vccd1 _16072_/X sky130_fd_sc_hd__and3_1
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13284_ _13481_/A _13481_/B vssd1 vssd1 vccd1 vccd1 _13289_/A sky130_fd_sc_hd__xor2_1
XFILLER_155_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19900_ _19900_/A vssd1 vssd1 vccd1 vccd1 _19901_/B sky130_fd_sc_hd__clkbuf_2
X_15023_ _15213_/A _15023_/B vssd1 vssd1 vccd1 vccd1 _15023_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12526__B2 _22824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12235_ _15536_/A _12235_/B _22660_/B vssd1 vssd1 vccd1 vccd1 _15445_/B sky130_fd_sc_hd__nand3_1
XFILLER_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17465__A1 _17083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19831_ _19831_/A _19887_/B vssd1 vssd1 vccd1 vccd1 _19832_/A sky130_fd_sc_hd__and2_1
XFILLER_151_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12166_ _19016_/B _19016_/C vssd1 vssd1 vccd1 vccd1 _18855_/A sky130_fd_sc_hd__nand2_1
XFILLER_150_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19762_ _19814_/B vssd1 vssd1 vccd1 vccd1 _19764_/C sky130_fd_sc_hd__inv_2
X_16974_ _16768_/B _16768_/C _16768_/A _16777_/A _16971_/B vssd1 vssd1 vccd1 vccd1
+ _16980_/A sky130_fd_sc_hd__a32oi_4
XANTENNA__11556__C _11712_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ _11859_/A _11861_/A _15557_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _12097_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_77_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18713_ _18713_/A _18713_/B _18836_/A vssd1 vssd1 vccd1 vccd1 _18741_/C sky130_fd_sc_hd__nand3_2
XANTENNA__21013__A2 _20972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15925_ _16009_/C _15898_/Y _16010_/B vssd1 vssd1 vccd1 vccd1 _15967_/B sky130_fd_sc_hd__o21ai_1
XFILLER_110_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19693_ _12207_/X _19624_/A _19692_/Y vssd1 vssd1 vccd1 vccd1 _19697_/D sky130_fd_sc_hd__o21ai_2
Xinput8 wb_adr_i[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12949__A _20579_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11853__A _18107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15325__A _15325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18644_ _18465_/X _18467_/Y _18474_/B _18462_/A vssd1 vssd1 vccd1 vccd1 _18646_/C
+ sky130_fd_sc_hd__a2bb2o_2
X_15856_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15856_/Y sky130_fd_sc_hd__clkinv_2
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14807_ _13923_/X _14562_/X _14708_/D vssd1 vssd1 vccd1 vccd1 _14815_/B sky130_fd_sc_hd__o21ai_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18575_ _18574_/X _18575_/B _18761_/A vssd1 vssd1 vccd1 vccd1 _18578_/B sky130_fd_sc_hd__nand3b_1
X_15787_ _16192_/B _12689_/A _17133_/A _15991_/D vssd1 vssd1 vccd1 vccd1 _15788_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18717__A1 _18681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ _12997_/Y _12963_/D _12998_/X vssd1 vssd1 vccd1 vccd1 _13037_/A sky130_fd_sc_hd__o21ai_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18636__A _18636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16991__A3 _16822_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17526_ _17634_/A vssd1 vssd1 vccd1 vccd1 _17526_/X sky130_fd_sc_hd__clkbuf_4
X_14738_ _14738_/A _14738_/B vssd1 vssd1 vccd1 vccd1 _14740_/C sky130_fd_sc_hd__nand2_1
XANTENNA__16728__B1 _15932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17457_ _17457_/A _17523_/C _17457_/C _17457_/D vssd1 vssd1 vccd1 vccd1 _17458_/C
+ sky130_fd_sc_hd__nand4_1
X_14669_ _14669_/A vssd1 vssd1 vccd1 vccd1 _14670_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12684__A _20593_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16408_ _15877_/X _16210_/B _15957_/C vssd1 vssd1 vccd1 vccd1 _16408_/Y sky130_fd_sc_hd__o21ai_2
X_17388_ _17388_/A vssd1 vssd1 vccd1 vccd1 _17388_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19127_ _19121_/B _19122_/Y _19114_/X vssd1 vssd1 vccd1 vccd1 _19129_/B sky130_fd_sc_hd__a21o_1
X_16339_ _16301_/Y _16305_/Y _16309_/Y vssd1 vssd1 vccd1 vccd1 _16617_/A sky130_fd_sc_hd__a21o_2
XFILLER_173_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18371__A _18371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19693__A2 _19624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19058_ _18798_/Y _18804_/B _19052_/Y vssd1 vssd1 vccd1 vccd1 _19063_/A sky130_fd_sc_hd__a21boi_1
XFILLER_146_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18009_ _17851_/X _17850_/Y _17866_/A _17864_/Y vssd1 vssd1 vccd1 vccd1 _18009_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21020_ _21020_/A _21020_/B vssd1 vssd1 vccd1 vccd1 _21021_/B sky130_fd_sc_hd__xor2_1
XANTENNA__16322__C _22700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22621__A _22643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1071 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15219__B1 _15188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20212__B1 _20341_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21922_ _21922_/A _21922_/B vssd1 vssd1 vccd1 vccd1 _21922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21853_ _21853_/A vssd1 vssd1 vccd1 vccd1 _21853_/X sky130_fd_sc_hd__buf_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18708__A1 _12009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17450__A _17457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20804_ _20844_/A _15919_/X _20717_/B _20717_/A _20683_/B vssd1 vssd1 vccd1 vccd1
+ _20804_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12453__B1 _20323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20515__A1 _20514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21784_ _21846_/A _21763_/A _21763_/B vssd1 vssd1 vccd1 vccd1 _21784_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20735_ _20735_/A _20735_/B vssd1 vssd1 vccd1 vccd1 _20735_/Y sky130_fd_sc_hd__nand2_1
XFILLER_196_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17392__B1 _17532_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16066__A _18328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12594__A _15558_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_678 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15942__A1 _15918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15401__C _16712_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20666_ _20768_/A _22934_/Q _20768_/C vssd1 vssd1 vccd1 vccd1 _20666_/X sky130_fd_sc_hd__and3_1
XANTENNA__15942__B2 _15935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22405_ _20069_/A input41/X _22413_/S vssd1 vssd1 vccd1 vccd1 _22406_/A sky130_fd_sc_hd__mux2_1
X_20597_ _20603_/C vssd1 vssd1 vccd1 vccd1 _20702_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_87_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22336_ _22336_/A vssd1 vssd1 vccd1 vccd1 _22341_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13705__B1 _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22267_ _22302_/A _22302_/B _22266_/Y vssd1 vssd1 vccd1 vccd1 _22308_/C sky130_fd_sc_hd__o21ai_1
XFILLER_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12020_ _11972_/Y _11976_/Y _11986_/A vssd1 vssd1 vccd1 vccd1 _12020_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_183_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11657__B _15435_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21218_ _21638_/C vssd1 vssd1 vccd1 vccd1 _21219_/C sky130_fd_sc_hd__clkbuf_2
X_22198_ _22215_/A _22215_/B vssd1 vssd1 vccd1 vccd1 _22198_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_105_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21149_ _21149_/A vssd1 vssd1 vccd1 vccd1 _21165_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__22888__D input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14130__B1 _13873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13971_ _13907_/X _13970_/X _14581_/B _14699_/B vssd1 vssd1 vccd1 vccd1 _14475_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_24_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15710_ _16712_/C vssd1 vssd1 vccd1 vccd1 _15711_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12922_ _16059_/A vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__buf_2
XFILLER_111_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16690_ _16690_/A _22891_/Q _16690_/C vssd1 vssd1 vccd1 vccd1 _16697_/A sky130_fd_sc_hd__nand3_1
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15641_ _15347_/X _15343_/X _15636_/Y _15640_/Y _15336_/Y vssd1 vssd1 vccd1 vccd1
+ _15660_/C sky130_fd_sc_hd__o2111ai_4
XANTENNA__17080__C1 _17462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ _12853_/A _12859_/B vssd1 vssd1 vccd1 vccd1 _12856_/A sky130_fd_sc_hd__nand2_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _17421_/A _17422_/A _11345_/X _11351_/X vssd1 vssd1 vccd1 vccd1 _18360_/X
+ sky130_fd_sc_hd__a211o_1
X_11804_ _11964_/A _11964_/B _11964_/C vssd1 vssd1 vccd1 vccd1 _11810_/C sky130_fd_sc_hd__nand3_1
XFILLER_33_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _19465_/A vssd1 vssd1 vccd1 vccd1 _17436_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15799__B _15799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12784_ _12374_/A _12374_/B _12391_/Y vssd1 vssd1 vccd1 vccd1 _12792_/B sky130_fd_sc_hd__o21ai_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17311_/A _17311_/B _17311_/C vssd1 vssd1 vccd1 vccd1 _17311_/X sky130_fd_sc_hd__and3_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11798__A2 _11639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14523_/A _14523_/B vssd1 vssd1 vccd1 vccd1 _14540_/B sky130_fd_sc_hd__nand2_2
XFILLER_159_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18291_ _18291_/A _18291_/B _18291_/C vssd1 vssd1 vccd1 vccd1 _18305_/D sky130_fd_sc_hd__nand3_4
X_11735_ _15559_/B vssd1 vssd1 vccd1 vccd1 _18093_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17242_ _17242_/A _17242_/B vssd1 vssd1 vccd1 vccd1 _17242_/Y sky130_fd_sc_hd__nand2_1
X_14454_ _22658_/A _15435_/B _14448_/A vssd1 vssd1 vccd1 vccd1 _22669_/D sky130_fd_sc_hd__a21o_1
X_11666_ _16257_/A vssd1 vssd1 vccd1 vccd1 _11666_/X sky130_fd_sc_hd__buf_4
X_13405_ _13413_/B _13413_/A vssd1 vssd1 vccd1 vccd1 _13405_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17173_ _17178_/A _17178_/B _17173_/C _17173_/D vssd1 vssd1 vccd1 vccd1 _17177_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19287__A _22916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14385_ _18258_/A _14381_/X _14382_/X _14361_/X _14863_/C vssd1 vssd1 vccd1 vccd1
+ _14385_/X sky130_fd_sc_hd__a32o_1
XANTENNA__12009__A _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11597_ _11533_/B _11578_/Y _11529_/Y vssd1 vssd1 vccd1 vccd1 _11600_/B sky130_fd_sc_hd__o21ai_1
X_16124_ _19336_/A vssd1 vssd1 vccd1 vccd1 _16124_/X sky130_fd_sc_hd__buf_4
X_13336_ _13329_/X _13337_/B _13337_/C vssd1 vssd1 vccd1 vccd1 _21234_/A sky130_fd_sc_hd__a21oi_1
XFILLER_41_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11848__A _15714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16055_ _15900_/B _15983_/Y _15997_/X _16005_/A vssd1 vssd1 vccd1 vccd1 _16055_/Y
+ sky130_fd_sc_hd__o211ai_4
X_13267_ _22847_/Q vssd1 vssd1 vccd1 vccd1 _21448_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_108_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15006_ _15006_/A _15006_/B _15006_/C vssd1 vssd1 vccd1 vccd1 _15006_/Y sky130_fd_sc_hd__nand3_1
XFILLER_155_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12218_ _18830_/A _12052_/A _19772_/C _12217_/X vssd1 vssd1 vccd1 vccd1 _12221_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13198_ _21173_/A _21609_/B _21173_/C vssd1 vssd1 vccd1 vccd1 _13199_/B sky130_fd_sc_hd__nand3_1
XANTENNA__22441__A input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15449__B1 _12117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19814_ _19814_/A _19814_/B _19814_/C vssd1 vssd1 vccd1 vccd1 _19815_/B sky130_fd_sc_hd__nor3_1
XFILLER_151_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12149_ _12146_/Y _12148_/Y _11619_/B vssd1 vssd1 vccd1 vccd1 _18128_/A sky130_fd_sc_hd__o21ai_4
XFILLER_29_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19745_ _19814_/B _19683_/Y _19764_/B vssd1 vssd1 vccd1 vccd1 _19760_/A sky130_fd_sc_hd__o21ai_1
X_16957_ _16946_/X _16948_/X _16956_/Y vssd1 vssd1 vccd1 vccd1 _16959_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__14672__A1 _13814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11583__A _18663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15908_ _15903_/X _15906_/Y _15907_/Y vssd1 vssd1 vccd1 vccd1 _15978_/A sky130_fd_sc_hd__o21ai_4
X_19676_ _19571_/A _19571_/B _22918_/Q vssd1 vssd1 vccd1 vccd1 _19676_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16888_ _17076_/C _17048_/D vssd1 vssd1 vccd1 vccd1 _16889_/C sky130_fd_sc_hd__nand2_2
XFILLER_92_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18627_ _15538_/X _15541_/X _18636_/A _18626_/Y vssd1 vssd1 vccd1 vccd1 _18627_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15839_ _15839_/A vssd1 vssd1 vccd1 vccd1 _15840_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19141__A_N _22915_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18558_ _18407_/A _18407_/B _18396_/C vssd1 vssd1 vccd1 vccd1 _18559_/B sky130_fd_sc_hd__o21ai_1
XFILLER_80_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17509_ _17500_/Y _17501_/X _17508_/Y vssd1 vssd1 vccd1 vccd1 _17719_/B sky130_fd_sc_hd__o21ai_1
XFILLER_61_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18489_ _12009_/X _18333_/X _18340_/B _18482_/Y _18705_/A vssd1 vssd1 vccd1 vccd1
+ _18490_/C sky130_fd_sc_hd__o221ai_4
XFILLER_61_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17913__A2 _17227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1097 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20520_ _20623_/A _20623_/B _20491_/Y _20501_/A vssd1 vssd1 vccd1 vccd1 _20522_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19197__A _19197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20451_ _16179_/X _20728_/A _20449_/Y _20450_/X vssd1 vssd1 vccd1 vccd1 _20532_/A
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__13022__B _13022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17126__B1 _17125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20382_ _20371_/A _20371_/B _20366_/B _20366_/C vssd1 vssd1 vccd1 vccd1 _20382_/X
+ sky130_fd_sc_hd__a22o_1
X_22121_ _22171_/A _22171_/B _22173_/D vssd1 vssd1 vccd1 vccd1 _22190_/A sky130_fd_sc_hd__nand3b_1
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput120 _22668_/Q vssd1 vssd1 vccd1 vccd1 y[4] sky130_fd_sc_hd__buf_2
XFILLER_133_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17429__A1 _17427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22052_ _22039_/Y _22044_/X _22046_/X vssd1 vssd1 vccd1 vccd1 _22100_/C sky130_fd_sc_hd__a21o_1
XANTENNA__18626__B1 _18810_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21003_ _20905_/B _20959_/A _20905_/A _20959_/B _21002_/Y vssd1 vssd1 vccd1 vccd1
+ _21004_/B sky130_fd_sc_hd__a41oi_4
XFILLER_87_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16101__A1 _12716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16101__B2 _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11493__A _18130_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19051__B1 _15530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22954_ _22959_/CLK _22954_/D vssd1 vssd1 vccd1 vccd1 _22954_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14300__C _14300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21905_ _21801_/A _21721_/A _21721_/B vssd1 vssd1 vccd1 vccd1 _21906_/A sky130_fd_sc_hd__o21bai_1
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22885_ _22922_/CLK input79/X vssd1 vssd1 vccd1 vccd1 _22885_/Q sky130_fd_sc_hd__dfxtp_1
X_21836_ _21836_/A vssd1 vssd1 vccd1 vccd1 _21836_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19354__A1 _17381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18157__A2 _11905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21767_ _21767_/A vssd1 vssd1 vccd1 vccd1 _21767_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14309__A input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ _18339_/C vssd1 vssd1 vccd1 vccd1 _18875_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14718__A2 _15114_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20718_ _20718_/A _20717_/Y vssd1 vssd1 vccd1 vccd1 _20718_/X sky130_fd_sc_hd__or2b_1
XFILLER_169_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21698_ _21695_/C _21698_/B _21698_/C vssd1 vssd1 vccd1 vccd1 _21702_/B sky130_fd_sc_hd__nand3b_2
XANTENNA__12729__A1 _12988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11451_ _18303_/C vssd1 vssd1 vccd1 vccd1 _11454_/A sky130_fd_sc_hd__inv_2
X_20649_ _20650_/A _20650_/B _20650_/C vssd1 vssd1 vccd1 vccd1 _20652_/A sky130_fd_sc_hd__a21o_1
XFILLER_183_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11937__C1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14170_ _14167_/A _14167_/B _14167_/C vssd1 vssd1 vccd1 vccd1 _14170_/X sky130_fd_sc_hd__a21o_1
X_11382_ _11995_/B vssd1 vssd1 vccd1 vccd1 _11772_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11952__A2 _11774_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13121_ _13105_/Y _21750_/C _21362_/A _13120_/Y vssd1 vssd1 vccd1 vccd1 _13122_/C
+ sky130_fd_sc_hd__a31o_1
X_22319_ _22336_/A _22341_/A _22320_/A vssd1 vssd1 vccd1 vccd1 _22323_/A sky130_fd_sc_hd__o21bai_1
XFILLER_139_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13052_ _22724_/Q vssd1 vssd1 vccd1 vccd1 _13158_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input54_A wb_dat_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12003_ _12003_/A _12003_/B _12003_/C vssd1 vssd1 vccd1 vccd1 _12004_/B sky130_fd_sc_hd__and3_1
X_17860_ _17860_/A _17860_/B vssd1 vssd1 vccd1 vccd1 _17861_/B sky130_fd_sc_hd__nand2_1
XFILLER_105_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_868 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18632__A3 _18626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16643__A2 _17039_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16811_ _19012_/C _17108_/B _16810_/C _16810_/D vssd1 vssd1 vccd1 vccd1 _16812_/C
+ sky130_fd_sc_hd__a22o_1
X_17791_ _17790_/Y _18044_/A _17788_/X vssd1 vssd1 vccd1 vccd1 _17793_/C sky130_fd_sc_hd__a21oi_1
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19530_ _19530_/A _19530_/B _19530_/C _19530_/D vssd1 vssd1 vccd1 vccd1 _19530_/X
+ sky130_fd_sc_hd__and4_1
X_16742_ _16743_/A _16743_/C _16743_/B vssd1 vssd1 vccd1 vccd1 _16742_/Y sky130_fd_sc_hd__a21oi_4
X_13954_ _13954_/A _13954_/B _14613_/A _14203_/B vssd1 vssd1 vccd1 vccd1 _14026_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_98_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19593__A1 _17730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12905_ _20133_/B vssd1 vssd1 vccd1 vccd1 _16078_/B sky130_fd_sc_hd__buf_2
X_16673_ _16673_/A vssd1 vssd1 vccd1 vccd1 _16673_/Y sky130_fd_sc_hd__inv_2
X_19461_ _19461_/A _19461_/B _19461_/C vssd1 vssd1 vccd1 vccd1 _19461_/X sky130_fd_sc_hd__and3_1
XFILLER_47_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13885_ _13881_/Y _13883_/Y _13884_/X vssd1 vssd1 vccd1 vccd1 _13920_/B sky130_fd_sc_hd__o21ai_1
XFILLER_59_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18412_ _18401_/X _18403_/X _18394_/Y _18399_/Y vssd1 vssd1 vccd1 vccd1 _18415_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_59_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15624_ _15624_/A _20593_/B _20678_/B _16563_/C vssd1 vssd1 vccd1 vccd1 _16431_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12836_ _12820_/Y _12832_/Y _16708_/A _12718_/A vssd1 vssd1 vccd1 vccd1 _12838_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _19458_/A _19392_/B vssd1 vssd1 vccd1 vccd1 _19398_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_768 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19345__A1 _11598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22955__CLK _22959_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19345__B2 _11474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_943 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15555_ _16253_/B _15543_/Y _15547_/X _15554_/X vssd1 vssd1 vccd1 vccd1 _15583_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_18343_ _18484_/A vssd1 vssd1 vccd1 vccd1 _18343_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16159__A1 _16157_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12767_/A vssd1 vssd1 vccd1 vccd1 _20177_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_431 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14219__A _15004_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14510_/C _14506_/B _14506_/C vssd1 vssd1 vccd1 vccd1 _14506_/Y sky130_fd_sc_hd__nand3_1
XFILLER_188_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18274_ _18772_/A _18772_/B _18772_/D vssd1 vssd1 vccd1 vccd1 _18274_/Y sky130_fd_sc_hd__nand3_2
X_11718_ _11718_/A vssd1 vssd1 vccd1 vccd1 _12046_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11640__A1 _11504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15486_ _15486_/A _15486_/B _15486_/C vssd1 vssd1 vccd1 vccd1 _16226_/A sky130_fd_sc_hd__nand3_2
XANTENNA__11640__B2 _11625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15906__A1 _15904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12698_ _12696_/X _13022_/C _12605_/Y _12592_/Y vssd1 vssd1 vccd1 vccd1 _12737_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_175_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17225_ _17225_/A _17225_/B vssd1 vssd1 vccd1 vccd1 _22956_/D sky130_fd_sc_hd__xnor2_1
X_14437_ _22965_/Q vssd1 vssd1 vccd1 vccd1 _16241_/D sky130_fd_sc_hd__clkinv_2
Xinput11 wb_adr_i[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11649_ _11644_/X _11646_/Y _11689_/A _11648_/Y vssd1 vssd1 vccd1 vccd1 _11649_/Y
+ sky130_fd_sc_hd__o211ai_1
Xinput22 wb_adr_i[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_1
Xinput33 wb_clk_i vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_6
XFILLER_190_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17156_ _17168_/B vssd1 vssd1 vccd1 vccd1 _17180_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput44 wb_dat_i[18] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14368_ _22700_/Q _14344_/X _14351_/X _21307_/B _14367_/X vssd1 vssd1 vccd1 vccd1
+ _14368_/X sky130_fd_sc_hd__a221o_1
Xinput55 wb_dat_i[28] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput66 wb_dat_i[9] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_4
Xinput77 x[6] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__16153__B _17006_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16107_ _16106_/C _12681_/A _12681_/B _19000_/A _16067_/D vssd1 vssd1 vccd1 vccd1
+ _16107_/X sky130_fd_sc_hd__a32o_1
X_13319_ _13319_/A vssd1 vssd1 vccd1 vccd1 _13319_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11578__A _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17087_ _17087_/A _17087_/B vssd1 vssd1 vccd1 vccd1 _17087_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14299_ input7/X input6/X input28/X input27/X vssd1 vssd1 vccd1 vccd1 _14300_/D sky130_fd_sc_hd__or4_1
XFILLER_171_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16038_ _16038_/A _16038_/B _16038_/C vssd1 vssd1 vccd1 vccd1 _16421_/C sky130_fd_sc_hd__nand3_4
XFILLER_192_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20966__A1 _17423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_bq_clk_i clkbuf_4_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _22850_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_97_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17989_ _17989_/A _17991_/A _17989_/C vssd1 vssd1 vccd1 vccd1 _18062_/D sky130_fd_sc_hd__nand3_1
XFILLER_96_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19728_ _19735_/B _19735_/C _19735_/A vssd1 vssd1 vccd1 vccd1 _19728_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__19480__A _19480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12202__A _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19584__B2 _11639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19659_ _19561_/A _19564_/Y _19577_/A vssd1 vssd1 vccd1 vccd1 _19659_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16398__A1 _16400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22670_ _22968_/CLK _22670_/D vssd1 vssd1 vccd1 vccd1 _22670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17431__C _17431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21621_ _21725_/A _21725_/B _21621_/C vssd1 vssd1 vccd1 vccd1 _21766_/B sky130_fd_sc_hd__and3_1
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14129__A _14191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21552_ _21406_/A _21406_/B _21406_/C _21416_/A vssd1 vssd1 vccd1 vccd1 _21553_/D
+ sky130_fd_sc_hd__a31o_2
XFILLER_178_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20503_ _20359_/A _20514_/A _20359_/C _20326_/Y vssd1 vssd1 vccd1 vccd1 _20503_/Y
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__13908__B1 _22761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20792__C _20792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21483_ _13050_/X _21192_/A _21478_/X _21486_/A _21482_/Y vssd1 vssd1 vccd1 vccd1
+ _21504_/C sky130_fd_sc_hd__o221ai_4
XFILLER_165_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19358__C _19358_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18847__B1 _19014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20434_ _20553_/A _20553_/B _20309_/A vssd1 vssd1 vccd1 vccd1 _20434_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_180_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20365_ _20224_/A _20224_/B _20224_/C _20364_/Y _20211_/Y vssd1 vssd1 vccd1 vccd1
+ _20365_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_164_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22104_ _22122_/C _22223_/A vssd1 vssd1 vccd1 vccd1 _22119_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14333__B1 _14313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20296_ _20319_/B _20319_/A _20295_/Y _20181_/A vssd1 vssd1 vccd1 vccd1 _20296_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22035_ _22131_/B vssd1 vssd1 vccd1 vccd1 _22196_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22231__D _22231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__B _11935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22937_ _22937_/CLK _22937_/D vssd1 vssd1 vccd1 vccd1 _22937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15423__A _18716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13670_ _13660_/X _13665_/Y _13669_/Y vssd1 vssd1 vccd1 vccd1 _13671_/B sky130_fd_sc_hd__o21ai_1
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17341__C _17341_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22868_ _22916_/CLK _22868_/D vssd1 vssd1 vccd1 vccd1 _22868_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_188_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_256 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19327__B2 _18856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12621_ _12621_/A _12621_/B vssd1 vssd1 vccd1 vccd1 _12621_/Y sky130_fd_sc_hd__nand2_1
XFILLER_188_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21819_ _21816_/Y _21817_/Y _21818_/Y vssd1 vssd1 vccd1 vccd1 _21834_/D sky130_fd_sc_hd__o21ai_2
X_22799_ _22799_/CLK _22799_/D vssd1 vssd1 vccd1 vccd1 _22799_/Q sky130_fd_sc_hd__dfxtp_2
X_15340_ _15797_/A vssd1 vssd1 vccd1 vccd1 _15891_/A sky130_fd_sc_hd__clkbuf_4
X_12552_ _12565_/A _12567_/A vssd1 vssd1 vccd1 vccd1 _12790_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18453__B _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ _11503_/A vssd1 vssd1 vccd1 vccd1 _11503_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15271_ _22878_/Q _15271_/B _15279_/A vssd1 vssd1 vccd1 vccd1 _15273_/A sky130_fd_sc_hd__nand3b_1
XFILLER_184_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12782__A _16488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12483_ _12487_/B vssd1 vssd1 vccd1 vccd1 _12792_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_184_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17010_ _16828_/B _16836_/X _16990_/Y vssd1 vssd1 vccd1 vccd1 _17010_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14222_ _14222_/A _14494_/C vssd1 vssd1 vccd1 vccd1 _14222_/Y sky130_fd_sc_hd__nand2_1
X_11434_ _11434_/A vssd1 vssd1 vccd1 vccd1 _14429_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__14572__B1 _14362_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11398__A _18876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20207__C _20207_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153_ _14153_/A _14285_/C vssd1 vssd1 vccd1 vccd1 _14248_/C sky130_fd_sc_hd__nor2_1
X_11365_ _18116_/A _11430_/B _12003_/B vssd1 vssd1 vccd1 vccd1 _11366_/A sky130_fd_sc_hd__o21ai_2
XFILLER_180_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13104_ _13330_/A _21595_/B _21448_/C vssd1 vssd1 vccd1 vccd1 _13105_/B sky130_fd_sc_hd__nand3_1
XFILLER_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14324__B1 _14313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18961_ _19279_/A _19279_/B _19281_/A vssd1 vssd1 vccd1 vccd1 _18965_/A sky130_fd_sc_hd__nand3_1
XANTENNA__16864__A2 _16753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14084_ _14161_/B _14149_/B _14161_/C vssd1 vssd1 vccd1 vccd1 _14147_/D sky130_fd_sc_hd__nand3_1
X_11296_ _11968_/B vssd1 vssd1 vccd1 vccd1 _18691_/C sky130_fd_sc_hd__buf_2
XANTENNA__22398__A0 _22700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12006__B _12006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ _17959_/A _17959_/B vssd1 vssd1 vccd1 vccd1 _17914_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _13037_/B _13035_/B vssd1 vssd1 vccd1 vccd1 _13036_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18892_ _19587_/D vssd1 vssd1 vccd1 vccd1 _19771_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_105_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_676 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17843_ _17843_/A _17904_/A vssd1 vssd1 vccd1 vccd1 _17869_/A sky130_fd_sc_hd__xor2_4
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17235__D _20870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19015__B1 _15690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17774_ _17777_/C _17776_/A _17785_/B vssd1 vssd1 vccd1 vccd1 _17778_/A sky130_fd_sc_hd__a21boi_2
XANTENNA__13835__C1 _14112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14986_ _15039_/A _15047_/B _14985_/X vssd1 vssd1 vccd1 vccd1 _15046_/B sky130_fd_sc_hd__o21ba_2
XFILLER_19_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19513_ _19521_/A _19581_/A _19521_/D vssd1 vssd1 vccd1 vccd1 _19513_/Y sky130_fd_sc_hd__nand3_1
X_16725_ _16312_/X _16714_/X _16720_/Y vssd1 vssd1 vccd1 vccd1 _16725_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__17532__B _17532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13937_ _13937_/A _13937_/B _13937_/C _13937_/D vssd1 vssd1 vccd1 vccd1 _13957_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_170_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19444_ _19681_/A _19681_/C _19680_/A vssd1 vssd1 vccd1 vccd1 _19447_/A sky130_fd_sc_hd__a21oi_1
XFILLER_34_234 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16656_ _16206_/A _15879_/A _16432_/Y _16433_/Y _16210_/Y vssd1 vssd1 vccd1 vccd1
+ _16657_/A sky130_fd_sc_hd__o2111a_1
X_13868_ _13861_/Y _13862_/X _14169_/A vssd1 vssd1 vccd1 vccd1 _13868_/X sky130_fd_sc_hd__o21a_1
XFILLER_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15052__A1 _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15607_ _16323_/A _16323_/B _16323_/C _16319_/B vssd1 vssd1 vccd1 vccd1 _15608_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ _12852_/B vssd1 vssd1 vccd1 vccd1 _12859_/A sky130_fd_sc_hd__clkbuf_2
X_19375_ _19356_/X _19363_/Y _19369_/Y _19379_/B vssd1 vssd1 vccd1 vccd1 _19376_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_50_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16587_ _16599_/C _16599_/B _16578_/X _16586_/X vssd1 vssd1 vccd1 vccd1 _16594_/A
+ sky130_fd_sc_hd__o2bb2ai_4
X_13799_ _22758_/Q vssd1 vssd1 vccd1 vccd1 _13799_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_163_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18326_ _11904_/X _11905_/X _19496_/B _15415_/C _19496_/C vssd1 vssd1 vccd1 vccd1
+ _18326_/Y sky130_fd_sc_hd__o2111ai_4
X_15538_ _15548_/A vssd1 vssd1 vccd1 vccd1 _15538_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18257_ _18257_/A _18257_/B _18257_/C vssd1 vssd1 vccd1 vccd1 _18257_/Y sky130_fd_sc_hd__nand3_1
X_15469_ _11568_/A _11568_/B _12606_/X _12607_/X vssd1 vssd1 vccd1 vccd1 _15470_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12692__A _20471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17208_ _17208_/A _17208_/B _17208_/C vssd1 vssd1 vccd1 vccd1 _17513_/C sky130_fd_sc_hd__nand3_1
XFILLER_163_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18188_ _12189_/Y _12186_/Y _12182_/C vssd1 vssd1 vccd1 vccd1 _18188_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_144_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20636__B1 _20631_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17139_ _17139_/A vssd1 vssd1 vccd1 vccd1 _17532_/C sky130_fd_sc_hd__buf_2
XFILLER_144_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17501__B1 _22898_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18844__A3 _19587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18810__C _19507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20150_ _20150_/A _20150_/B _20150_/C vssd1 vssd1 vccd1 vccd1 _20167_/B sky130_fd_sc_hd__nand3_2
XFILLER_143_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19194__B _19490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22389__A0 _12343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20081_ _20728_/A _13022_/D _20077_/B _20293_/A vssd1 vssd1 vccd1 vccd1 _20161_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16068__B1 _16098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20133__B _20133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16607__A2 _16377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11755__B _19461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12629__B1 _12630_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19557__A1 _12064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20983_ _20933_/Y _20935_/Y _20938_/Y vssd1 vssd1 vccd1 vccd1 _20985_/A sky130_fd_sc_hd__a21bo_1
XFILLER_26_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22722_ input33/X _22722_/D vssd1 vssd1 vccd1 vccd1 _22722_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11852__A1 _11566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15043__A1 _14845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16058__B _19000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22653_ _22653_/A vssd1 vssd1 vccd1 vccd1 _22813_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16791__A1 _16778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21604_ _21604_/A _21604_/B _21604_/C vssd1 vssd1 vccd1 vccd1 _21645_/B sky130_fd_sc_hd__nand3_1
XFILLER_178_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22584_ _22783_/Q input59/X _22584_/S vssd1 vssd1 vccd1 vccd1 _22585_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13698__A _22871_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21535_ _21535_/A _21535_/B _21535_/C vssd1 vssd1 vccd1 vccd1 _21535_/X sky130_fd_sc_hd__and3_1
XFILLER_167_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21466_ _21466_/A _21466_/B vssd1 vssd1 vccd1 vccd1 _21466_/X sky130_fd_sc_hd__or2_1
XFILLER_153_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14306__B input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20417_ _20844_/A _15890_/X _20155_/B _20144_/Y _20155_/C vssd1 vssd1 vccd1 vccd1
+ _20429_/C sky130_fd_sc_hd__o221a_2
XFILLER_162_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19493__B1 _19490_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21397_ _21442_/A _21445_/C _21445_/A vssd1 vssd1 vccd1 vccd1 _21399_/B sky130_fd_sc_hd__a21o_1
XFILLER_175_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12580__A2 _12577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20348_ _20340_/Y _20343_/Y _20344_/Y _20347_/Y vssd1 vssd1 vccd1 vccd1 _20349_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_108_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15418__A _20355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_1099 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20279_ _12525_/A _12525_/B _20177_/A vssd1 vssd1 vccd1 vccd1 _20281_/A sky130_fd_sc_hd__a21o_1
XFILLER_103_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22018_ _22016_/A _22017_/X _22679_/Q vssd1 vssd1 vccd1 vccd1 _22018_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14041__B _22863_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14840_ _14758_/C _14660_/B _14759_/Y _14757_/B vssd1 vssd1 vccd1 vccd1 _14840_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12096__A1 _11705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input17_A wb_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771_ _14771_/A vssd1 vssd1 vccd1 vccd1 _15107_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11983_ _11793_/B _11974_/Y _12137_/A vssd1 vssd1 vccd1 vccd1 _11984_/A sky130_fd_sc_hd__o21ai_1
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13832__A2 _13746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16510_ _16489_/X _16509_/Y _15542_/X _16494_/X vssd1 vssd1 vccd1 vccd1 _16510_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_13722_ _22869_/Q vssd1 vssd1 vccd1 vccd1 _14110_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_543 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17490_ _17490_/A _17490_/B _17490_/C vssd1 vssd1 vccd1 vccd1 _17491_/B sky130_fd_sc_hd__nand3_1
XANTENNA__16767__D1 _19687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16441_ _16433_/C _16439_/Y _16440_/Y vssd1 vssd1 vccd1 vccd1 _16441_/X sky130_fd_sc_hd__o21a_1
X_13653_ _21489_/A _13572_/B _13657_/A _13657_/B vssd1 vssd1 vccd1 vccd1 _13655_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18464__A _18464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _12785_/B vssd1 vssd1 vccd1 vccd1 _12938_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_176_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16372_ _15601_/Y _15602_/X _15644_/Y _15654_/Y vssd1 vssd1 vccd1 vccd1 _16372_/X
+ sky130_fd_sc_hd__o211a_1
X_19160_ _19160_/A vssd1 vssd1 vccd1 vccd1 _19517_/A sky130_fd_sc_hd__clkbuf_4
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13584_ _21595_/B vssd1 vssd1 vccd1 vccd1 _21195_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_169_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _19046_/C _18849_/D _12098_/Y _18110_/X vssd1 vssd1 vccd1 vccd1 _18278_/B
+ sky130_fd_sc_hd__a31o_2
X_15323_ _17532_/B _18690_/B _17532_/A vssd1 vssd1 vccd1 vccd1 _15324_/A sky130_fd_sc_hd__and3_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _22824_/Q vssd1 vssd1 vccd1 vccd1 _20128_/A sky130_fd_sc_hd__buf_2
XFILLER_33_70 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19091_ _19091_/A _19091_/B _19091_/C vssd1 vssd1 vccd1 vccd1 _19091_/X sky130_fd_sc_hd__or3_1
XFILLER_184_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18042_ _18042_/A vssd1 vssd1 vccd1 vccd1 _18042_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15254_ _15240_/A _15224_/A _15238_/B _15238_/A vssd1 vssd1 vccd1 vccd1 _15266_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12466_ _12802_/A _12813_/A _12579_/C vssd1 vssd1 vccd1 vccd1 _20210_/A sky130_fd_sc_hd__nand3_4
XFILLER_184_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14205_ _14868_/C _14203_/B _14157_/A _14861_/C vssd1 vssd1 vccd1 vccd1 _14205_/Y
+ sky130_fd_sc_hd__a22oi_1
X_11417_ _22789_/Q vssd1 vssd1 vccd1 vccd1 _11418_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17808__A _17833_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15185_ _15213_/A _15185_/B _15160_/A vssd1 vssd1 vccd1 vccd1 _15186_/C sky130_fd_sc_hd__or3b_1
X_12397_ _12586_/A vssd1 vssd1 vccd1 vccd1 _15466_/C sky130_fd_sc_hd__buf_2
XANTENNA__16712__A _20471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21291__B1 _22673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14136_ _14134_/Y _14135_/X _14111_/X vssd1 vssd1 vccd1 vccd1 _14231_/C sky130_fd_sc_hd__o21ai_1
X_11348_ _22788_/Q vssd1 vssd1 vccd1 vccd1 _18115_/C sky130_fd_sc_hd__clkbuf_2
X_19993_ _20037_/C _19992_/C _19992_/B vssd1 vssd1 vccd1 vccd1 _19994_/B sky130_fd_sc_hd__o21ai_1
XFILLER_181_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20234__A _20234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16431__B _16431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11856__A _15991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18944_ _18763_/A _18764_/B _18754_/X vssd1 vssd1 vccd1 vccd1 _18945_/C sky130_fd_sc_hd__a21boi_2
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14067_ _14564_/C vssd1 vssd1 vccd1 vccd1 _14868_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11279_ _22799_/Q vssd1 vssd1 vccd1 vccd1 _11496_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17246__C _17532_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_602 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13018_ _12579_/X _13016_/X _13017_/X _12989_/B vssd1 vssd1 vccd1 vccd1 _13018_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11575__B _11899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18875_ _18876_/A _18876_/B _18875_/C _18875_/D vssd1 vssd1 vccd1 vccd1 _18875_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_121_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_646 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17826_ _17826_/A _17826_/B _17826_/C vssd1 vssd1 vccd1 vccd1 _17827_/C sky130_fd_sc_hd__nand3_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19461__C _19461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17757_ _17753_/A _17753_/B _17755_/Y _17756_/Y vssd1 vssd1 vccd1 vccd1 _17760_/C
+ sky130_fd_sc_hd__o22ai_2
XFILLER_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16578__A2_N _16879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22543__A0 _14366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14969_ _14969_/A _14969_/B vssd1 vssd1 vccd1 vccd1 _14971_/B sky130_fd_sc_hd__xor2_1
X_16708_ _16708_/A vssd1 vssd1 vccd1 vccd1 _16708_/X sky130_fd_sc_hd__clkbuf_4
X_17688_ _17688_/A _17688_/B _17688_/C vssd1 vssd1 vccd1 vccd1 _17690_/A sky130_fd_sc_hd__nand3_1
X_19427_ _19434_/A _19427_/B _19427_/C _19427_/D vssd1 vssd1 vccd1 vccd1 _19561_/A
+ sky130_fd_sc_hd__nand4_2
X_16639_ _16378_/X _16636_/Y _16637_/Y _16638_/Y vssd1 vssd1 vccd1 vccd1 _16895_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13587__A1 _21445_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19358_ _19358_/A _19358_/B _19358_/C _19358_/D vssd1 vssd1 vccd1 vccd1 _19359_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_188_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18093__B _18093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18514__A2 _11988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18309_ _18309_/A _18309_/B _18442_/B vssd1 vssd1 vccd1 vccd1 _18309_/X sky130_fd_sc_hd__and3_1
XANTENNA__15328__A2 _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19289_ _19289_/A _19288_/Y vssd1 vssd1 vccd1 vccd1 _19290_/C sky130_fd_sc_hd__or2b_1
XFILLER_175_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22673__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21320_ _21320_/A _21320_/B _21320_/C vssd1 vssd1 vccd1 vccd1 _21321_/A sky130_fd_sc_hd__nand3_2
XFILLER_163_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20609__B1 _20241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12011__A1 _12009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21251_ _21251_/A _21251_/B _21251_/C vssd1 vssd1 vccd1 vccd1 _21251_/X sky130_fd_sc_hd__and3_1
XFILLER_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20085__A1 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20202_ _20115_/A _20115_/B _20115_/C vssd1 vssd1 vccd1 vccd1 _20202_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21182_ _21245_/A _21245_/B vssd1 vssd1 vccd1 vccd1 _21240_/A sky130_fd_sc_hd__xnor2_1
XFILLER_143_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16341__B _16617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11766__A _22792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20133_ _20133_/A _20133_/B _20323_/D vssd1 vssd1 vccd1 vccd1 _20133_/Y sky130_fd_sc_hd__nand3_2
XFILLER_98_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20064_ _12894_/A _12894_/B _13011_/A vssd1 vssd1 vccd1 vccd1 _20064_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A wb_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22534__A0 _13896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16069__A _19470_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11932__C _11932_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20966_ _17423_/X _17424_/X _21082_/B vssd1 vssd1 vccd1 vccd1 _20966_/X sky130_fd_sc_hd__a21o_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22705_ _22801_/CLK _22705_/D vssd1 vssd1 vccd1 vccd1 _22705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16764__A1 _15546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _20897_/A _20897_/B vssd1 vssd1 vccd1 vccd1 _20961_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15701__A _20678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22636_ _22636_/A vssd1 vssd1 vccd1 vccd1 _22805_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__21422__B _21422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15972__C1 _15901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16516__A1 _18203_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22567_ _22775_/Q input50/X _22569_/S vssd1 vssd1 vccd1 vccd1 _22568_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12320_ _12320_/A _12369_/A vssd1 vssd1 vccd1 vccd1 _12320_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21518_ _13373_/A _13373_/B _21689_/A vssd1 vssd1 vccd1 vccd1 _21539_/A sky130_fd_sc_hd__a21o_1
XFILLER_142_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22498_ _22498_/A vssd1 vssd1 vccd1 vccd1 _22744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ _12251_/A _12251_/B _12251_/C vssd1 vssd1 vccd1 vccd1 _18261_/A sky130_fd_sc_hd__nand3_1
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19466__B1 _11672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21449_ _21449_/A _21449_/B vssd1 vssd1 vccd1 vccd1 _21449_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17477__C1 _17466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ _12189_/A _18208_/B _12182_/C _12182_/D vssd1 vssd1 vccd1 vccd1 _12188_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_134_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11761__B1 _11932_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16990_ _16822_/B _16822_/C _16822_/A vssd1 vssd1 vccd1 vccd1 _16990_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15941_ _15941_/A vssd1 vssd1 vccd1 vccd1 _15941_/X sky130_fd_sc_hd__buf_4
XFILLER_95_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18459__A _18459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18660_ _19199_/A _19320_/A _18865_/A _18659_/B vssd1 vssd1 vccd1 vccd1 _18661_/C
+ sky130_fd_sc_hd__a22o_1
X_15872_ _15952_/A _15952_/B _15952_/C _16034_/C vssd1 vssd1 vccd1 vccd1 _15951_/A
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__15255__A1 _14990_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12003__C _12003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17611_ _17611_/A _17611_/B vssd1 vssd1 vccd1 vccd1 _17611_/X sky130_fd_sc_hd__and2_1
XANTENNA__18992__A2 _18984_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14823_ _14738_/B _14737_/B _14737_/A vssd1 vssd1 vccd1 vccd1 _14825_/A sky130_fd_sc_hd__a21bo_1
X_18591_ _18773_/A _18774_/A _18274_/Y _18772_/C vssd1 vssd1 vccd1 vccd1 _18591_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__22525__A0 _13826_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _20870_/A _20870_/B _19768_/C _17539_/Y _17535_/Y vssd1 vssd1 vccd1 vccd1
+ _17544_/B sky130_fd_sc_hd__a32o_1
X_11966_ _11945_/A _11777_/Y _11951_/Y vssd1 vssd1 vccd1 vccd1 _11966_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20536__C1 _20263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14754_ _14655_/A _14655_/B _14752_/B vssd1 vssd1 vccd1 vccd1 _14756_/B sky130_fd_sc_hd__o21ai_2
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15007__A1 _14818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ _13776_/B _13849_/C _13776_/A vssd1 vssd1 vccd1 vccd1 _14258_/B sky130_fd_sc_hd__a21oi_1
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17473_ _17486_/A _17473_/B vssd1 vssd1 vccd1 vccd1 _17474_/C sky130_fd_sc_hd__nand2_1
XANTENNA__11292__A2 _22953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16129__D _16192_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14685_ _14685_/A _14685_/B vssd1 vssd1 vccd1 vccd1 _14685_/Y sky130_fd_sc_hd__nand2_1
X_11897_ _11909_/A _11909_/B _11909_/C vssd1 vssd1 vccd1 vccd1 _11897_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__16755__B2 _16740_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19212_ _19507_/A _19587_/C _19687_/D _19587_/A vssd1 vssd1 vccd1 vccd1 _19218_/B
+ sky130_fd_sc_hd__nand4_2
X_16424_ _16424_/A _16424_/B _16424_/C vssd1 vssd1 vccd1 vccd1 _16424_/Y sky130_fd_sc_hd__nand3_1
X_13636_ _13657_/C _13634_/X _13657_/A vssd1 vssd1 vccd1 vccd1 _13666_/C sky130_fd_sc_hd__o21ai_1
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19143_ _18788_/A _18969_/X _18968_/A _18970_/Y vssd1 vssd1 vccd1 vccd1 _19143_/Y
+ sky130_fd_sc_hd__o211ai_2
X_16355_ _16355_/A _16355_/B _16355_/C vssd1 vssd1 vccd1 vccd1 _16627_/A sky130_fd_sc_hd__nand3_4
XFILLER_13_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13567_ _13527_/Y _13530_/X _13524_/X vssd1 vssd1 vccd1 vccd1 _13567_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14227__A _15114_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15306_ _16256_/A _16256_/B _15306_/C _15776_/D vssd1 vssd1 vccd1 vccd1 _15306_/Y
+ sky130_fd_sc_hd__nand4_4
X_12518_ _12518_/A vssd1 vssd1 vccd1 vccd1 _12549_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19074_ _19074_/A _19074_/B _19074_/C _19074_/D vssd1 vssd1 vccd1 vccd1 _19148_/C
+ sky130_fd_sc_hd__nand4_1
X_16286_ _16286_/A vssd1 vssd1 vccd1 vccd1 _16286_/Y sky130_fd_sc_hd__inv_2
X_13498_ _13498_/A _13498_/B _13498_/C vssd1 vssd1 vccd1 vccd1 _21280_/A sky130_fd_sc_hd__nand3_1
XFILLER_172_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22444__A _22512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18025_ _21048_/B _18023_/X _21048_/C _18778_/D _21081_/B vssd1 vssd1 vccd1 vccd1
+ _18025_/X sky130_fd_sc_hd__o32a_1
XANTENNA__17538__A _19507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15237_ _15238_/A _15212_/A _15238_/B vssd1 vssd1 vccd1 vccd1 _15240_/D sky130_fd_sc_hd__o21a_1
X_12449_ _16465_/A _12411_/A _20255_/C _12307_/Y vssd1 vssd1 vccd1 vccd1 _12449_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_172_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15168_ _15168_/A _15181_/A _15168_/C vssd1 vssd1 vccd1 vccd1 _15181_/B sky130_fd_sc_hd__nor3_2
XFILLER_158_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11752__B1 _11751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11897__B1_N _11909_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _14203_/A _14564_/C vssd1 vssd1 vccd1 vccd1 _14119_/Y sky130_fd_sc_hd__nand2_1
X_19976_ _19976_/A _19976_/B _19976_/C vssd1 vssd1 vccd1 vccd1 _19976_/Y sky130_fd_sc_hd__nand3_1
X_15099_ _15098_/A _15098_/B _15098_/C vssd1 vssd1 vccd1 vccd1 _15100_/B sky130_fd_sc_hd__a21o_1
XFILLER_68_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15494__A1 _17379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18927_ _18938_/A _18937_/A _18938_/B vssd1 vssd1 vccd1 vccd1 _18927_/Y sky130_fd_sc_hd__nand3_2
XFILLER_140_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18858_ _18858_/A vssd1 vssd1 vccd1 vccd1 _19481_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17809_ _19901_/A _21017_/A _21017_/B _20972_/B _19901_/D vssd1 vssd1 vccd1 vccd1
+ _17811_/D sky130_fd_sc_hd__a32o_1
XFILLER_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18789_ _18970_/B _18789_/B vssd1 vssd1 vccd1 vccd1 _18792_/A sky130_fd_sc_hd__nand2_1
XANTENNA__21319__A1 _13662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20790__A2 _16580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20820_ _20748_/A _20748_/C _20748_/B vssd1 vssd1 vccd1 vccd1 _20822_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__18196__B1 _11634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20751_ _20751_/A _20751_/B _20751_/C vssd1 vssd1 vccd1 vccd1 _20758_/B sky130_fd_sc_hd__nor3_1
XFILLER_165_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16617__A _16617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20682_ _20682_/A _20682_/B _20682_/C vssd1 vssd1 vccd1 vccd1 _20683_/B sky130_fd_sc_hd__nand3_2
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22421_ _22421_/A vssd1 vssd1 vccd1 vccd1 _22710_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12232__A1 _22658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14509__B1 _14503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13041__A _13045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22352_ _22352_/A _22352_/B vssd1 vssd1 vccd1 vccd1 _22354_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12783__A2 _15455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21303_ _22730_/Q _22731_/Q vssd1 vssd1 vccd1 vccd1 _21304_/D sky130_fd_sc_hd__nor2_1
XANTENNA__11991__B1 _12107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22283_ _22300_/B _22284_/C _22300_/A vssd1 vssd1 vccd1 vccd1 _22285_/A sky130_fd_sc_hd__a21oi_1
XFILLER_85_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1022 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21234_ _21234_/A _21233_/Y vssd1 vssd1 vccd1 vccd1 _21234_/X sky130_fd_sc_hd__or2b_1
XFILLER_132_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11496__A _22790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21165_ _21165_/A _22947_/Q vssd1 vssd1 vccd1 vccd1 _21165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20116_ _20116_/A vssd1 vssd1 vccd1 vccd1 _20154_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21096_ _21061_/A _21061_/B _21094_/Y _21095_/Y vssd1 vssd1 vccd1 vccd1 _21115_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__18279__A _18279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20047_ _22927_/Q _20059_/A _20059_/B vssd1 vssd1 vccd1 vccd1 _20049_/B sky130_fd_sc_hd__or3_1
XFILLER_19_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15415__B _20675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1111 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11820_/A vssd1 vssd1 vccd1 vccd1 _16014_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21998_ _21987_/Y _21989_/Y _22075_/B _21994_/A _22029_/A vssd1 vssd1 vccd1 vccd1
+ _21998_/X sky130_fd_sc_hd__o2111a_1
XFILLER_61_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_bq_clk_i clkbuf_3_7_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _22951_/CLK
+ sky130_fd_sc_hd__clkbuf_8
X_11751_ _17421_/A _17422_/A _11454_/A vssd1 vssd1 vccd1 vccd1 _11751_/X sky130_fd_sc_hd__a21o_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20949_ _20949_/A _20949_/B _20949_/C vssd1 vssd1 vccd1 vccd1 _20952_/A sky130_fd_sc_hd__or3_1
XFILLER_18_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15431__A _15707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18445__C _18445_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14470_ _14274_/A _14562_/A _13986_/A vssd1 vssd1 vccd1 vccd1 _14470_/X sky130_fd_sc_hd__o21a_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _14438_/A _15297_/A _11734_/A vssd1 vssd1 vccd1 vccd1 _11702_/A sky130_fd_sc_hd__o21ai_2
XFILLER_144_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16246__B _19197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13421_ _13421_/A vssd1 vssd1 vccd1 vccd1 _22041_/B sky130_fd_sc_hd__clkbuf_4
X_22619_ _22798_/Q input40/X _22619_/S vssd1 vssd1 vccd1 vccd1 _22620_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19838__A _19838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16140_ _16143_/B _16143_/C vssd1 vssd1 vccd1 vccd1 _16140_/Y sky130_fd_sc_hd__nand2_1
X_13352_ _13349_/X _13351_/Y _13315_/X _13354_/B vssd1 vssd1 vccd1 vccd1 _13352_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_128_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12303_ _12303_/A vssd1 vssd1 vccd1 vccd1 _16328_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_182_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16071_ _16056_/Y _16064_/Y _16070_/Y vssd1 vssd1 vccd1 vccd1 _16126_/C sky130_fd_sc_hd__a21oi_2
XFILLER_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13283_ _13269_/X _13276_/X _13413_/B _13282_/Y vssd1 vssd1 vccd1 vccd1 _13481_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__15712__A2 _12727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15022_ _14954_/X _14955_/Y _14952_/Y vssd1 vssd1 vccd1 vccd1 _15023_/B sky130_fd_sc_hd__a21boi_1
XFILLER_170_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12234_ _15530_/A vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12526__A2 _12540_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19830_ _19827_/Y _19757_/Y _19890_/A _19890_/B _19891_/D vssd1 vssd1 vccd1 vccd1
+ _19887_/B sky130_fd_sc_hd__o2111ai_2
XANTENNA__17465__A2 _17728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ _12165_/A vssd1 vssd1 vccd1 vccd1 _15887_/A sky130_fd_sc_hd__buf_2
XFILLER_146_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11931__A2_N _11736_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19761_ _19761_/A _19761_/B _19880_/B _19761_/D vssd1 vssd1 vccd1 vccd1 _19761_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_110_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16973_ _16961_/Y _16966_/X _16970_/Y _16972_/Y vssd1 vssd1 vccd1 vccd1 _17188_/A
+ sky130_fd_sc_hd__o211ai_4
X_12096_ _11705_/X _11737_/A _11707_/A _11936_/A _11583_/B vssd1 vssd1 vccd1 vccd1
+ _12096_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_7_1011 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18712_ _18905_/A _18905_/B _18722_/C _18722_/D vssd1 vssd1 vccd1 vccd1 _18836_/A
+ sky130_fd_sc_hd__nand4_2
X_15924_ _15924_/A _15924_/B _15924_/C vssd1 vssd1 vccd1 vccd1 _16010_/B sky130_fd_sc_hd__nand3_2
X_19692_ _17380_/X _17381_/X _19461_/B _19461_/C _18197_/C vssd1 vssd1 vccd1 vccd1
+ _19692_/Y sky130_fd_sc_hd__o2111ai_1
XANTENNA__12695__D1 _16937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20757__C1 _20759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 wb_adr_i[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
X_18643_ _18933_/A _18933_/B _18933_/C vssd1 vssd1 vccd1 vccd1 _18646_/B sky130_fd_sc_hd__nand3_1
XFILLER_49_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _15855_/A _15855_/B _15944_/C _15855_/D vssd1 vssd1 vccd1 vccd1 _15875_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17821__A _19896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14806_ _14806_/A _14806_/B _14806_/C vssd1 vssd1 vccd1 vccd1 _14902_/A sky130_fd_sc_hd__nand3_1
X_18574_ _18572_/C _18572_/A _18572_/B _18571_/X vssd1 vssd1 vccd1 vccd1 _18574_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__20509__C1 _20913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ _15911_/A vssd1 vssd1 vccd1 vccd1 _17133_/A sky130_fd_sc_hd__buf_4
XFILLER_33_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14451__A2 _11404_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _12960_/A _12997_/A _12960_/B vssd1 vssd1 vccd1 vccd1 _12998_/X sky130_fd_sc_hd__a21o_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17525_ _19772_/C _17739_/A _17525_/C _17525_/D vssd1 vssd1 vccd1 vccd1 _17531_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16728__A1 _16325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14737_ _14737_/A _14737_/B vssd1 vssd1 vccd1 vccd1 _14738_/A sky130_fd_sc_hd__nand2_1
XFILLER_178_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11949_ _18445_/C _18680_/D _19197_/A _11949_/D vssd1 vssd1 vccd1 vccd1 _11949_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_17_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12462__B2 _15569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16437__A _16669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17456_ _17304_/B _17307_/B _17266_/Y _17262_/X vssd1 vssd1 vccd1 vccd1 _17458_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_14668_ _14561_/D _14561_/Y _14655_/A _14655_/B vssd1 vssd1 vccd1 vccd1 _14752_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16407_ _15881_/Y _16212_/Y _16406_/Y vssd1 vssd1 vccd1 vccd1 _16664_/C sky130_fd_sc_hd__o21bai_2
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _13617_/C _13617_/A _13601_/A _13618_/X vssd1 vssd1 vccd1 vccd1 _13674_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_17387_ _17383_/Y _17385_/Y _17386_/X vssd1 vssd1 vccd1 vccd1 _17550_/A sky130_fd_sc_hd__a21oi_1
X_14599_ _14468_/Y _13873_/X _15069_/A _14461_/Y vssd1 vssd1 vccd1 vccd1 _14600_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_192_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19126_ _18952_/B _18946_/X _18975_/Y vssd1 vssd1 vccd1 vccd1 _19129_/A sky130_fd_sc_hd__a21oi_1
XFILLER_146_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16338_ _16336_/Y _16337_/X _15566_/X vssd1 vssd1 vccd1 vccd1 _16342_/B sky130_fd_sc_hd__o21ai_2
XFILLER_118_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_532 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19057_ _19231_/A _19231_/B _19231_/C vssd1 vssd1 vccd1 vccd1 _19074_/A sky130_fd_sc_hd__nand3_2
X_16269_ _16266_/X _16267_/X _11568_/B _11568_/A _16268_/X vssd1 vssd1 vccd1 vccd1
+ _16269_/X sky130_fd_sc_hd__a221o_2
XFILLER_173_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18008_ _17967_/C _17967_/A _22904_/Q vssd1 vssd1 vccd1 vccd1 _18012_/A sky130_fd_sc_hd__a21o_1
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19483__A _19630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13190__A2 _21580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15467__A1 _15465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19959_ _19959_/A _19959_/B vssd1 vssd1 vccd1 vccd1 _19960_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22861__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21921_ _21931_/B _21931_/A _22089_/A vssd1 vssd1 vccd1 vccd1 _21927_/C sky130_fd_sc_hd__and3_1
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11763__B _22790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19930__B _22923_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17731__A _17731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21852_ _21964_/A _21455_/X _21957_/A vssd1 vssd1 vccd1 vccd1 _21852_/Y sky130_fd_sc_hd__o21ai_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18708__A2 _19160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20803_ _20803_/A _20869_/B _20803_/C vssd1 vssd1 vccd1 vccd1 _20810_/B sky130_fd_sc_hd__nand3_2
XANTENNA__17450__B _17523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21783_ _21485_/X _21649_/A _21645_/Y _21646_/Y vssd1 vssd1 vccd1 vccd1 _21783_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20515__A2 _15935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20734_ _20734_/A _20734_/B _20734_/C _20928_/C vssd1 vssd1 vccd1 vccd1 _20735_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_168_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17392__A1 _16778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12594__B _20130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20665_ _20768_/C _20768_/A _22934_/Q vssd1 vssd1 vccd1 vccd1 _20770_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__15942__A2 _15941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20279__A1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22404_ _22426_/A vssd1 vssd1 vccd1 vccd1 _22413_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20596_ _20596_/A _20702_/A _20596_/C vssd1 vssd1 vccd1 vccd1 _20603_/C sky130_fd_sc_hd__nand3_1
XFILLER_52_1098 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22335_ _22335_/A _22335_/B vssd1 vssd1 vccd1 vccd1 _22338_/A sky130_fd_sc_hd__xnor2_2
XFILLER_87_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16352__C1 _16351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22266_ _22306_/B _21594_/Y _22264_/Y _22302_/A vssd1 vssd1 vccd1 vccd1 _22266_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_3_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21217_ _21183_/X _21212_/Y _21369_/A vssd1 vssd1 vccd1 vccd1 _21237_/B sky130_fd_sc_hd__o21ai_1
XFILLER_151_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19841__B1 _19176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22197_ _22196_/Y _22137_/C _22137_/D vssd1 vssd1 vccd1 vccd1 _22215_/B sky130_fd_sc_hd__a21bo_1
XFILLER_183_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16810__A _19619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20451__A1 _16179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21148_ _21157_/B vssd1 vssd1 vccd1 vccd1 _21149_/A sky130_fd_sc_hd__inv_2
XFILLER_116_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13970_ _14583_/D vssd1 vssd1 vccd1 vccd1 _13970_/X sky130_fd_sc_hd__buf_2
XFILLER_59_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21079_ _21079_/A _21079_/B vssd1 vssd1 vccd1 vccd1 _21079_/Y sky130_fd_sc_hd__nor2_2
XFILLER_101_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12769__B _12769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _12921_/A vssd1 vssd1 vccd1 vccd1 _16059_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17080__B1 _16711_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17641__A _18629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15640_ _15891_/A _15938_/A _15639_/Y vssd1 vssd1 vccd1 vccd1 _15640_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_74_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12852_/A _12852_/B vssd1 vssd1 vccd1 vccd1 _12853_/A sky130_fd_sc_hd__nand2_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _11595_/X _11589_/X _11793_/A _11528_/Y vssd1 vssd1 vccd1 vccd1 _11964_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_55_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15571_ _15571_/A _15571_/B _15571_/C _15571_/D vssd1 vssd1 vccd1 vccd1 _15571_/Y
+ sky130_fd_sc_hd__nand4_4
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12516_/X _15455_/A _20502_/C _15696_/D _12526_/X vssd1 vssd1 vccd1 vccd1
+ _12783_/X sky130_fd_sc_hd__o2111a_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15799__C _16313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_602 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16257__A _16257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17310_ _17310_/A vssd1 vssd1 vccd1 vccd1 _17341_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11734_/A vssd1 vssd1 vccd1 vccd1 _15559_/B sky130_fd_sc_hd__buf_6
XFILLER_25_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14522_ _14522_/A _14522_/B _14522_/C _14522_/D vssd1 vssd1 vccd1 vccd1 _14540_/C
+ sky130_fd_sc_hd__nand4_4
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _17636_/A _18281_/Y _18296_/B _18289_/Y vssd1 vssd1 vccd1 vccd1 _18291_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17383__A1 _15919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_994 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _19047_/B _20928_/A _20928_/B vssd1 vssd1 vccd1 vccd1 _17242_/B sky130_fd_sc_hd__and3_1
X_14453_ _14443_/X _11438_/B _14448_/X vssd1 vssd1 vccd1 vccd1 _22668_/D sky130_fd_sc_hd__a21o_1
X_11665_ _11732_/A vssd1 vssd1 vccd1 vccd1 _16257_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_186_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13404_ _13659_/C _21990_/B vssd1 vssd1 vccd1 vccd1 _13419_/A sky130_fd_sc_hd__nand2_2
XFILLER_70_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17172_ _17172_/A vssd1 vssd1 vccd1 vccd1 _17173_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_14384_ _14593_/B vssd1 vssd1 vccd1 vccd1 _14863_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__17135__A1 _12207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11596_ _11589_/X _11583_/Y _11595_/X vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__a21bo_1
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11955__B1 _11633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16123_ _19012_/C vssd1 vssd1 vccd1 vccd1 _19336_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13335_ _21713_/A _13456_/A _21713_/C vssd1 vssd1 vccd1 vccd1 _13337_/C sky130_fd_sc_hd__and3_1
XFILLER_6_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12614__A2_N _12601_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15697__A1 _18666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20690__A1 _20793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16054_ _18984_/A _18984_/B _16498_/D vssd1 vssd1 vccd1 vccd1 _16110_/B sky130_fd_sc_hd__and3_2
X_13266_ _13650_/B vssd1 vssd1 vccd1 vccd1 _13572_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__20690__B2 _17530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12217_ _12204_/X _12207_/X _11818_/A _12216_/X vssd1 vssd1 vccd1 vccd1 _12217_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15005_ _15006_/A _15005_/B _15006_/C vssd1 vssd1 vccd1 vccd1 _15005_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__17816__A _17816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18635__A1 _18625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ _13521_/A _21494_/B _13521_/C vssd1 vssd1 vccd1 vccd1 _13199_/A sky130_fd_sc_hd__nand3_1
XFILLER_194_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15449__A1 _12929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16720__A _20781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22884__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22441__B input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19813_ _19813_/A _19813_/B vssd1 vssd1 vccd1 vccd1 _19815_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15449__B2 _15455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ _12148_/A _12148_/B _18677_/A vssd1 vssd1 vccd1 vccd1 _12148_/Y sky130_fd_sc_hd__nand3_4
XFILLER_29_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11864__A _18875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19744_ _19741_/X _19808_/B _19747_/A vssd1 vssd1 vccd1 vccd1 _19764_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16956_ _16956_/A _17138_/A vssd1 vssd1 vccd1 vccd1 _16956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12079_ _12079_/A _12079_/B _12079_/C vssd1 vssd1 vccd1 vccd1 _18238_/B sky130_fd_sc_hd__nand3_1
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14672__A2 _13814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19060__A1 _17388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ _15988_/B _16781_/B _18985_/C vssd1 vssd1 vccd1 vccd1 _15907_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__11583__B _11583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19675_ _19675_/A _19827_/A vssd1 vssd1 vccd1 vccd1 _19757_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11486__A2 _11349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16949__A1 _15450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16887_ _17049_/A _17049_/B _16886_/B vssd1 vssd1 vccd1 vccd1 _17048_/D sky130_fd_sc_hd__a21o_1
X_18626_ _16225_/X _16227_/X _18810_/D _17401_/D vssd1 vssd1 vccd1 vccd1 _18626_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _15838_/A vssd1 vssd1 vccd1 vccd1 _15839_/A sky130_fd_sc_hd__buf_2
XFILLER_53_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15621__A1 _15792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14424__A2 _14418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15621__B2 _16397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17270__B _17270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18557_ _18557_/A _18557_/B vssd1 vssd1 vccd1 vccd1 _18561_/A sky130_fd_sc_hd__nand2_1
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15769_ _15769_/A _15769_/B _15769_/C vssd1 vssd1 vccd1 vccd1 _15773_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13632__B1 _21874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17508_ _17508_/A _22898_/Q _17508_/C vssd1 vssd1 vccd1 vccd1 _17508_/Y sky130_fd_sc_hd__nand3_1
XFILLER_177_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18488_ _18488_/A vssd1 vssd1 vccd1 vccd1 _18705_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17439_ _17732_/A vssd1 vssd1 vccd1 vccd1 _17439_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12199__B1 _11727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14118__C _14765_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13935__A1 _13814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20450_ _20449_/A _20449_/B _20449_/C vssd1 vssd1 vccd1 vccd1 _20450_/X sky130_fd_sc_hd__o21a_1
XANTENNA__19197__B _19496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13022__C _13022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11946__B1 _11935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19109_ _18823_/A _18823_/B _18823_/C _18833_/Y vssd1 vssd1 vccd1 vccd1 _19112_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_118_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17677__A2 _17678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20381_ _20403_/C _20378_/B _20379_/X _20380_/Y vssd1 vssd1 vccd1 vccd1 _20381_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_173_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22120_ _22171_/B _22115_/A _22171_/A vssd1 vssd1 vccd1 vccd1 _22190_/B sky130_fd_sc_hd__a21bo_1
XFILLER_161_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput110 _14343_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__22632__A _22643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput121 _22669_/Q vssd1 vssd1 vccd1 vccd1 y[5] sky130_fd_sc_hd__buf_2
XANTENNA__17429__A2 _17111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22051_ _22047_/Y _22049_/X _22099_/A vssd1 vssd1 vccd1 vccd1 _22051_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_161_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21002_ _20961_/Y _20959_/B _21001_/Y vssd1 vssd1 vccd1 vccd1 _21002_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13973__B _13973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16101__A2 _11912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11774__A _19197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19941__A _19941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11493__B _18797_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22953_ _22964_/CLK _22953_/D vssd1 vssd1 vccd1 vccd1 _22953_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__19051__A1 _12157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19051__B2 _15531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21904_ _21909_/B vssd1 vssd1 vccd1 vccd1 _22007_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22884_ _22916_/CLK input78/X vssd1 vssd1 vccd1 vccd1 _22884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21835_ _21837_/A _21837_/D _21837_/C vssd1 vssd1 vccd1 vccd1 _21836_/A sky130_fd_sc_hd__a21boi_2
XFILLER_71_758 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19354__A2 _17380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21766_ _21766_/A _21766_/B vssd1 vssd1 vccd1 vccd1 _21769_/A sky130_fd_sc_hd__nand2_1
XFILLER_196_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20717_ _20717_/A _20717_/B vssd1 vssd1 vccd1 vccd1 _20717_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18292__A _18292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21697_ _21440_/Y _21415_/A _21559_/A _21695_/A _21559_/B vssd1 vssd1 vccd1 vccd1
+ _21698_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12729__A2 _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11450_ _11450_/A vssd1 vssd1 vccd1 vccd1 _18303_/C sky130_fd_sc_hd__buf_2
XFILLER_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20972__D _20972_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20648_ _20648_/A vssd1 vssd1 vccd1 vccd1 _20650_/C sky130_fd_sc_hd__inv_2
XFILLER_165_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11949__A _18445_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _11633_/A vssd1 vssd1 vccd1 vccd1 _11381_/X sky130_fd_sc_hd__clkbuf_4
X_20579_ _20579_/A _20579_/B _20579_/C vssd1 vssd1 vccd1 vccd1 _20579_/X sky130_fd_sc_hd__and3_1
XFILLER_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _13120_/A _13120_/B vssd1 vssd1 vccd1 vccd1 _13120_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_1064 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22318_ _22318_/A _22318_/B vssd1 vssd1 vccd1 vccd1 _22320_/A sky130_fd_sc_hd__xnor2_1
XFILLER_11_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20672__A1 _15941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13586__D _21878_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _22722_/Q _22721_/Q _22720_/Q vssd1 vssd1 vccd1 vccd1 _13067_/A sky130_fd_sc_hd__nor3_4
XANTENNA__17636__A _17636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18617__A1 _17635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22249_ _22250_/C _22250_/A _22683_/Q vssd1 vssd1 vccd1 vccd1 _22294_/A sky130_fd_sc_hd__a21o_1
XFILLER_127_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12002_ _11425_/Y _18508_/A _12001_/Y vssd1 vssd1 vccd1 vccd1 _12017_/A sky130_fd_sc_hd__o21ai_1
XFILLER_105_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input47_A wb_dat_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16810_ _19619_/B _17385_/C _16810_/C _16810_/D vssd1 vssd1 vccd1 vccd1 _16812_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11684__A _12117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17790_ _17800_/D _17800_/A _17790_/C _17790_/D vssd1 vssd1 vccd1 vccd1 _17790_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__16643__A3 _16879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22177__A1 _22176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16741_ _16842_/A _16842_/C _16842_/B vssd1 vssd1 vccd1 vccd1 _16741_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13953_ _14117_/A _22859_/D _14107_/A _14203_/A vssd1 vssd1 vccd1 vccd1 _13954_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19593__A2 _19176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19460_ _14432_/A _15808_/X _11672_/A _19614_/B _19614_/C vssd1 vssd1 vccd1 vccd1
+ _19625_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_35_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12904_ _12904_/A vssd1 vssd1 vccd1 vccd1 _20133_/B sky130_fd_sc_hd__clkbuf_4
X_16672_ _16672_/A vssd1 vssd1 vccd1 vccd1 _16672_/X sky130_fd_sc_hd__clkbuf_2
X_13884_ _13851_/A _13851_/B _13831_/A vssd1 vssd1 vccd1 vccd1 _13884_/X sky130_fd_sc_hd__a21o_1
XFILLER_185_1035 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18411_ _18411_/A _18411_/B _18411_/C vssd1 vssd1 vccd1 vccd1 _18417_/A sky130_fd_sc_hd__nand3_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ _20477_/A vssd1 vssd1 vccd1 vccd1 _20678_/B sky130_fd_sc_hd__clkbuf_4
X_19391_ _19530_/A _19530_/B _19530_/C _19530_/D vssd1 vssd1 vccd1 vccd1 _19392_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12417__A1 _16465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12835_ _20213_/A _20092_/B vssd1 vssd1 vccd1 vccd1 _16708_/A sky130_fd_sc_hd__nand2_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12417__B2 _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19345__A2 _16758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _11541_/A _19464_/A _18349_/A vssd1 vssd1 vccd1 vccd1 _18345_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__13404__A _13659_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15554_ _12913_/A _19687_/B _16215_/A _16215_/B vssd1 vssd1 vccd1 vccd1 _15554_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17356__A1 _17226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16159__A2 _16997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _22827_/Q vssd1 vssd1 vccd1 vccd1 _12767_/A sky130_fd_sc_hd__inv_2
XANTENNA__17356__B2 _17215_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _14818_/A _13924_/X _13926_/Y _13933_/X _14504_/X vssd1 vssd1 vccd1 vccd1
+ _14505_/X sky130_fd_sc_hd__o32a_1
X_11717_ _15536_/A _22658_/B vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__nand2_1
X_18273_ _18271_/Y _18272_/Y _12251_/A vssd1 vssd1 vccd1 vccd1 _18772_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__15367__B1 _15358_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15485_ _15522_/A _15521_/A vssd1 vssd1 vccd1 vccd1 _16217_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15906__A2 _15905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11640__A2 _11505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ _12697_/A vssd1 vssd1 vccd1 vccd1 _13022_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__16715__A _16715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17224_ _22895_/Q _17222_/A _17222_/B _17223_/Y vssd1 vssd1 vccd1 vccd1 _17225_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_175_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14436_ _22966_/Q vssd1 vssd1 vccd1 vccd1 _16242_/B sky130_fd_sc_hd__clkbuf_2
X_11648_ _11647_/A _11647_/B _11635_/X _11641_/X vssd1 vssd1 vccd1 vccd1 _11648_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__21340__B _21498_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 wb_adr_i[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__22101__A1 _21683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput23 wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_2
Xinput34 wb_cyc_i vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_2
XFILLER_190_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17155_ _17155_/A _17155_/B _17155_/C vssd1 vssd1 vccd1 vccd1 _17168_/B sky130_fd_sc_hd__nand3_1
XFILLER_155_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput45 wb_dat_i[19] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
X_11579_ _15357_/A _18663_/A _11529_/Y _11578_/Y vssd1 vssd1 vccd1 vccd1 _11591_/A
+ sky130_fd_sc_hd__a31o_1
X_14367_ _22796_/Q _14354_/X _14355_/X _14361_/X _14366_/X vssd1 vssd1 vccd1 vccd1
+ _14367_/X sky130_fd_sc_hd__a32o_1
Xinput56 wb_dat_i[29] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput67 wb_stb_i vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_2
XANTENNA__12681__C _20101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput78 x[7] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_1
X_16106_ _16106_/A _16106_/B _16106_/C _16106_/D vssd1 vssd1 vccd1 vccd1 _16166_/A
+ sky130_fd_sc_hd__nand4_4
X_13318_ _13633_/A _21220_/A _13316_/X _13317_/X vssd1 vssd1 vccd1 vccd1 _13318_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17086_ _17081_/Y _17084_/X _17085_/Y vssd1 vssd1 vccd1 vccd1 _17086_/Y sky130_fd_sc_hd__o21ai_1
X_14298_ input30/X input29/X input12/X input1/X vssd1 vssd1 vccd1 vccd1 _14300_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_171_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14342__A1 _11980_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16037_ _15962_/X _15959_/X _15947_/Y _15949_/A vssd1 vssd1 vccd1 vccd1 _16038_/C
+ sky130_fd_sc_hd__o211ai_2
X_13249_ _13273_/B vssd1 vssd1 vccd1 vccd1 _21250_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14342__B2 _12413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16450__A _19318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20966__A2 _17424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17988_ _17988_/A _17988_/B vssd1 vssd1 vccd1 vccd1 _17989_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__22168__A1 _13305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19727_ _19605_/B _19605_/C _19605_/A _19611_/X vssd1 vssd1 vccd1 vccd1 _19735_/A
+ sky130_fd_sc_hd__a31o_1
X_16939_ _16934_/X _16937_/Y _16976_/B vssd1 vssd1 vccd1 vccd1 _16939_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__12202__B _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19584__A2 _17400_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17281__A _18659_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19658_ _19658_/A _19658_/B vssd1 vssd1 vccd1 vccd1 _19814_/B sky130_fd_sc_hd__nor2_1
XFILLER_93_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16398__A2 _21050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18609_ _18556_/A _18556_/B _18556_/C _18765_/B _18565_/A vssd1 vssd1 vccd1 vccd1
+ _18609_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_65_596 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19589_ _12207_/X _19464_/A _19500_/X vssd1 vssd1 vccd1 vccd1 _19596_/C sky130_fd_sc_hd__o21ai_2
XFILLER_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21620_ _21383_/X _21606_/X _21766_/A vssd1 vssd1 vccd1 vccd1 _21620_/X sky130_fd_sc_hd__o21a_1
XFILLER_178_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21551_ _21551_/A _21551_/B vssd1 vssd1 vccd1 vccd1 _21695_/A sky130_fd_sc_hd__nand2_2
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20502_ _20502_/A _20502_/B _20502_/C vssd1 vssd1 vccd1 vccd1 _20502_/X sky130_fd_sc_hd__and3_1
XANTENNA__13908__A1 _13820_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21482_ _21482_/A _21482_/B vssd1 vssd1 vccd1 vccd1 _21482_/Y sky130_fd_sc_hd__nand2_2
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19358__D _19358_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20433_ _20834_/A _20835_/A vssd1 vssd1 vccd1 vccd1 _21066_/A sky130_fd_sc_hd__nor2_2
XANTENNA__18847__A1 _11702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20364_ _20364_/A _20446_/A vssd1 vssd1 vccd1 vccd1 _20364_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18206__A_N _18204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22103_ _13305_/A _13305_/B _22102_/Y _22167_/A vssd1 vssd1 vccd1 vccd1 _22129_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14333__A1 _13725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14333__B2 _13202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20295_ _20165_/A _20165_/B _20165_/C vssd1 vssd1 vccd1 vccd1 _20295_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_161_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21603__B1 _21750_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22034_ _22034_/A _22196_/A _22034_/C _22229_/B vssd1 vssd1 vccd1 vccd1 _22131_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_115_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_700 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15833__A1 _16613_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15833__B2 _15834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19024__A1 _19350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19024__B2 _19015_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22936_ _22937_/CLK _22936_/D vssd1 vssd1 vccd1 vccd1 _22936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_708 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15423__B _15774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22867_ _22944_/CLK _22867_/D vssd1 vssd1 vccd1 vccd1 _22867_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17341__D _17341_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13224__A _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12620_ _12456_/Y _12463_/Y _12478_/Y _12479_/X vssd1 vssd1 vccd1 vccd1 _12620_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_189_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21818_ _21837_/C _21837_/D vssd1 vssd1 vccd1 vccd1 _21818_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12804__D1 _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_588 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22798_ _22799_/CLK _22798_/D vssd1 vssd1 vccd1 vccd1 _22798_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18535__B1 _18534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21134__A2 _21086_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12551_ _12669_/A _12528_/A _16328_/A _12470_/X vssd1 vssd1 vccd1 vccd1 _12567_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_157_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21749_ _21749_/A vssd1 vssd1 vccd1 vccd1 _21877_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11622__A2 _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11502_ _11502_/A vssd1 vssd1 vccd1 vccd1 _11502_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_615 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18453__C _18453_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12482_ _17144_/A vssd1 vssd1 vccd1 vccd1 _15774_/C sky130_fd_sc_hd__clkbuf_4
X_15270_ _22876_/D vssd1 vssd1 vccd1 vccd1 _15271_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11679__A _19316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11433_ _11942_/A vssd1 vssd1 vccd1 vccd1 _18288_/A sky130_fd_sc_hd__clkbuf_2
X_14221_ _14255_/A _14255_/C _14255_/B _14256_/A _14256_/B vssd1 vssd1 vccd1 vccd1
+ _14282_/A sky130_fd_sc_hd__a32o_1
XFILLER_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14055__A _14165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_980 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14152_ _14165_/B _14115_/B _14115_/C vssd1 vssd1 vccd1 vccd1 _14153_/A sky130_fd_sc_hd__a21oi_1
XFILLER_164_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11364_ _11429_/A _11421_/A _18115_/C vssd1 vssd1 vccd1 vccd1 _12003_/B sky130_fd_sc_hd__a21o_2
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17510__B2 _17719_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13103_ _22842_/Q vssd1 vssd1 vccd1 vccd1 _21595_/B sky130_fd_sc_hd__buf_2
XANTENNA__14324__A1 _12876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13894__A _22761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18960_ _19138_/D _18960_/B _18960_/C vssd1 vssd1 vccd1 vccd1 _19279_/B sky130_fd_sc_hd__nand3_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14324__B2 _13659_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14083_ _14083_/A vssd1 vssd1 vccd1 vccd1 _14161_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_180_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11295_ _11295_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11968_/B sky130_fd_sc_hd__nand2_2
XANTENNA__22398__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ _17226_/X _17227_/X _17959_/A _17959_/B _17910_/Y vssd1 vssd1 vccd1 vccd1
+ _17915_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_180_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _12944_/X _12991_/X _12993_/X _12990_/A _13031_/A vssd1 vssd1 vccd1 vccd1
+ _13035_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_152_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18891_ _11636_/X _18889_/X _18890_/X _19587_/B _18980_/A vssd1 vssd1 vccd1 vccd1
+ _18891_/X sky130_fd_sc_hd__o311a_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16077__A1 _15972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17842_ _17842_/A _17842_/B vssd1 vssd1 vccd1 vccd1 _17904_/A sky130_fd_sc_hd__xnor2_2
XFILLER_26_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19015__A1 _14431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17773_ _17701_/A _17701_/C _17701_/B vssd1 vssd1 vccd1 vccd1 _17785_/B sky130_fd_sc_hd__a21boi_1
XFILLER_120_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14985_ _14924_/A _14927_/B _15039_/A _14984_/Y _14982_/B vssd1 vssd1 vccd1 vccd1
+ _14985_/X sky130_fd_sc_hd__o221a_1
XANTENNA__22922__CLK _22922_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19512_ _19512_/A _19512_/B vssd1 vssd1 vccd1 vccd1 _19521_/D sky130_fd_sc_hd__nand2_1
X_16724_ _19470_/B _19470_/D _17385_/C _20593_/A vssd1 vssd1 vccd1 vccd1 _16724_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__15614__A _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13936_ _13935_/X _13931_/X _13933_/X vssd1 vssd1 vccd1 vccd1 _13937_/D sky130_fd_sc_hd__a21o_1
XANTENNA__17532__C _17532_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19443_ _19443_/A vssd1 vssd1 vccd1 vccd1 _19680_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16655_ _16441_/X _17078_/A _16659_/A vssd1 vssd1 vccd1 vccd1 _16889_/B sky130_fd_sc_hd__o21bai_2
XFILLER_62_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13867_ _13867_/A vssd1 vssd1 vccd1 vccd1 _14169_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15606_ _20461_/A vssd1 vssd1 vccd1 vccd1 _20463_/A sky130_fd_sc_hd__buf_2
X_19374_ _19374_/A _19374_/B vssd1 vssd1 vccd1 vccd1 _19379_/B sky130_fd_sc_hd__nand2_1
X_12818_ _12818_/A _12818_/B _12818_/C vssd1 vssd1 vccd1 vccd1 _12852_/B sky130_fd_sc_hd__nand3_1
X_16586_ _16586_/A _16586_/B _17313_/B _16879_/A vssd1 vssd1 vccd1 vccd1 _16586_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20425__A2_N _20432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13798_ _13798_/A vssd1 vssd1 vccd1 vccd1 _13820_/A sky130_fd_sc_hd__buf_2
XFILLER_43_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18325_ _18325_/A vssd1 vssd1 vccd1 vccd1 _19496_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_163_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15537_ _14430_/A _16241_/C _16226_/B _15536_/X vssd1 vssd1 vccd1 vccd1 _15548_/A
+ sky130_fd_sc_hd__o211ai_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12749_/A _12749_/B vssd1 vssd1 vccd1 vccd1 _12750_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18256_ _18249_/A _12249_/A _18772_/B _18772_/C vssd1 vssd1 vccd1 vccd1 _18257_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15468_ _15308_/A _15472_/A _15574_/C vssd1 vssd1 vccd1 vccd1 _15477_/A sky130_fd_sc_hd__o21ai_1
XFILLER_124_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17207_ _17208_/A _17208_/B _17208_/C vssd1 vssd1 vccd1 vccd1 _17603_/C sky130_fd_sc_hd__a21oi_2
XFILLER_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14419_ _22811_/Q _14411_/X _14412_/X _14413_/X _22779_/Q vssd1 vssd1 vccd1 vccd1
+ _14419_/X sky130_fd_sc_hd__a32o_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18187_ _18404_/A _18187_/B vssd1 vssd1 vccd1 vccd1 _18187_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13220__D1 _21638_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15399_ _16257_/C vssd1 vssd1 vccd1 vccd1 _20502_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__20097__C1 _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17138_ _17138_/A vssd1 vssd1 vccd1 vccd1 _17138_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18844__A4 _16062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17069_ _22893_/Q _16702_/Y _16899_/Y _16901_/Y vssd1 vssd1 vccd1 vccd1 _17070_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__18810__D _18810_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19194__C _19490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22389__A1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20080_ _20080_/A vssd1 vssd1 vccd1 vccd1 _20293_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17426__D _19614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16068__B2 _16155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11755__C _18303_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12629__A1 _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20982_ _20982_/A _20982_/B _20982_/C vssd1 vssd1 vccd1 vccd1 _20985_/C sky130_fd_sc_hd__or3_1
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15579__B1 _15546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22721_ input33/X _22721_/D vssd1 vssd1 vccd1 vccd1 _22721_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11852__A2 _11845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16058__C _16058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1096 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22652_ _22813_/Q input56/X _22652_/S vssd1 vssd1 vccd1 vccd1 _22653_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16791__A2 _16779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21603_ _21482_/B _21751_/A _21750_/C _21758_/A _22184_/A vssd1 vssd1 vccd1 vccd1
+ _21604_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22583_ _22583_/A vssd1 vssd1 vccd1 vccd1 _22782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21534_ _21545_/A _21545_/B vssd1 vssd1 vccd1 vccd1 _21534_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17740__A1 _15941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11499__A _12154_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21465_ _21805_/D _21514_/C _21666_/B vssd1 vssd1 vccd1 vccd1 _21465_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_193_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11368__A1 _15932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_991 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20416_ _20449_/A vssd1 vssd1 vccd1 vccd1 _20844_/A sky130_fd_sc_hd__clkbuf_4
X_21396_ _21245_/A _21395_/Y _21181_/A vssd1 vssd1 vccd1 vccd1 _21445_/A sky130_fd_sc_hd__o21ai_1
XFILLER_146_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20347_ _20347_/A _20347_/B vssd1 vssd1 vccd1 vccd1 _20347_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14603__A _14892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20278_ _12761_/X _15890_/X _20155_/B _20144_/Y _20155_/C vssd1 vssd1 vccd1 vccd1
+ _20284_/C sky130_fd_sc_hd__o221ai_4
XANTENNA__22945__CLK _22948_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22017_ _22086_/A _22086_/B _22155_/A _22145_/A vssd1 vssd1 vccd1 vccd1 _22017_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12123__A _18208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15806__A1 _15810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15267__C1 _15260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13817__B1 _14122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17008__B1 _15936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14770_ _14770_/A vssd1 vssd1 vccd1 vccd1 _15107_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11982_ _11789_/X _11791_/X _11794_/A _11797_/B vssd1 vssd1 vccd1 vccd1 _11982_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1024 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13721_ _14065_/A vssd1 vssd1 vccd1 vccd1 _13728_/A sky130_fd_sc_hd__buf_2
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22919_ _22922_/CLK _22919_/D vssd1 vssd1 vccd1 vccd1 _22919_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__16767__C1 _15577_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18745__A _18933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_555 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16231__A1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16440_ _16206_/A _15879_/A _16433_/Y vssd1 vssd1 vccd1 vccd1 _16440_/Y sky130_fd_sc_hd__o21ai_1
X_13652_ _21398_/B _21195_/C _21398_/A _21195_/B _13650_/A vssd1 vssd1 vccd1 vccd1
+ _13657_/B sky130_fd_sc_hd__a32o_1
XFILLER_72_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12603_ _20338_/C vssd1 vssd1 vccd1 vccd1 _20463_/C sky130_fd_sc_hd__clkbuf_4
X_16371_ _15666_/A _15668_/X _15673_/C vssd1 vssd1 vccd1 vccd1 _16371_/Y sky130_fd_sc_hd__o21ai_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _21195_/C vssd1 vssd1 vccd1 vccd1 _13664_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15990__B1 _11911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18110_ _18810_/A _18848_/D _18367_/C _18848_/C vssd1 vssd1 vccd1 vccd1 _18110_/X
+ sky130_fd_sc_hd__and4_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _15315_/Y _15343_/A _15321_/Y vssd1 vssd1 vccd1 vccd1 _15339_/A sky130_fd_sc_hd__o21ai_2
X_19090_ _19033_/X _19039_/Y _19082_/Y _19106_/A vssd1 vssd1 vccd1 vccd1 _19117_/B
+ sky130_fd_sc_hd__o211ai_2
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12970_/A vssd1 vssd1 vccd1 vccd1 _16759_/A sky130_fd_sc_hd__buf_2
XFILLER_12_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18041_ _18019_/Y _17999_/A _18042_/A _18040_/Y vssd1 vssd1 vccd1 vccd1 _18049_/A
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__14545__A1 _14561_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15253_ _15238_/A _15224_/A _15238_/B vssd1 vssd1 vccd1 vccd1 _15253_/Y sky130_fd_sc_hd__o21ai_1
X_12465_ _20086_/A _20207_/C _20478_/C _17141_/A vssd1 vssd1 vccd1 vccd1 _12479_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_172_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20618__A1 _17407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14204_ _14693_/D vssd1 vssd1 vccd1 vccd1 _14861_/C sky130_fd_sc_hd__buf_2
XFILLER_184_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11416_ _18115_/C vssd1 vssd1 vccd1 vccd1 _11420_/D sky130_fd_sc_hd__inv_2
XFILLER_193_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15184_ _15217_/A _15056_/A _15056_/B _15160_/A vssd1 vssd1 vccd1 vccd1 _15186_/B
+ sky130_fd_sc_hd__a31o_1
X_12396_ _12396_/A _12520_/B _12396_/C vssd1 vssd1 vccd1 vccd1 _12586_/A sky130_fd_sc_hd__nand3_1
XFILLER_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12017__B _18367_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16712__B _20471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ _13948_/X _13949_/X _13748_/X vssd1 vssd1 vccd1 vccd1 _14135_/X sky130_fd_sc_hd__a21o_1
X_11347_ _11496_/B vssd1 vssd1 vccd1 vccd1 _18099_/A sky130_fd_sc_hd__buf_2
XFILLER_193_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19992_ _20037_/C _19992_/B _19992_/C vssd1 vssd1 vccd1 vccd1 _19994_/A sky130_fd_sc_hd__or3_1
XFILLER_4_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18943_ _18937_/Y _18938_/Y _18932_/Y _18935_/A vssd1 vssd1 vccd1 vccd1 _18945_/B
+ sky130_fd_sc_hd__o211ai_4
X_14066_ _13857_/X _13725_/Y _14684_/B _14834_/A vssd1 vssd1 vccd1 vccd1 _14126_/B
+ sky130_fd_sc_hd__o211a_1
X_11278_ _11306_/A _11385_/C _11273_/X _11783_/C _11420_/C vssd1 vssd1 vccd1 vccd1
+ _11285_/A sky130_fd_sc_hd__o311ai_4
XFILLER_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13017_ _13024_/B _12681_/A _12681_/B _12989_/A _12975_/D vssd1 vssd1 vccd1 vccd1
+ _13017_/X sky130_fd_sc_hd__a32o_1
X_18874_ _18695_/X _18696_/X _18707_/B _18692_/Y vssd1 vssd1 vccd1 vccd1 _18883_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17825_ _17826_/A _17826_/B _17826_/C vssd1 vssd1 vccd1 vccd1 _17890_/A sky130_fd_sc_hd__a21o_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_658 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12968__A _12968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17756_ _17745_/X _17826_/B _17744_/A vssd1 vssd1 vccd1 vccd1 _17756_/Y sky130_fd_sc_hd__a21oi_1
X_14968_ _14968_/A _14968_/B vssd1 vssd1 vccd1 vccd1 _14969_/B sky130_fd_sc_hd__nor2_1
XFILLER_94_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22543__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12687__B _12687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16707_ _16620_/A _16620_/B _16620_/C _16706_/Y vssd1 vssd1 vccd1 vccd1 _16707_/Y
+ sky130_fd_sc_hd__a31oi_2
X_13919_ _13881_/A _13986_/A _13873_/A _13877_/Y _14808_/A vssd1 vssd1 vccd1 vccd1
+ _13920_/C sky130_fd_sc_hd__o2111ai_1
X_17687_ _17687_/A _17687_/B _17687_/C vssd1 vssd1 vccd1 vccd1 _17688_/C sky130_fd_sc_hd__nand3_1
XFILLER_62_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14899_ _14899_/A _14899_/B vssd1 vssd1 vccd1 vccd1 _14901_/C sky130_fd_sc_hd__nor2_1
X_19426_ _19255_/Y _19303_/Y _19253_/Y _19434_/B vssd1 vssd1 vccd1 vccd1 _19427_/D
+ sky130_fd_sc_hd__a31o_1
X_16638_ _16637_/A _16637_/B _16630_/B _16630_/A vssd1 vssd1 vccd1 vccd1 _16638_/Y
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_63_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19357_ _19357_/A _19357_/B vssd1 vssd1 vccd1 vccd1 _19357_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13587__A2 _21489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16569_ _11800_/X _17874_/A _17875_/A _16563_/Y vssd1 vssd1 vccd1 vccd1 _16570_/A
+ sky130_fd_sc_hd__o31ai_1
XANTENNA__19172__B1 _19334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22818__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18308_ _18571_/D _18442_/B _18309_/A vssd1 vssd1 vccd1 vccd1 _18308_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18093__C _18093_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19288_ _22916_/Q _19288_/B vssd1 vssd1 vccd1 vccd1 _19288_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18239_ _18272_/A _18239_/B _18239_/C vssd1 vssd1 vccd1 vccd1 _18240_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13311__B _21476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21250_ _21250_/A _22850_/Q _21250_/C vssd1 vssd1 vccd1 vccd1 _21251_/C sky130_fd_sc_hd__and3_1
XANTENNA__21806__B1 _21805_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19475__A1 _19476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12011__A2 _19350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20201_ _20198_/Y _20158_/B _20167_/B _20200_/X vssd1 vssd1 vccd1 vccd1 _20286_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20085__A2 _20359_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21181_ _21181_/A _21181_/B vssd1 vssd1 vccd1 vccd1 _21245_/B sky130_fd_sc_hd__nand2_1
XFILLER_143_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20132_ _20249_/B _15899_/B _20134_/B _20129_/Y _20131_/Y vssd1 vssd1 vccd1 vccd1
+ _20132_/X sky130_fd_sc_hd__a32o_2
XFILLER_131_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17238__B1 _18203_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20063_ _20063_/A _20063_/B vssd1 vssd1 vccd1 vccd1 _22908_/D sky130_fd_sc_hd__nor2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15264__A2 _15260_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22534__A1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20965_ _20843_/X _15941_/X _20933_/B _20930_/Y _17928_/A vssd1 vssd1 vccd1 vccd1
+ _20987_/A sky130_fd_sc_hd__o32a_2
XFILLER_65_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22704_ _22800_/CLK _22704_/D vssd1 vssd1 vccd1 vccd1 _22704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__A1 _13022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20896_ _20906_/C vssd1 vssd1 vccd1 vccd1 _20897_/B sky130_fd_sc_hd__inv_2
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16764__A2 _16758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22635_ _22805_/Q input48/X _22641_/S vssd1 vssd1 vccd1 vccd1 _22636_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15972__B1 _12772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19702__A2 _17388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22566_ _22566_/A vssd1 vssd1 vccd1 vccd1 _22774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1085 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16516__A2 _12696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21517_ _21538_/A _21537_/A _21538_/B vssd1 vssd1 vccd1 vccd1 _21531_/A sky130_fd_sc_hd__nand3_1
XFILLER_6_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22497_ _22744_/Q input51/X _22497_/S vssd1 vssd1 vccd1 vccd1 _22498_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16813__A _16831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12118__A _12118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12250_ _18249_/A _18236_/B _18272_/B _12250_/D vssd1 vssd1 vccd1 vccd1 _12251_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19466__A1 _14432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21448_ _21448_/A _21448_/B _21448_/C vssd1 vssd1 vccd1 vccd1 _21449_/B sky130_fd_sc_hd__nand3_2
XFILLER_170_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _12181_/A _12181_/B _12181_/C vssd1 vssd1 vccd1 vccd1 _12182_/D sky130_fd_sc_hd__nand3_2
X_21379_ _21379_/A _21393_/C vssd1 vssd1 vccd1 vccd1 _21535_/A sky130_fd_sc_hd__nand2_1
XFILLER_122_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15940_ _15940_/A vssd1 vssd1 vccd1 vccd1 _15941_/A sky130_fd_sc_hd__buf_2
XFILLER_27_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_912 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11513__A1 _11511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18459__B _19687_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14987__B _15046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15871_ _15415_/X _15870_/X _15703_/B vssd1 vssd1 vccd1 vccd1 _16034_/C sky130_fd_sc_hd__o21ai_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12788__A _16489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17610_ _17607_/X _17713_/A _22899_/Q vssd1 vssd1 vccd1 vccd1 _17610_/Y sky130_fd_sc_hd__a21oi_1
X_14822_ _14822_/A _14902_/A _14822_/C vssd1 vssd1 vccd1 vccd1 _14902_/B sky130_fd_sc_hd__nand3_1
X_18590_ _18590_/A vssd1 vssd1 vccd1 vccd1 _19294_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22525__A1 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _17394_/Y _17402_/Y _17536_/X _17540_/Y vssd1 vssd1 vccd1 vccd1 _17541_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12474__C1 _16319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14753_ _14750_/A _14750_/B _14751_/A vssd1 vssd1 vccd1 vccd1 _14756_/A sky130_fd_sc_hd__a21o_1
XFILLER_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _11846_/Y _11774_/Y _11945_/B vssd1 vssd1 vccd1 vccd1 _11965_/X sky130_fd_sc_hd__a21o_1
XANTENNA__20536__B1 _20263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output116_A _22952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13704_ _13707_/A vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__buf_2
X_17472_ _17486_/B _17472_/B vssd1 vssd1 vccd1 vccd1 _17473_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13018__A1 _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14684_ _14684_/A _14684_/B _14684_/C vssd1 vssd1 vccd1 vccd1 _14685_/B sky130_fd_sc_hd__nand3_4
XFILLER_60_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16755__A2 _16753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11896_ _11896_/A _11896_/B _11896_/C vssd1 vssd1 vccd1 vccd1 _11909_/C sky130_fd_sc_hd__nand3_4
X_19211_ _19211_/A _19418_/B _19211_/C vssd1 vssd1 vccd1 vccd1 _19211_/X sky130_fd_sc_hd__and3_1
X_16423_ _16038_/B _15964_/Y _16203_/Y _16422_/Y vssd1 vssd1 vccd1 vccd1 _16424_/C
+ sky130_fd_sc_hd__o211ai_2
X_13635_ _13635_/A _21878_/C _13664_/A _13650_/A vssd1 vssd1 vccd1 vccd1 _13657_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__15963__B1 _15959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19142_ _19290_/A _19142_/B vssd1 vssd1 vccd1 vccd1 _19145_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16354_ _16354_/A _16617_/A _16354_/C vssd1 vssd1 vccd1 vccd1 _16355_/C sky130_fd_sc_hd__nand3_1
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ _13565_/Y _13524_/X _13526_/A _13526_/B vssd1 vssd1 vccd1 vccd1 _13566_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15305_ _15298_/Y _15309_/A _15304_/Y vssd1 vssd1 vccd1 vccd1 _15313_/A sky130_fd_sc_hd__o21ai_1
XFILLER_118_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19073_ _11625_/X _11626_/X _19585_/D _19046_/A _19065_/X vssd1 vssd1 vccd1 vccd1
+ _19074_/D sky130_fd_sc_hd__o2111ai_4
X_12517_ _22825_/Q vssd1 vssd1 vccd1 vccd1 _20134_/C sky130_fd_sc_hd__clkbuf_2
X_16285_ _16606_/A _16606_/B _16606_/C vssd1 vssd1 vccd1 vccd1 _16377_/A sky130_fd_sc_hd__nand3_1
XFILLER_9_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13497_ _13498_/A _13498_/B _13498_/C vssd1 vssd1 vccd1 vccd1 _13497_/X sky130_fd_sc_hd__and3_1
X_18024_ _19983_/B vssd1 vssd1 vccd1 vccd1 _18778_/D sky130_fd_sc_hd__buf_2
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15236_ _15217_/A _15217_/B _15217_/C _15224_/D vssd1 vssd1 vccd1 vccd1 _15243_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12448_ _15394_/A _16257_/C _16256_/D _20694_/A vssd1 vssd1 vccd1 vccd1 _12448_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_154_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15339__A _15339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11867__A _19154_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ _15181_/A _15168_/C _15168_/A vssd1 vssd1 vccd1 vccd1 _15169_/B sky130_fd_sc_hd__o21a_1
XFILLER_141_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12379_ _12379_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _15352_/A sky130_fd_sc_hd__nand2_2
XFILLER_158_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14118_ _14765_/A _14118_/B _14765_/C vssd1 vssd1 vccd1 vccd1 _14118_/Y sky130_fd_sc_hd__nand3_1
XFILLER_125_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19975_ _19975_/A vssd1 vssd1 vccd1 vccd1 _19975_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15098_ _15098_/A _15098_/B _15098_/C vssd1 vssd1 vccd1 vccd1 _15100_/A sky130_fd_sc_hd__nand3_1
XANTENNA__16691__A1 _16669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15494__A2 _12719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18926_ _18929_/A _18929_/B _18978_/A _18931_/B vssd1 vssd1 vccd1 vccd1 _18938_/B
+ sky130_fd_sc_hd__a22o_1
X_14049_ _14049_/A _14049_/B vssd1 vssd1 vccd1 vccd1 _14103_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18857_ _18857_/A vssd1 vssd1 vccd1 vccd1 _19480_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_926 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17808_ _17833_/C vssd1 vssd1 vccd1 vccd1 _21017_/B sky130_fd_sc_hd__buf_2
X_18788_ _18788_/A _18969_/A _18969_/B vssd1 vssd1 vccd1 vccd1 _18789_/B sky130_fd_sc_hd__or3_1
XANTENNA__14454__B1 _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17739_ _17739_/A _19769_/B _19768_/D _20806_/C vssd1 vssd1 vccd1 vccd1 _17826_/A
+ sky130_fd_sc_hd__nand4_4
XANTENNA__18196__A1 _15530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12210__B _22662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20750_ _20751_/A _20751_/C _20751_/B vssd1 vssd1 vccd1 vccd1 _20758_/A sky130_fd_sc_hd__o21a_1
XFILLER_126_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19409_ _19244_/Y _19400_/X _19407_/X _19408_/X vssd1 vssd1 vccd1 vccd1 _19410_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20681_ _20682_/C _20682_/A _20482_/A _20680_/X vssd1 vssd1 vccd1 vccd1 _20683_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_195_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22420_ _22710_/Q input49/X _22424_/S vssd1 vssd1 vccd1 vccd1 _22421_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19696__B2 _17388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22351_ _22338_/A _22341_/A _22341_/C _22341_/B vssd1 vssd1 vccd1 vccd1 _22352_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13041__B _13045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21302_ _22729_/Q _22728_/Q vssd1 vssd1 vccd1 vccd1 _21583_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11991__A1 _22792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22282_ _22317_/B _22282_/B vssd1 vssd1 vccd1 vccd1 _22300_/A sky130_fd_sc_hd__nor2_1
XFILLER_191_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11777__A _18445_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21233_ _13346_/X _21216_/A _13329_/X _21944_/A _21805_/B vssd1 vssd1 vccd1 vccd1
+ _21233_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_191_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15249__A _15259_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1034 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21164_ _21164_/A _21164_/B vssd1 vssd1 vccd1 vccd1 _21164_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22370__A _22426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16682__A1 _17502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20115_ _20115_/A _20115_/B _20115_/C vssd1 vssd1 vccd1 vccd1 _20116_/A sky130_fd_sc_hd__nand3_1
X_21095_ _21095_/A _21095_/B _21095_/C vssd1 vssd1 vccd1 vccd1 _21095_/Y sky130_fd_sc_hd__nand3_1
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20046_ _20025_/X _20032_/B _20042_/Y _20044_/Y vssd1 vssd1 vccd1 vccd1 _20059_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19620__A1 _17436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19620__B2 _19614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15415__C _15415_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _22029_/A _21994_/A _22029_/B vssd1 vssd1 vccd1 vccd1 _21997_/Y sky130_fd_sc_hd__a21boi_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11750_ _11750_/A vssd1 vssd1 vccd1 vccd1 _17422_/A sky130_fd_sc_hd__buf_2
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21433__B _22674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20949_/B _20949_/C _20949_/A vssd1 vssd1 vccd1 vccd1 _20992_/A sky130_fd_sc_hd__o21ai_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15431__B _15700_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11681_ _11675_/A _11675_/B _15482_/B _11560_/C _11667_/Y vssd1 vssd1 vccd1 vccd1
+ _15297_/A sky130_fd_sc_hd__a41o_2
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20879_ _20879_/A _20941_/A _20879_/C vssd1 vssd1 vccd1 vccd1 _20941_/B sky130_fd_sc_hd__nand3_1
XFILLER_81_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16246__C _16515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13420_ _13494_/B _13495_/B _13495_/A vssd1 vssd1 vccd1 vccd1 _13491_/B sky130_fd_sc_hd__nand3_1
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22618_ _22618_/A vssd1 vssd1 vccd1 vccd1 _22797_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18344__D1 _15624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13351_ _13147_/A _13147_/B _13329_/X _13337_/B _21767_/A vssd1 vssd1 vccd1 vccd1
+ _13351_/Y sky130_fd_sc_hd__a221oi_4
XFILLER_194_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22549_ _22571_/A vssd1 vssd1 vccd1 vccd1 _22558_/S sky130_fd_sc_hd__buf_2
XFILLER_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21125__A1_N _22942_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12302_ _12396_/C vssd1 vssd1 vccd1 vccd1 _12387_/B sky130_fd_sc_hd__buf_2
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16070_ _16068_/Y _16055_/Y _16069_/X vssd1 vssd1 vccd1 vccd1 _16070_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_155_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input77_A x[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13282_ _13413_/A _13282_/B vssd1 vssd1 vccd1 vccd1 _13282_/Y sky130_fd_sc_hd__nand2_1
XFILLER_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ _15018_/X _15019_/Y _14959_/C _14960_/B vssd1 vssd1 vccd1 vccd1 _15030_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ _15445_/A vssd1 vssd1 vccd1 vccd1 _15530_/A sky130_fd_sc_hd__buf_2
XFILLER_136_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18111__A1 _19046_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12931__B1 _12718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ _12156_/X _12162_/Y _12163_/X vssd1 vssd1 vccd1 vccd1 _12164_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_162_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14998__A _14998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19760_ _19760_/A _19760_/B vssd1 vssd1 vccd1 vccd1 _19880_/B sky130_fd_sc_hd__nand2_1
X_16972_ _16972_/A _16972_/B vssd1 vssd1 vccd1 vccd1 _16972_/Y sky130_fd_sc_hd__nand2_1
X_12095_ _12090_/X _12094_/Y _12001_/Y vssd1 vssd1 vccd1 vccd1 _12102_/A sky130_fd_sc_hd__a21boi_2
XFILLER_123_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18711_ _18491_/A _18916_/A _18916_/B vssd1 vssd1 vccd1 vccd1 _18713_/B sky130_fd_sc_hd__a21o_1
X_15923_ _16011_/A _16011_/B vssd1 vssd1 vccd1 vccd1 _16009_/C sky130_fd_sc_hd__nand2_1
X_19691_ _19590_/X _19596_/B _19690_/X vssd1 vssd1 vccd1 vccd1 _19698_/A sky130_fd_sc_hd__a21oi_1
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20757__B1 _20759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14510__B _14629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18642_ _18635_/X _18637_/X _18619_/Y _18835_/A vssd1 vssd1 vccd1 vccd1 _18933_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _15854_/A _15854_/B _15864_/B vssd1 vssd1 vccd1 vccd1 _15855_/D sky130_fd_sc_hd__nand3_1
XFILLER_188_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14805_ _14805_/A _14895_/B _14805_/C _14805_/D vssd1 vssd1 vccd1 vccd1 _14806_/C
+ sky130_fd_sc_hd__nand4_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _18761_/A _18575_/B _18571_/X _18572_/X vssd1 vssd1 vccd1 vccd1 _18578_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _11295_/A _11295_/B _16465_/A vssd1 vssd1 vccd1 vccd1 _16192_/B sky130_fd_sc_hd__a21oi_4
X_12997_ _12997_/A vssd1 vssd1 vccd1 vccd1 _12997_/Y sky130_fd_sc_hd__inv_2
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17524_ _17452_/A _17457_/D _17457_/C vssd1 vssd1 vccd1 vccd1 _17524_/Y sky130_fd_sc_hd__a21boi_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _14740_/A _14740_/B _14734_/Y _14735_/X vssd1 vssd1 vccd1 vccd1 _14745_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_11948_ _15633_/A vssd1 vssd1 vccd1 vccd1 _18680_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_73_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16728__A2 _16325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_620 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16437__B _16670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17455_ _17457_/A _17523_/C _17457_/C _17457_/D vssd1 vssd1 vccd1 vccd1 _17458_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _14843_/A _14843_/B _14843_/C _14845_/B vssd1 vssd1 vccd1 vccd1 _14762_/A
+ sky130_fd_sc_hd__a31o_1
X_11879_ _11429_/A _18258_/A _11420_/D vssd1 vssd1 vccd1 vccd1 _11879_/Y sky130_fd_sc_hd__a21oi_2
X_16406_ _16406_/A _16406_/B vssd1 vssd1 vccd1 vccd1 _16406_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17446__A1_N _17523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13618_ _13618_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _13618_/X sky130_fd_sc_hd__and2_1
X_17386_ _19694_/A _17386_/B _20675_/B vssd1 vssd1 vccd1 vccd1 _17386_/X sky130_fd_sc_hd__and3_1
X_14598_ _14468_/B _14685_/A _15010_/A _13873_/X _14568_/Y vssd1 vssd1 vccd1 vccd1
+ _14600_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__22455__A _22512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19125_ _18975_/Y _18950_/A _19121_/Y _19124_/X vssd1 vssd1 vccd1 vccd1 _19147_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_146_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16337_ _12114_/X _16179_/A _15309_/B _15470_/B _15579_/X vssd1 vssd1 vccd1 vccd1
+ _16337_/X sky130_fd_sc_hd__o32a_1
XFILLER_186_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13549_ _13614_/C _13614_/B _13614_/A vssd1 vssd1 vccd1 vccd1 _13551_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__12981__A _15577_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19056_ _12216_/X _19048_/Y _17632_/A _19651_/A _19055_/Y vssd1 vssd1 vccd1 vccd1
+ _19231_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_173_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16268_ _16268_/A vssd1 vssd1 vccd1 vccd1 _16268_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18007_ _18007_/A _18007_/B _18007_/C _18007_/D vssd1 vssd1 vccd1 vccd1 _18053_/A
+ sky130_fd_sc_hd__nand4_1
X_15219_ _15115_/A _15115_/B _15154_/A _15188_/A vssd1 vssd1 vccd1 vccd1 _15224_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_127_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16199_ _15966_/X _15921_/X _16198_/Y _16024_/Y vssd1 vssd1 vccd1 vccd1 _16201_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_114_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19483__B _19630_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19958_ _19959_/A _19959_/B vssd1 vssd1 vccd1 vccd1 _20001_/A sky130_fd_sc_hd__or2_1
XFILLER_113_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17715__C _22900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18909_ _18909_/A vssd1 vssd1 vccd1 vccd1 _18912_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_1081 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19889_ _19889_/A _19889_/B vssd1 vssd1 vccd1 vccd1 _22902_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21920_ _21931_/B _22089_/A _21931_/A vssd1 vssd1 vccd1 vccd1 _21927_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12221__A _12221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21851_ _21851_/A _22041_/B _21851_/C vssd1 vssd1 vccd1 vccd1 _21957_/A sky130_fd_sc_hd__nand3_4
XANTENNA__18169__A1 _19470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18546__C _18546_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20802_ _20869_/B _20803_/C _20803_/A vssd1 vssd1 vccd1 vccd1 _20810_/A sky130_fd_sc_hd__a21o_1
XFILLER_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_683 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21782_ _21799_/B _21802_/C vssd1 vssd1 vccd1 vccd1 _21782_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20733_ _20928_/C _16129_/C _16078_/B _20734_/B _20734_/C vssd1 vssd1 vccd1 vccd1
+ _20735_/A sky130_fd_sc_hd__a32o_1
XFILLER_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17392__A2 _16779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20664_ _20827_/A _20827_/B _20827_/C _20764_/A vssd1 vssd1 vccd1 vccd1 _20768_/A
+ sky130_fd_sc_hd__nand4b_2
XFILLER_196_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18326__D1 _19496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22403_ _22403_/A vssd1 vssd1 vccd1 vccd1 _22702_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__20279__A2 _12525_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20595_ _20595_/A _20682_/B vssd1 vssd1 vccd1 vccd1 _20596_/C sky130_fd_sc_hd__nor2_1
XFILLER_13_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15155__A1 _15188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22334_ _22316_/A _22318_/B _22316_/B vssd1 vssd1 vccd1 vccd1 _22335_/B sky130_fd_sc_hd__o21bai_2
XANTENNA__15155__B2 _14503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22265_ _22264_/Y _22265_/B _22265_/C vssd1 vssd1 vccd1 vccd1 _22302_/B sky130_fd_sc_hd__nand3b_1
XFILLER_151_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21216_ _21216_/A _21216_/B vssd1 vssd1 vccd1 vccd1 _21369_/A sky130_fd_sc_hd__nand2_2
XFILLER_144_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22196_ _22196_/A _22196_/B vssd1 vssd1 vccd1 vccd1 _22196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16810__B _17385_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22686__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20451__A2 _20728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21147_ _21147_/A _21151_/B vssd1 vssd1 vccd1 vccd1 _22925_/D sky130_fd_sc_hd__xor2_1
XFILLER_160_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14611__A _14611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21078_ _21124_/B _21124_/A vssd1 vssd1 vccd1 vccd1 _22921_/D sky130_fd_sc_hd__xor2_1
XFILLER_24_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20739__B1 _20735_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20029_ _20042_/B _20029_/B _20029_/C vssd1 vssd1 vccd1 vccd1 _20030_/A sky130_fd_sc_hd__nand3_1
XANTENNA__17922__A _17922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12920_ _13002_/A _13002_/B _12920_/C vssd1 vssd1 vccd1 vccd1 _12963_/B sky130_fd_sc_hd__nand3_1
XFILLER_100_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17080__A1 _16580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12851_ _12851_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12851_/Y sky130_fd_sc_hd__nand2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11970__A _18648_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15442__A _16473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11802_ _11789_/X _11791_/X _18665_/A _15624_/A _11976_/A vssd1 vssd1 vccd1 vccd1
+ _11964_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_15_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15580_/A _16039_/A _15559_/Y _15558_/Y _15563_/Y vssd1 vssd1 vccd1 vccd1
+ _15571_/D sky130_fd_sc_hd__o221ai_4
XFILLER_15_823 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _16488_/A vssd1 vssd1 vccd1 vccd1 _15696_/D sky130_fd_sc_hd__buf_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16257__B _16257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14499_/Y _14607_/B _14492_/Y _14497_/Y vssd1 vssd1 vccd1 vccd1 _14522_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11733_ _15557_/A vssd1 vssd1 vccd1 vccd1 _18093_/C sky130_fd_sc_hd__buf_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17383__A2 _17388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _17133_/Y _17235_/Y _17237_/Y _17129_/Y vssd1 vssd1 vccd1 vccd1 _17242_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_30_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14443_/X _11404_/A _14448_/X vssd1 vssd1 vccd1 vccd1 _22667_/D sky130_fd_sc_hd__a21o_1
XFILLER_187_658 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _18459_/C _18666_/B _18839_/B _11664_/D vssd1 vssd1 vccd1 vccd1 _11932_/C
+ sky130_fd_sc_hd__and4_4
XFILLER_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13403_ _22851_/Q vssd1 vssd1 vccd1 vccd1 _21990_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_70_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17171_ _16966_/X _17164_/Y _17167_/Y _17170_/Y vssd1 vssd1 vccd1 vccd1 _17172_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14383_ _14383_/A vssd1 vssd1 vccd1 vccd1 _14593_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__13944__A2 _14181_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17135__A2 _15919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11595_ _15904_/A _15905_/A _18131_/B _18131_/C vssd1 vssd1 vccd1 vccd1 _11595_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11955__A1 _11285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16122_ _16070_/Y _16121_/X _16073_/Y _16076_/Y vssd1 vssd1 vccd1 vccd1 _16122_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_31_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13334_ _13450_/C vssd1 vssd1 vccd1 vccd1 _21713_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_127_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15697__A2 _15774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16894__A1 _16397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16053_ _11459_/A _11459_/B _11778_/A _11778_/B _12988_/A vssd1 vssd1 vccd1 vccd1
+ _16053_/X sky130_fd_sc_hd__a221o_4
XFILLER_155_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13265_ _13265_/A vssd1 vssd1 vccd1 vccd1 _21632_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater131_A _22846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20690__A2 _17833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15004_ _15114_/A _15064_/C _15070_/A _15004_/D vssd1 vssd1 vccd1 vccd1 _15013_/A
+ sky130_fd_sc_hd__and4_1
X_12216_ _18282_/A vssd1 vssd1 vccd1 vccd1 _12216_/X sky130_fd_sc_hd__buf_2
XFILLER_29_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18635__A2 _18627_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17816__B _17816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13196_ _13375_/A vssd1 vssd1 vccd1 vccd1 _13521_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_68_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15449__A2 _16274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16720__B _20781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19812_ _19763_/Y _19765_/Y _19817_/A vssd1 vssd1 vccd1 vccd1 _19823_/A sky130_fd_sc_hd__o21bai_2
XFILLER_97_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22441__C input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12147_ _22792_/Q _22793_/Q vssd1 vssd1 vccd1 vccd1 _18677_/A sky130_fd_sc_hd__nor2_4
XFILLER_110_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19743_ _19746_/A _19808_/B _19746_/C vssd1 vssd1 vccd1 vccd1 _19747_/A sky130_fd_sc_hd__a21oi_1
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16955_ _16225_/A _16227_/A _16947_/A _17144_/C vssd1 vssd1 vccd1 vccd1 _17138_/A
+ sky130_fd_sc_hd__o211ai_2
X_12078_ _11903_/B _11903_/C _11909_/C vssd1 vssd1 vccd1 vccd1 _12079_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13137__A _22843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15906_ _15904_/X _15905_/X _20502_/B vssd1 vssd1 vccd1 vccd1 _15906_/Y sky130_fd_sc_hd__o21ai_1
X_19674_ _19674_/A _19674_/B _22919_/Q vssd1 vssd1 vccd1 vccd1 _19827_/A sky130_fd_sc_hd__nand3_1
X_16886_ _17049_/A _16886_/B _17049_/B vssd1 vssd1 vccd1 vccd1 _17076_/C sky130_fd_sc_hd__nand3_4
XANTENNA__19060__A2 _18371_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12041__A _22660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11583__C _16313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18625_ _19043_/A _17391_/A _17647_/A _18636_/A vssd1 vssd1 vccd1 vccd1 _18625_/X
+ sky130_fd_sc_hd__o22a_1
X_15837_ _15828_/X _15826_/Y _15836_/X vssd1 vssd1 vccd1 vccd1 _15944_/A sky130_fd_sc_hd__a21o_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15621__A2 _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15352__A _15352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15768_ _15862_/A _15864_/D _15766_/X _15767_/X vssd1 vssd1 vccd1 vccd1 _15769_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_18556_ _18556_/A _18556_/B _18556_/C vssd1 vssd1 vccd1 vccd1 _18568_/B sky130_fd_sc_hd__nand3_2
XFILLER_75_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17507_ _17507_/A _17726_/D _17726_/C _17959_/C vssd1 vssd1 vccd1 vccd1 _17508_/C
+ sky130_fd_sc_hd__nand4_1
X_14719_ _13851_/A _13851_/B _13748_/X vssd1 vssd1 vccd1 vccd1 _14719_/X sky130_fd_sc_hd__a21o_1
XFILLER_75_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18487_ _18487_/A _18487_/B vssd1 vssd1 vccd1 vccd1 _18490_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15699_ _15748_/A vssd1 vssd1 vccd1 vccd1 _15740_/B sky130_fd_sc_hd__inv_2
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18663__A _18663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17438_ _17430_/Y _17437_/X _17433_/C vssd1 vssd1 vccd1 vccd1 _17449_/C sky130_fd_sc_hd__o21bai_2
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17369_ _17719_/A _17719_/C vssd1 vssd1 vccd1 vccd1 _22957_/D sky130_fd_sc_hd__xor2_2
XFILLER_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13935__A2 _13814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17126__A2 _17122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19197__C _19197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11946__A1 _18292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13022__D _13022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19108_ _19303_/A _19116_/A vssd1 vssd1 vccd1 vccd1 _19111_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20380_ _20240_/C _20240_/A _20240_/B _20398_/A vssd1 vssd1 vccd1 vccd1 _20380_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_119_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039_ _19034_/Y _18908_/A _19095_/C _18908_/B vssd1 vssd1 vccd1 vccd1 _19039_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_173_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput100 _14417_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_115_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput111 _14346_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[7] sky130_fd_sc_hd__buf_2
Xoutput122 _22670_/Q vssd1 vssd1 vccd1 vccd1 y[6] sky130_fd_sc_hd__buf_2
XFILLER_161_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22050_ _21964_/X _21970_/X _21957_/A _21972_/C vssd1 vssd1 vccd1 vccd1 _22099_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_86_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16630__B _16630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21001_ _20958_/A _20958_/B _22938_/Q vssd1 vssd1 vccd1 vccd1 _21001_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14431__A _14431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11774__B _11949_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22952_ _22952_/CLK _22952_/D vssd1 vssd1 vccd1 vccd1 _22952_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19051__A2 _12158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__C _18453_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21903_ _21802_/A _21792_/X _21802_/C _21901_/Y _21902_/Y vssd1 vssd1 vccd1 vccd1
+ _21909_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_44_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22883_ _22915_/CLK input77/X vssd1 vssd1 vccd1 vccd1 _22883_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16358__A _20471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21834_ _21834_/A _21834_/B _21834_/C _21834_/D vssd1 vssd1 vccd1 vccd1 _21931_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_55_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21697__A1 _21440_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_664 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21765_ _21765_/A vssd1 vssd1 vccd1 vccd1 _21846_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20716_ _20630_/A _20602_/Y _20634_/C vssd1 vssd1 vccd1 vccd1 _20721_/A sky130_fd_sc_hd__o21ai_1
XFILLER_184_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20608__A _20608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21696_ _21560_/A _21556_/A _21838_/A vssd1 vssd1 vccd1 vccd1 _21698_/B sky130_fd_sc_hd__a21o_1
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20647_ _20452_/A _20452_/B _20454_/C _20928_/C _20449_/Y vssd1 vssd1 vccd1 vccd1
+ _20648_/A sky130_fd_sc_hd__a41o_1
XFILLER_177_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11937__A1 _11704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20657__C1 _20551_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ _11380_/A _11380_/B vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__nand2_2
XANTENNA__11949__B _18680_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20578_ _12967_/A _17874_/A _17875_/A _20462_/A vssd1 vssd1 vccd1 vccd1 _20578_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_125_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14336__C1 _14335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22317_ _22317_/A _22317_/B vssd1 vssd1 vccd1 vccd1 _22318_/B sky130_fd_sc_hd__nor2_1
XFILLER_124_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13050_ _13176_/A vssd1 vssd1 vccd1 vccd1 _13050_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21439__A _22675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18617__A2 _12116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22248_ _22245_/X _22246_/Y _22155_/A _22212_/Y vssd1 vssd1 vccd1 vccd1 _22250_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12001_ _12001_/A _12001_/B vssd1 vssd1 vccd1 vccd1 _12001_/Y sky130_fd_sc_hd__nand2_2
XFILLER_3_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22179_ _22179_/A vssd1 vssd1 vccd1 vccd1 _22186_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17652__A _19585_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16740_ _16734_/X _16735_/X _16739_/Y vssd1 vssd1 vccd1 vccd1 _16740_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_115_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1000 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20188__A1 _20064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13952_ _13728_/A _22859_/D _13727_/A _13763_/A _22872_/Q vssd1 vssd1 vccd1 vccd1
+ _13954_/A sky130_fd_sc_hd__a32o_1
XFILLER_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _20133_/A vssd1 vssd1 vccd1 vccd1 _16129_/C sky130_fd_sc_hd__buf_2
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16671_ _16659_/B _16659_/C _16659_/A vssd1 vssd1 vccd1 vccd1 _16672_/A sky130_fd_sc_hd__a21oi_2
X_13883_ _14722_/A _13876_/A _14721_/B _14184_/C vssd1 vssd1 vccd1 vccd1 _13883_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_62_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16800__A1 _16177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18410_ _18401_/X _18403_/X _18406_/Y _18409_/Y vssd1 vssd1 vccd1 vccd1 _18411_/C
+ sky130_fd_sc_hd__o211ai_1
X_15622_ _11911_/A _16300_/A _12009_/A _15378_/A vssd1 vssd1 vccd1 vccd1 _15647_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_185_1047 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19390_ _19457_/A _19389_/B _19389_/C vssd1 vssd1 vccd1 vccd1 _19390_/Y sky130_fd_sc_hd__a21oi_1
X_12834_ _20213_/B vssd1 vssd1 vccd1 vccd1 _20092_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12417__A2 _12967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _18337_/X _18484_/A _18340_/Y vssd1 vssd1 vccd1 vccd1 _18349_/A sky130_fd_sc_hd__o21ai_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _19358_/A _19358_/B _15774_/D vssd1 vssd1 vccd1 vccd1 _16215_/B sky130_fd_sc_hd__and3_1
XANTENNA__13404__B _21990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _13022_/A vssd1 vssd1 vccd1 vccd1 _12765_/X sky130_fd_sc_hd__buf_2
XANTENNA__18483__A _18690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17356__A2 _17227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_612 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14818_/A _14057_/X _14503_/X _13924_/X vssd1 vssd1 vccd1 vccd1 _14504_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_70_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11716_ _15481_/A vssd1 vssd1 vccd1 vccd1 _22658_/B sky130_fd_sc_hd__buf_2
X_18272_ _18272_/A _18272_/B _18272_/C vssd1 vssd1 vccd1 vccd1 _18272_/Y sky130_fd_sc_hd__nand3_1
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19298__B _19298_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15484_ _15484_/A _15486_/B vssd1 vssd1 vccd1 vccd1 _15521_/A sky130_fd_sc_hd__nor2_1
XANTENNA__15367__B2 _15378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21621__B _21725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12921_/A vssd1 vssd1 vccd1 vccd1 _12696_/X sky130_fd_sc_hd__buf_4
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17223_ _17221_/Y _17222_/Y _17070_/B _17070_/A vssd1 vssd1 vccd1 vccd1 _17223_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_187_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14435_ _14439_/A _22967_/Q vssd1 vssd1 vccd1 vccd1 _14435_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11647_ _11647_/A _11647_/B _11647_/C _11647_/D vssd1 vssd1 vccd1 vccd1 _11689_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_128_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21340__C _21741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 wb_adr_i[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22851__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17154_ _16959_/B _16956_/Y _16948_/X _16946_/X vssd1 vssd1 vccd1 vccd1 _17155_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_156_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput24 wb_adr_i[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
X_14366_ _22764_/Q vssd1 vssd1 vccd1 vccd1 _14366_/X sky130_fd_sc_hd__clkbuf_4
Xinput35 wb_dat_i[0] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_4
XANTENNA__20112__A1 _12928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11578_ _11578_/A _11581_/A vssd1 vssd1 vccd1 vccd1 _11578_/Y sky130_fd_sc_hd__nor2_1
Xinput46 wb_dat_i[1] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__20112__B2 _20110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput57 wb_dat_i[2] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_4
X_16105_ _16069_/X _16099_/X _16104_/Y vssd1 vssd1 vccd1 vccd1 _16111_/A sky130_fd_sc_hd__o21ai_2
Xinput68 wb_we_i vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__20640__A2_N _20737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13317_ _21202_/A vssd1 vssd1 vccd1 vccd1 _13317_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput79 x[8] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17085_ _20584_/A _20584_/B _17085_/C vssd1 vssd1 vccd1 vccd1 _17085_/Y sky130_fd_sc_hd__nand3_4
XFILLER_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14297_ input25/X input24/X input32/X input31/X vssd1 vssd1 vccd1 vccd1 _14300_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_143_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16036_ _15949_/A _15947_/Y _15942_/X _15937_/X vssd1 vssd1 vccd1 vccd1 _16038_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13248_ _13273_/A vssd1 vssd1 vccd1 vccd1 _21250_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17277__D1 _20781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21612__A1 _21383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ _13105_/A _13105_/B _13120_/B _13120_/A vssd1 vssd1 vccd1 vccd1 _13216_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_35_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21571__A1_N _22674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17987_ _17987_/A _17987_/B vssd1 vssd1 vccd1 vccd1 _17988_/B sky130_fd_sc_hd__nor2_1
XFILLER_85_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12105__A1 _11771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18658__A _18797_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22168__A2 _13305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19726_ _19726_/A vssd1 vssd1 vccd1 vccd1 _19735_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16938_ _17133_/A _19490_/B _19490_/A vssd1 vssd1 vccd1 vccd1 _16976_/B sky130_fd_sc_hd__and3_2
XANTENNA__20179__A1 _12765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17281__B _17281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19657_ _19656_/Y _19652_/Y _19555_/C _19545_/Y vssd1 vssd1 vccd1 vccd1 _19658_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16869_ _16869_/A _16869_/B vssd1 vssd1 vccd1 vccd1 _16869_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16178__A _16178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16398__A3 _16400_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15082__A _15082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18608_ _18556_/B _18556_/C _18556_/A vssd1 vssd1 vccd1 vccd1 _18608_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_19_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19588_ _19588_/A vssd1 vssd1 vccd1 vccd1 _19596_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18539_ _18528_/X _18529_/Y _18535_/Y _18538_/X vssd1 vssd1 vccd1 vccd1 _18553_/A
+ sky130_fd_sc_hd__o2bb2ai_4
XANTENNA__18544__A1 _11979_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18544__B2 _11474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15810__A _15810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21550_ _21410_/B _21410_/C _21410_/A _21417_/B _21417_/C vssd1 vssd1 vccd1 vccd1
+ _21551_/B sky130_fd_sc_hd__a32o_2
XFILLER_194_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20501_ _20501_/A vssd1 vssd1 vccd1 vccd1 _20501_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21481_ _21490_/A _21481_/B vssd1 vssd1 vccd1 vccd1 _21504_/B sky130_fd_sc_hd__nand2_2
XFILLER_119_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11919__A1 _11606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20432_ _20549_/B _20432_/B _20549_/C _20549_/D vssd1 vssd1 vccd1 vccd1 _20554_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_146_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22643__A _22643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17737__A _18305_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16063__D _16586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20363_ _20224_/C _20224_/A _20224_/B vssd1 vssd1 vccd1 vccd1 _20363_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__11488__C _11980_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16641__A _20972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22102_ _22102_/A _22102_/B vssd1 vssd1 vccd1 vccd1 _22102_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13984__B _14564_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20294_ _20298_/A _20294_/B vssd1 vssd1 vccd1 vccd1 _20319_/A sky130_fd_sc_hd__nand2_1
XFILLER_115_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12344__A1 _16318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22033_ _21683_/A _21724_/D _21724_/A _22196_/A _22034_/C vssd1 vssd1 vccd1 vccd1
+ _22131_/A sky130_fd_sc_hd__a32o_2
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15833__A2 _17652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19024__A2 _17434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22935_ _22937_/CLK _22935_/D vssd1 vssd1 vccd1 vccd1 _22935_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15423__C _20129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22866_ _22916_/CLK _22866_/D vssd1 vssd1 vccd1 vccd1 _22866_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21817_ _21698_/B _21698_/C _21695_/C vssd1 vssd1 vccd1 vccd1 _21817_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_169_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22797_ _22797_/CLK _22797_/D vssd1 vssd1 vccd1 vccd1 _22797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22874__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ _12550_/A _12550_/B _12550_/C vssd1 vssd1 vccd1 vccd1 _12565_/A sky130_fd_sc_hd__nand3_2
XFILLER_196_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21748_ _21936_/A _21757_/A _21937_/A vssd1 vssd1 vccd1 vccd1 _21748_/Y sky130_fd_sc_hd__nand3_1
XFILLER_169_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11501_ _11381_/X _11636_/A _11500_/Y vssd1 vssd1 vccd1 vccd1 _11501_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_19_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22619__A0 _22798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ _12683_/A vssd1 vssd1 vccd1 vccd1 _20250_/C sky130_fd_sc_hd__buf_2
XFILLER_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21679_ _21648_/X _21657_/Y _21664_/X _21677_/X vssd1 vssd1 vccd1 vccd1 _21680_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_7_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14220_ _14917_/C _14276_/D _15118_/A _14220_/D vssd1 vssd1 vccd1 vccd1 _14256_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_156_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18299__B1 _18778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12032__B1 _11685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ _18663_/A vssd1 vssd1 vccd1 vccd1 _19061_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_149_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16849__A1 _16742_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_992 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21842__A1 _21269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ _14151_/A _14151_/B _14151_/C vssd1 vssd1 vccd1 vccd1 _14248_/A sky130_fd_sc_hd__nand3_2
XANTENNA__17647__A _17647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11363_ _11471_/C vssd1 vssd1 vccd1 vccd1 _11430_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_152_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16551__A _18680_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13102_ _13105_/A _13300_/A _13591_/A _13322_/A _21343_/A vssd1 vssd1 vccd1 vccd1
+ _13122_/B sky130_fd_sc_hd__o2111ai_4
XANTENNA__21169__A _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14082_ _14082_/A vssd1 vssd1 vccd1 vccd1 _14161_/B sky130_fd_sc_hd__clkbuf_1
X_11294_ _11325_/B _11404_/D vssd1 vssd1 vccd1 vccd1 _11295_/B sky130_fd_sc_hd__nand2_4
XFILLER_106_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17910_ _17910_/A _17910_/B _17910_/C _17910_/D vssd1 vssd1 vccd1 vccd1 _17910_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_117_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _13028_/Y _13029_/Y _13032_/X vssd1 vssd1 vccd1 vccd1 _13038_/B sky130_fd_sc_hd__o21ai_1
XFILLER_133_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18890_ _18890_/A vssd1 vssd1 vccd1 vccd1 _18890_/X sky130_fd_sc_hd__buf_2
XANTENNA__17085__C _17085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15809__C1 _11672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17841_ _17839_/X _17736_/B _19793_/C _18030_/B vssd1 vssd1 vccd1 vccd1 _17842_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14088__A1 _14147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18478__A _18765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12099__B1 _12098_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17772_ _17626_/X _17627_/X _17697_/C _17727_/X _17769_/Y vssd1 vssd1 vccd1 vccd1
+ _17776_/A sky130_fd_sc_hd__a311o_1
XANTENNA__19015__A2 _15808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14984_ _14980_/A _15035_/B _14980_/C vssd1 vssd1 vccd1 vccd1 _14984_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13835__A1 _13736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18197__B _19351_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19511_ _19511_/A _19511_/B _19580_/A vssd1 vssd1 vccd1 vccd1 _19581_/A sky130_fd_sc_hd__nand3_2
X_16723_ _16743_/A _16743_/C _16743_/B vssd1 vssd1 vccd1 vccd1 _16723_/X sky130_fd_sc_hd__a21o_2
X_13935_ _13814_/A _13814_/B _13926_/Y _14502_/A vssd1 vssd1 vccd1 vccd1 _13935_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17532__D _17532_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19442_ _19442_/A vssd1 vssd1 vccd1 vccd1 _19442_/Y sky130_fd_sc_hd__inv_2
X_16654_ _17076_/A _17076_/B vssd1 vssd1 vccd1 vccd1 _16659_/A sky130_fd_sc_hd__nand2_1
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13866_ _13830_/Y _13866_/B _13866_/C vssd1 vssd1 vccd1 vccd1 _13867_/A sky130_fd_sc_hd__nand3b_1
XFILLER_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15605_ _16319_/B _16318_/A _16319_/D _15370_/A vssd1 vssd1 vccd1 vccd1 _20461_/A
+ sky130_fd_sc_hd__o211ai_4
X_12817_ _12817_/A _12817_/B vssd1 vssd1 vccd1 vccd1 _12818_/C sky130_fd_sc_hd__nand2_1
X_19373_ _19190_/C _19372_/X _19190_/B vssd1 vssd1 vccd1 vccd1 _19376_/B sky130_fd_sc_hd__o21ai_1
X_16585_ _16585_/A _16585_/B vssd1 vssd1 vccd1 vccd1 _17313_/B sky130_fd_sc_hd__nand2_2
XFILLER_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13797_ _13959_/A _13989_/A _14506_/C vssd1 vssd1 vccd1 vccd1 _13808_/A sky130_fd_sc_hd__nand3_2
XFILLER_62_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15536_ _15536_/A vssd1 vssd1 vccd1 vccd1 _15536_/X sky130_fd_sc_hd__clkbuf_2
X_18324_ _18324_/A _22796_/Q vssd1 vssd1 vccd1 vccd1 _18495_/B sky130_fd_sc_hd__nand2_2
XFILLER_176_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _13007_/A vssd1 vssd1 vccd1 vccd1 _12749_/B sky130_fd_sc_hd__inv_2
XFILLER_148_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18255_ _18231_/Y _18234_/X _18250_/B vssd1 vssd1 vccd1 vccd1 _18257_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15467_ _15465_/X _15466_/Y _15306_/Y vssd1 vssd1 vccd1 vccd1 _15574_/C sky130_fd_sc_hd__o21ai_4
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12679_ _16257_/D vssd1 vssd1 vccd1 vccd1 _17401_/B sky130_fd_sc_hd__clkbuf_4
X_17206_ _17206_/A _17206_/B vssd1 vssd1 vccd1 vccd1 _17208_/C sky130_fd_sc_hd__nand2_1
XFILLER_147_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14418_ _22369_/D vssd1 vssd1 vccd1 vccd1 _14418_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18186_ _18395_/B _18395_/C vssd1 vssd1 vccd1 vccd1 _18187_/B sky130_fd_sc_hd__nand2_1
X_15398_ _15331_/Y _15329_/X _15426_/B _15344_/X vssd1 vssd1 vccd1 vccd1 _15513_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_156_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20097__B1 _12687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17137_ _17137_/A vssd1 vssd1 vccd1 vccd1 _17400_/A sky130_fd_sc_hd__buf_4
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14349_ _12107_/C _14338_/X _14339_/X _14331_/X _12378_/C vssd1 vssd1 vccd1 vccd1
+ _14349_/X sky130_fd_sc_hd__a32o_1
XFILLER_7_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16461__A _20086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17068_ _17222_/A _17222_/B _22895_/Q vssd1 vssd1 vccd1 vccd1 _17071_/B sky130_fd_sc_hd__a21o_1
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16019_ _16133_/A _16134_/B vssd1 vssd1 vccd1 vccd1 _16020_/B sky130_fd_sc_hd__nand2_1
XANTENNA__19772__A _19900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22402__S _22402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17292__A _19336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21349__B1 _13350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19709_ _19704_/Y _19789_/B _19709_/C vssd1 vssd1 vccd1 vccd1 _19864_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__19557__A3 _18023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20981_ _20982_/A _20982_/B _20982_/C vssd1 vssd1 vccd1 vccd1 _20985_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__17568__A2 _17412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22897__CLK _22952_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22720_ input33/X _22720_/D vssd1 vssd1 vccd1 vccd1 _22720_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15579__A1 _15465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16058__D _16100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22651_ _22651_/A vssd1 vssd1 vccd1 vccd1 _22812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19714__B1 _16016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19012__A _19687_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21602_ _21739_/C _21738_/A vssd1 vssd1 vccd1 vccd1 _22184_/A sky130_fd_sc_hd__and2_1
X_22582_ _22782_/Q input58/X _22584_/S vssd1 vssd1 vccd1 vccd1 _22583_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17029__A2_N _16740_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21533_ _21401_/Y _21390_/Y _21404_/Y _21403_/Y vssd1 vssd1 vccd1 vccd1 _21545_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_22_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17740__A2 _17817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21464_ _21805_/D _21514_/C _21666_/B vssd1 vssd1 vccd1 vccd1 _21464_/X sky130_fd_sc_hd__and3_1
XFILLER_182_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11368__A2 _18795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17467__A _17467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20415_ _20415_/A vssd1 vssd1 vccd1 vccd1 _20449_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_174_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21395_ _21179_/C _21179_/B _21179_/A vssd1 vssd1 vccd1 vccd1 _21395_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_107_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12107__C _12107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20605__B _20605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20346_ _20463_/A _20463_/B _20346_/C vssd1 vssd1 vccd1 vccd1 _20347_/B sky130_fd_sc_hd__and3_1
XFILLER_190_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20277_ _20284_/B vssd1 vssd1 vccd1 vccd1 _20281_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22016_ _22016_/A _22679_/Q vssd1 vssd1 vccd1 vccd1 _22016_/X sky130_fd_sc_hd__and2_1
XFILLER_89_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12123__B _12123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11540__A2 _18367_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15806__A2 _15810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17633__C _17833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17008__B2 _17728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11981_ _11526_/A _11979_/Y _11980_/X _11372_/A _18330_/A vssd1 vssd1 vccd1 vccd1
+ _11981_/X sky130_fd_sc_hd__o32a_1
XFILLER_57_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14490__A1 _14857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13720_ _13821_/B _13897_/A _13810_/C vssd1 vssd1 vccd1 vccd1 _14065_/A sky130_fd_sc_hd__o21ai_1
XFILLER_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_832 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22918_ _22922_/CLK _22918_/D vssd1 vssd1 vccd1 vccd1 _22918_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16231__A2 _12774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13651_ _13649_/X _21757_/A _13401_/A _13650_/X vssd1 vssd1 vccd1 vccd1 _13658_/C
+ sky130_fd_sc_hd__a31oi_1
XFILLER_44_567 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22849_ _22850_/CLK _22861_/Q vssd1 vssd1 vccd1 vccd1 _22849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15450__A _15450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12602_ _12445_/Y _12595_/Y _12436_/Y vssd1 vssd1 vccd1 vccd1 _12602_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_169_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16370_ _16377_/A _16370_/B _16377_/B _16377_/C vssd1 vssd1 vccd1 vccd1 _16370_/Y
+ sky130_fd_sc_hd__nand4_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_228 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13582_ _21588_/B vssd1 vssd1 vccd1 vccd1 _21195_/C sky130_fd_sc_hd__buf_2
XANTENNA__15990__A1 _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20068__A _20069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _20611_/A _16712_/C vssd1 vssd1 vccd1 vccd1 _15321_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _12540_/C vssd1 vssd1 vccd1 vccd1 _15776_/D sky130_fd_sc_hd__buf_2
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18040_ _18040_/A vssd1 vssd1 vccd1 vccd1 _18040_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15252_ _15252_/A _15262_/A vssd1 vssd1 vccd1 vccd1 _22685_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12464_ _12579_/C vssd1 vssd1 vccd1 vccd1 _20478_/C sky130_fd_sc_hd__buf_2
XFILLER_184_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14203_ _14203_/A _14203_/B _14785_/B _14786_/B vssd1 vssd1 vccd1 vccd1 _14203_/X
+ sky130_fd_sc_hd__and4_1
X_11415_ _11415_/A vssd1 vssd1 vccd1 vccd1 _11636_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__20618__A2 _17131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15183_ _15240_/A _14854_/X _15148_/A _15152_/C vssd1 vssd1 vccd1 vccd1 _15210_/A
+ sky130_fd_sc_hd__o31a_1
X_12395_ _12467_/A vssd1 vssd1 vccd1 vccd1 _15466_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_193_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12017__C _17312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16712__C _16712_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14134_ _13736_/B _13833_/X _14489_/C _14963_/A vssd1 vssd1 vccd1 vccd1 _14134_/Y
+ sky130_fd_sc_hd__o211ai_4
X_11346_ _12148_/A _11764_/B vssd1 vssd1 vccd1 vccd1 _11429_/A sky130_fd_sc_hd__nand2_2
X_19991_ _19991_/A _19991_/B vssd1 vssd1 vccd1 vccd1 _19992_/C sky130_fd_sc_hd__nor2_1
XFILLER_193_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18942_ _18933_/X _18646_/X _18927_/Y _18932_/Y vssd1 vssd1 vccd1 vccd1 _18945_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14702__C1 _22765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14065_ _14065_/A vssd1 vssd1 vccd1 vccd1 _14834_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11277_ _11277_/A vssd1 vssd1 vccd1 vccd1 _11420_/C sky130_fd_sc_hd__buf_2
X_13016_ _13024_/A _13024_/B _13016_/C _16153_/A vssd1 vssd1 vccd1 vccd1 _13016_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_140_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18873_ _18722_/D _18721_/B _18722_/C vssd1 vssd1 vccd1 vccd1 _18899_/A sky130_fd_sc_hd__a21boi_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17824_ _17886_/B _17824_/B vssd1 vssd1 vccd1 vccd1 _17826_/C sky130_fd_sc_hd__nand2_1
XANTENNA__17107__A1_N _16976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20250__B _20502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12968__B _12968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17755_ _17755_/A _17755_/B vssd1 vssd1 vccd1 vccd1 _17755_/Y sky130_fd_sc_hd__nor2_1
X_14967_ _14966_/A _14966_/C _14966_/B vssd1 vssd1 vccd1 vccd1 _14968_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__17840__A _17840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16706_ _16706_/A vssd1 vssd1 vccd1 vccd1 _16706_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13918_ _13984_/A vssd1 vssd1 vccd1 vccd1 _14808_/A sky130_fd_sc_hd__buf_2
X_17686_ _17687_/C _17687_/A _17687_/B vssd1 vssd1 vccd1 vccd1 _17688_/B sky130_fd_sc_hd__a21o_1
X_14898_ _14966_/A _14965_/A _14965_/B vssd1 vssd1 vccd1 vccd1 _14899_/B sky130_fd_sc_hd__and3_1
XFILLER_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19425_ _19419_/X _19418_/X _19556_/A _19422_/A vssd1 vssd1 vccd1 vccd1 _19427_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16637_ _16637_/A _16637_/B _16706_/A vssd1 vssd1 vccd1 vccd1 _16637_/Y sky130_fd_sc_hd__nand3_2
X_13849_ _13892_/B _13849_/B _13849_/C vssd1 vssd1 vccd1 vccd1 _13851_/A sky130_fd_sc_hd__nand3_4
XFILLER_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12984__A _15799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19356_ _19350_/X _15840_/A _19352_/X _19368_/B _19355_/Y vssd1 vssd1 vccd1 vccd1
+ _19356_/X sky130_fd_sc_hd__o311a_2
XFILLER_50_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21081__B _21081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16568_ _16568_/A vssd1 vssd1 vccd1 vccd1 _17875_/A sky130_fd_sc_hd__buf_2
XFILLER_149_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18307_ _18307_/A vssd1 vssd1 vccd1 vccd1 _18442_/B sky130_fd_sc_hd__clkbuf_1
X_15519_ _15738_/B vssd1 vssd1 vccd1 vccd1 _15859_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18093__D _18093_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19287_ _22916_/Q _19288_/B vssd1 vssd1 vccd1 vccd1 _19289_/A sky130_fd_sc_hd__nor2_1
XFILLER_149_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16499_ _15495_/X _15435_/D _11660_/A _16226_/B _18258_/B vssd1 vssd1 vccd1 vccd1
+ _16499_/X sky130_fd_sc_hd__o311a_1
XFILLER_31_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18238_ _18238_/A _18238_/B vssd1 vssd1 vccd1 vccd1 _18239_/C sky130_fd_sc_hd__nand2_1
XANTENNA__22059__B2 _22062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21806__A1 _22229_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18169_ _19470_/B _19504_/D _18363_/A _18130_/Y vssd1 vssd1 vccd1 vccd1 _18310_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16191__A _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20200_ _20200_/A _20199_/Y vssd1 vssd1 vccd1 vccd1 _20200_/X sky130_fd_sc_hd__or2b_1
XFILLER_143_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21180_ _21179_/C _21176_/A _21179_/A vssd1 vssd1 vccd1 vccd1 _21181_/B sky130_fd_sc_hd__a21o_1
XANTENNA__20085__A3 _20359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15497__B1 _12672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20131_ _12671_/A _12844_/A _20242_/A vssd1 vssd1 vccd1 vccd1 _20131_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_171_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20062_ _20049_/B _20061_/Y _20055_/Y vssd1 vssd1 vccd1 vccd1 _20063_/B sky130_fd_sc_hd__a21oi_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18986__A1 _15797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__A2 _18445_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16069__C _16106_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13055__A _13055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20964_ _20946_/A _20946_/B _20945_/B vssd1 vssd1 vccd1 vccd1 _21008_/A sky130_fd_sc_hd__o21a_2
XANTENNA__22368__A _22368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22703_ _22800_/CLK _22703_/D vssd1 vssd1 vccd1 vccd1 _22703_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20895_ _20842_/X _20892_/Y _20894_/Y vssd1 vssd1 vccd1 vccd1 _20906_/C sky130_fd_sc_hd__o21ai_4
XFILLER_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22634_ _22634_/A vssd1 vssd1 vccd1 vccd1 _22804_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__19699__C1 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15972__A1 _16241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15972__B2 _12774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19163__A1 _11636_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19163__B2 _15888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17174__B1 _17123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22565_ _22774_/Q input49/X _22569_/S vssd1 vssd1 vccd1 vccd1 _22566_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18910__A1 _19602_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21516_ _21507_/Y _21512_/Y _21514_/X _21515_/Y vssd1 vssd1 vccd1 vccd1 _21538_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_182_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22496_ _22496_/A vssd1 vssd1 vccd1 vccd1 _22743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22912__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21447_ _21990_/A _21629_/B _21990_/C vssd1 vssd1 vccd1 vccd1 _21633_/A sky130_fd_sc_hd__nand3_2
XFILLER_182_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19466__A2 _15808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12180_ _12164_/Y _12168_/X _18162_/A _18165_/A vssd1 vssd1 vccd1 vccd1 _12181_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_150_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21378_ _21378_/A _21378_/B vssd1 vssd1 vccd1 vccd1 _21393_/C sky130_fd_sc_hd__nor2_1
XFILLER_79_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20329_ _12721_/A _15718_/A _20210_/A _20210_/B vssd1 vssd1 vccd1 vccd1 _20364_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_62_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21025__A2 _17816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_924 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11513__A2 _18203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18459__C _18459_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15870_ _17039_/A _20806_/C _17816_/A _17039_/D vssd1 vssd1 vccd1 vccd1 _15870_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_114_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input22_A wb_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ _14821_/A _14821_/B vssd1 vssd1 vccd1 vccd1 _14822_/A sky130_fd_sc_hd__nor2_1
XFILLER_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _17539_/Y _17535_/Y _17533_/X vssd1 vssd1 vccd1 vccd1 _17540_/Y sky130_fd_sc_hd__a21oi_1
X_14752_ _14752_/A _14752_/B _14839_/A _14839_/B vssd1 vssd1 vccd1 vccd1 _14752_/X
+ sky130_fd_sc_hd__and4_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _11964_/A _11964_/B _11964_/C vssd1 vssd1 vccd1 vccd1 _11964_/X sky130_fd_sc_hd__and3_1
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12474__B1 _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20536__A1 _20844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _22753_/Q vssd1 vssd1 vccd1 vccd1 _13707_/A sky130_fd_sc_hd__buf_2
X_17471_ _17469_/A _17469_/B _17479_/A _17479_/B vssd1 vssd1 vccd1 vccd1 _17474_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_567 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14683_ _14684_/A _14693_/B _14684_/C vssd1 vssd1 vccd1 vccd1 _14793_/A sky130_fd_sc_hd__nand3_1
XFILLER_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11895_ _11895_/A _11895_/B _11895_/C vssd1 vssd1 vccd1 vccd1 _11896_/B sky130_fd_sc_hd__nand3_1
X_19210_ _19037_/A _19031_/X _19037_/B vssd1 vssd1 vccd1 vccd1 _19210_/Y sky130_fd_sc_hd__a21boi_1
X_16422_ _16422_/A _16657_/C vssd1 vssd1 vccd1 vccd1 _16422_/Y sky130_fd_sc_hd__nand2_1
X_13634_ _13361_/X _13319_/X _13126_/X _13434_/X vssd1 vssd1 vccd1 vccd1 _13634_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_60_846 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15963__B2 _15962_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12777__A1 _12765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19141_ _22915_/Q _19141_/B _19141_/C vssd1 vssd1 vccd1 vccd1 _19142_/B sky130_fd_sc_hd__nand3b_1
X_16353_ _16345_/X _16352_/Y _16310_/Y _16315_/X vssd1 vssd1 vccd1 vccd1 _16355_/B
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__19587__A _19587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13565_ _13523_/C _13565_/B _13565_/C vssd1 vssd1 vccd1 vccd1 _13565_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_34_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15304_ _15454_/A _15304_/B vssd1 vssd1 vccd1 vccd1 _15304_/Y sky130_fd_sc_hd__nand2_1
X_19072_ _11380_/A _11380_/B _18830_/D _19046_/A _19065_/A vssd1 vssd1 vccd1 vccd1
+ _19074_/C sky130_fd_sc_hd__a32o_1
XFILLER_157_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12516_ _12525_/A _12525_/B _20123_/A vssd1 vssd1 vccd1 vccd1 _12516_/X sky130_fd_sc_hd__a21o_1
X_16284_ _16287_/A _16287_/B _16286_/A vssd1 vssd1 vccd1 vccd1 _16606_/C sky130_fd_sc_hd__and3_1
XANTENNA__15715__A1 _16554_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13496_ _13556_/C _13496_/B vssd1 vssd1 vccd1 vccd1 _13498_/C sky130_fd_sc_hd__nand2_1
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18023_ _18023_/A vssd1 vssd1 vccd1 vccd1 _18023_/X sky130_fd_sc_hd__clkbuf_2
X_15235_ _15223_/Y _15242_/A _15227_/A _15225_/Y vssd1 vssd1 vccd1 vccd1 _15245_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12447_ _12447_/A vssd1 vssd1 vccd1 vccd1 _16257_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_172_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17468__A1 _17466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16125__D1 _12876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15166_ _15112_/A _15112_/B _15111_/B vssd1 vssd1 vccd1 vccd1 _15168_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__15339__B _15339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12378_ _12378_/A _12378_/B _12378_/C vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__nand3_2
XFILLER_125_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _14117_/A _14785_/B _14786_/B _14203_/A vssd1 vssd1 vccd1 vccd1 _14117_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_140_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11329_ _11420_/B _11302_/A _11860_/A _11277_/A vssd1 vssd1 vccd1 vccd1 _11371_/B
+ sky130_fd_sc_hd__o211ai_2
X_19974_ _19974_/A _19974_/B _19974_/C vssd1 vssd1 vccd1 vccd1 _19974_/Y sky130_fd_sc_hd__nand3_1
XFILLER_158_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15097_ _15097_/A _15097_/B vssd1 vssd1 vccd1 vccd1 _15098_/C sky130_fd_sc_hd__and2_1
XANTENNA__15058__C _15058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18925_ _18929_/A _18929_/B _18978_/A _18931_/B vssd1 vssd1 vccd1 vccd1 _18937_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__16691__A2 _16670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14048_ _14099_/B _14099_/C _14096_/C vssd1 vssd1 vccd1 vccd1 _14097_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20261__A _20261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15355__A _15355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18856_ _18856_/A vssd1 vssd1 vccd1 vccd1 _19695_/A sky130_fd_sc_hd__buf_2
XFILLER_121_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17640__A1 _15840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17807_ _17833_/B vssd1 vssd1 vccd1 vccd1 _21017_/A sky130_fd_sc_hd__buf_2
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18787_ _18969_/A _18969_/B _18788_/A vssd1 vssd1 vccd1 vccd1 _18970_/B sky130_fd_sc_hd__o21ai_1
XFILLER_95_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15999_ _15780_/B _15901_/Y _17085_/C _15900_/Y _15577_/D vssd1 vssd1 vccd1 vccd1
+ _16000_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_94_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17738_ _19689_/C vssd1 vssd1 vccd1 vccd1 _19769_/B sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_2_0_bq_clk_i_A clkbuf_4_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18196__A2 _15531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17669_ _16124_/X _17006_/A _17562_/Y _17564_/Y vssd1 vssd1 vccd1 vccd1 _17669_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19408_ _19408_/A vssd1 vssd1 vccd1 vccd1 _19408_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12217__B1 _11818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1078 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20680_ _17423_/X _17424_/X _12721_/X vssd1 vssd1 vccd1 vccd1 _20680_/X sky130_fd_sc_hd__a21o_1
XANTENNA__22935__CLK _22937_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19339_ _19326_/A _19512_/A _19512_/B vssd1 vssd1 vccd1 vccd1 _19342_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__12219__A _12219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22350_ _22341_/B _22338_/A _22338_/B _22352_/A vssd1 vssd1 vccd1 vccd1 _22354_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21301_ _21301_/A vssd1 vssd1 vccd1 vccd1 _21466_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22281_ _22244_/B _22280_/Y _22277_/X _22317_/A vssd1 vssd1 vccd1 vccd1 _22282_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14434__A _22964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21232_ _21238_/C _21238_/B _21226_/Y _21227_/X vssd1 vssd1 vccd1 vccd1 _21239_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_145_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11777__B _15714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11743__A2 _11721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21163_ _21164_/A _21164_/B _21161_/X _21162_/Y vssd1 vssd1 vccd1 vccd1 _21167_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20114_ _12810_/B _12810_/C _12810_/A _12859_/A _12859_/B vssd1 vssd1 vccd1 vccd1
+ _20115_/C sky130_fd_sc_hd__a32oi_4
X_21094_ _21138_/A _21094_/B vssd1 vssd1 vccd1 vccd1 _21094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_120_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20045_ _20042_/Y _20044_/Y _20025_/X _20032_/B vssd1 vssd1 vccd1 vccd1 _20059_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19620__A2 _20012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1120 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21996_ _21996_/A _21996_/B _21996_/C _21996_/D vssd1 vssd1 vccd1 vccd1 _21996_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__21715__B1 _21269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19384__A1 _19340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _20884_/A _20884_/B _20884_/C _20882_/B _20882_/A vssd1 vssd1 vccd1 vccd1
+ _20949_/A sky130_fd_sc_hd__o32a_1
XFILLER_26_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _15484_/A vssd1 vssd1 vccd1 vccd1 _14438_/A sky130_fd_sc_hd__buf_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20878_ _20941_/A _20879_/C _20879_/A vssd1 vssd1 vccd1 vccd1 _20880_/A sky130_fd_sc_hd__a21o_1
X_22617_ _18698_/A input39/X _22619_/S vssd1 vssd1 vccd1 vccd1 _22618_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16824__A _19320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18344__C1 _19587_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13350_ _13350_/A vssd1 vssd1 vccd1 vccd1 _21767_/A sky130_fd_sc_hd__buf_2
XFILLER_14_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18895__B1 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22548_ _22548_/A vssd1 vssd1 vccd1 vccd1 _22766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12301_ _12437_/A vssd1 vssd1 vccd1 vccd1 _20130_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13281_ _13281_/A _13281_/B vssd1 vssd1 vccd1 vccd1 _13413_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14344__A _14370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22479_ _22479_/A vssd1 vssd1 vccd1 vccd1 _22735_/D sky130_fd_sc_hd__clkbuf_1
X_15020_ _14959_/C _14960_/B _15018_/X _15019_/Y vssd1 vssd1 vccd1 vccd1 _15088_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_154_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12232_ _22658_/B _12046_/X _12043_/A _11721_/C vssd1 vssd1 vccd1 vccd1 _15445_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_136_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21246__A2 _21247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18111__A2 _18849_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12931__A1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _18093_/A _18093_/B _15714_/A vssd1 vssd1 vccd1 vccd1 _12163_/X sky130_fd_sc_hd__and3_2
XANTENNA__12931__B2 _16155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16971_ _16971_/A _16971_/B vssd1 vssd1 vccd1 vccd1 _16972_/B sky130_fd_sc_hd__nand2_1
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12094_ _12094_/A _19358_/D _19358_/C _12094_/D vssd1 vssd1 vccd1 vccd1 _12094_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_7_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20206__B1 _20086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18710_ _18905_/A _18905_/B _18722_/C _18722_/D vssd1 vssd1 vccd1 vccd1 _18713_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_122_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15922_ _15915_/A _15915_/B _15920_/X _15921_/X vssd1 vssd1 vccd1 vccd1 _15967_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_19690_ _12207_/X _19839_/D _19500_/X vssd1 vssd1 vccd1 vccd1 _19690_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12695__B1 _20584_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18641_ _18619_/Y _18624_/A _18633_/Y vssd1 vssd1 vccd1 vccd1 _18933_/A sky130_fd_sc_hd__a21o_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15853_ _15853_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15855_/B sky130_fd_sc_hd__nor2_1
XFILLER_49_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15402__A1_N _12094_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18486__A _18706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14804_ _14716_/C _14800_/X _14716_/B vssd1 vssd1 vccd1 vccd1 _14806_/B sky130_fd_sc_hd__o21ai_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18572_ _18572_/A _18572_/B _18572_/C vssd1 vssd1 vccd1 vccd1 _18572_/X sky130_fd_sc_hd__and3_1
XANTENNA__20509__A1 _16778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ _15915_/B vssd1 vssd1 vccd1 vccd1 _15784_/Y sky130_fd_sc_hd__inv_2
X_12996_ _12994_/X _12990_/A _13036_/A vssd1 vssd1 vccd1 vccd1 _12996_/X sky130_fd_sc_hd__a21o_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22958__CLK _22964_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17523_ _17523_/A _17523_/B _17523_/C vssd1 vssd1 vccd1 vccd1 _17585_/B sky130_fd_sc_hd__and3_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11947_ _11947_/A _11947_/B _11947_/C vssd1 vssd1 vccd1 vccd1 _12219_/A sky130_fd_sc_hd__nand3_4
XFILLER_17_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14735_ _14733_/A _14733_/B _14737_/A _14737_/B vssd1 vssd1 vccd1 vccd1 _14735_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13423__A _13423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17454_ _17454_/A _17454_/B _17454_/C vssd1 vssd1 vccd1 vccd1 _17479_/A sky130_fd_sc_hd__nand3_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _15176_/A vssd1 vssd1 vccd1 vccd1 _14845_/B sky130_fd_sc_hd__clkbuf_2
X_11878_ _18679_/C vssd1 vssd1 vccd1 vccd1 _18258_/A sky130_fd_sc_hd__buf_4
XFILLER_189_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16405_ _16433_/A _16433_/B _16433_/C vssd1 vssd1 vccd1 vccd1 _16406_/B sky130_fd_sc_hd__and3_1
X_13617_ _13617_/A _13617_/B _13617_/C vssd1 vssd1 vccd1 vccd1 _13617_/X sky130_fd_sc_hd__and3_1
XFILLER_189_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17385_ _19772_/C _17385_/B _17385_/C _17525_/D vssd1 vssd1 vccd1 vccd1 _17385_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14597_ _14576_/X _14578_/A _14575_/A vssd1 vssd1 vccd1 vccd1 _14600_/A sky130_fd_sc_hd__o21ai_1
XFILLER_9_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19124_ _19121_/B _19122_/Y _19123_/Y vssd1 vssd1 vccd1 vccd1 _19124_/X sky130_fd_sc_hd__a21o_1
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16336_ _15567_/A _15565_/B _15565_/C _15565_/D vssd1 vssd1 vccd1 vccd1 _16336_/Y
+ sky130_fd_sc_hd__a22oi_2
X_13548_ _13548_/A vssd1 vssd1 vccd1 vccd1 _13614_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_146_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18350__A2 _18135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11973__A2 _11639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19055_ _18330_/X _18203_/C _18797_/Y vssd1 vssd1 vccd1 vccd1 _19055_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16267_ _16267_/A vssd1 vssd1 vccd1 vccd1 _16267_/X sky130_fd_sc_hd__clkbuf_2
X_13479_ _13484_/A _13484_/B _13289_/A vssd1 vssd1 vccd1 vccd1 _13479_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18006_ _18055_/A _18055_/B _22905_/Q vssd1 vssd1 vccd1 vccd1 _18015_/C sky130_fd_sc_hd__a21o_1
XFILLER_145_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15218_ _15185_/B _15240_/A _15214_/X _15217_/X vssd1 vssd1 vccd1 vccd1 _15224_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18638__B1 _18619_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16198_ _16043_/A _16043_/B _16043_/C vssd1 vssd1 vccd1 vccd1 _16198_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _15149_/A vssd1 vssd1 vccd1 vccd1 _15217_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19957_ _19860_/Y _19863_/Y _19916_/A _19917_/A _19956_/X vssd1 vssd1 vccd1 vccd1
+ _19959_/B sky130_fd_sc_hd__o32ai_4
XANTENNA__14675__A1 _14670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15872__B1 _16034_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18908_ _18908_/A _18908_/B _18908_/C vssd1 vssd1 vccd1 vccd1 _18914_/B sky130_fd_sc_hd__nand3_2
XFILLER_19_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19888_ _19890_/A _19887_/B _19887_/C vssd1 vssd1 vccd1 vccd1 _19889_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18839_ _19194_/A _18839_/B _19465_/A _19194_/D vssd1 vssd1 vccd1 vccd1 _18839_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_83_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21850_ _21850_/A _22108_/C _22031_/A _22106_/A vssd1 vssd1 vccd1 vccd1 _21850_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18169__A2 _19504_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20801_ _20711_/Y _20718_/X _20720_/C vssd1 vssd1 vccd1 vccd1 _20803_/A sky130_fd_sc_hd__o21ai_1
XFILLER_24_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21781_ _21781_/A _21781_/B _21781_/C vssd1 vssd1 vccd1 vccd1 _21802_/C sky130_fd_sc_hd__nand3_2
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14429__A _14429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20732_ _20818_/B _20730_/B _20778_/B _20812_/A vssd1 vssd1 vccd1 vccd1 _20737_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20663_ _20827_/B _20827_/C _21066_/A _20827_/A vssd1 vssd1 vccd1 vccd1 _20768_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__18326__C1 _15415_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_698 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22402_ _22702_/Q input40/X _22402_/S vssd1 vssd1 vccd1 vccd1 _22403_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11413__A1 _15482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20594_ _20596_/A _20702_/A _20595_/A _20682_/B vssd1 vssd1 vccd1 vccd1 _20629_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22333_ _22333_/A _22333_/B vssd1 vssd1 vccd1 vccd1 _22335_/A sky130_fd_sc_hd__nor2_1
XANTENNA__16352__A1 _16103_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22264_ _22231_/D _22263_/B _22263_/C vssd1 vssd1 vccd1 vccd1 _22264_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21215_ _21724_/A _21609_/B _21724_/D vssd1 vssd1 vccd1 vccd1 _21216_/B sky130_fd_sc_hd__nand3_2
XFILLER_133_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22195_ _22195_/A _22195_/B vssd1 vssd1 vccd1 vccd1 _22215_/A sky130_fd_sc_hd__xor2_2
XFILLER_160_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21146_ _22945_/Q _21157_/B vssd1 vssd1 vccd1 vccd1 _21151_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15707__B _15707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13508__A _22041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12412__A _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21077_ _21076_/C _21075_/Y _21004_/B _21076_/Y vssd1 vssd1 vccd1 vccd1 _21124_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_76_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20028_ _20042_/B _20029_/B _20029_/C vssd1 vssd1 vccd1 vccd1 _20032_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__18801__B1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16819__A _18848_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15615__B1 _16304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17080__A2 _16579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ _20120_/A _12859_/A _12859_/B vssd1 vssd1 vccd1 vccd1 _12851_/B sky130_fd_sc_hd__a21o_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15723__A _15723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11801_ _11800_/X _11639_/A _11797_/A vssd1 vssd1 vccd1 vccd1 _11964_/A sky130_fd_sc_hd__o21ai_1
XFILLER_61_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _12886_/B _12781_/B _16160_/C _20452_/C vssd1 vssd1 vccd1 vccd1 _12781_/X
+ sky130_fd_sc_hd__and4b_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ _21934_/Y _21935_/Y _21977_/Y _21978_/X vssd1 vssd1 vccd1 vccd1 _22029_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14492_/Y _14611_/B _14497_/Y vssd1 vssd1 vccd1 vccd1 _14522_/A sky130_fd_sc_hd__a21o_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11732_/A vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__buf_4
XANTENNA__16257__C _16257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20911__A1 _20123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14443_/X _11404_/D _14448_/X vssd1 vssd1 vccd1 vccd1 _22666_/D sky130_fd_sc_hd__a21o_1
XFILLER_159_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _19322_/A vssd1 vssd1 vccd1 vccd1 _18839_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18317__C1 _22796_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13402_ _13664_/B vssd1 vssd1 vccd1 vccd1 _13659_/C sky130_fd_sc_hd__buf_2
X_17170_ _17170_/A _17180_/A vssd1 vssd1 vccd1 vccd1 _17170_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14382_ _22442_/B vssd1 vssd1 vccd1 vccd1 _14382_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17369__B _17719_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11594_ _11594_/A vssd1 vssd1 vccd1 vccd1 _15905_/A sky130_fd_sc_hd__buf_2
XANTENNA__13944__A3 _14181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16121_ _16081_/A _16081_/B _16056_/Y vssd1 vssd1 vccd1 vccd1 _16121_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11955__A2 _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13333_ _13450_/A vssd1 vssd1 vccd1 vccd1 _21713_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16052_ _16047_/A _16047_/B _16050_/Y _16051_/X vssd1 vssd1 vccd1 vccd1 _16126_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_183_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16894__A2 _15630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13264_ _21398_/B _21367_/C _13517_/C vssd1 vssd1 vccd1 vccd1 _13272_/B sky130_fd_sc_hd__nand3_1
XANTENNA__20690__A3 _17833_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15003_ _15062_/A vssd1 vssd1 vccd1 vccd1 _15114_/A sky130_fd_sc_hd__buf_2
X_12215_ _17380_/A _17381_/A _18445_/A vssd1 vssd1 vccd1 vccd1 _18282_/A sky130_fd_sc_hd__o21ai_2
XFILLER_29_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17385__A _19772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13195_ _13143_/A _13143_/B _13112_/D _21473_/A vssd1 vssd1 vccd1 vccd1 _13375_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_29_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19811_ _19811_/A _19833_/A vssd1 vssd1 vccd1 vccd1 _19817_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16720__C _16720_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15303__C1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ _12146_/A _12146_/B vssd1 vssd1 vccd1 vccd1 _12146_/Y sky130_fd_sc_hd__nand2_2
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19742_ _19742_/A _19742_/B _19808_/A vssd1 vssd1 vccd1 vccd1 _19808_/B sky130_fd_sc_hd__nand3_2
XFILLER_173_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16954_ _16954_/A _16954_/B vssd1 vssd1 vccd1 vccd1 _16954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12077_ _12075_/Y _12076_/X _12077_/C _12077_/D vssd1 vssd1 vccd1 vccd1 _12079_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15905_ _15905_/A vssd1 vssd1 vccd1 vccd1 _15905_/X sky130_fd_sc_hd__buf_4
X_19673_ _19674_/A _19674_/B _22919_/Q vssd1 vssd1 vccd1 vccd1 _19675_/A sky130_fd_sc_hd__a21o_1
XFILLER_37_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16885_ _16884_/X _16885_/B _17042_/A vssd1 vssd1 vccd1 vccd1 _17049_/B sky130_fd_sc_hd__nand3b_2
XANTENNA__11583__D _18875_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18624_ _18624_/A vssd1 vssd1 vccd1 vccd1 _18835_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15633__A _15633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _15915_/A _15914_/A _16414_/B _15784_/Y vssd1 vssd1 vccd1 vccd1 _15836_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_65_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18555_ _18557_/B _18555_/B vssd1 vssd1 vccd1 vccd1 _18556_/C sky130_fd_sc_hd__nand2_2
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _15860_/A _15860_/B _15758_/C vssd1 vssd1 vccd1 vccd1 _15767_/X sky130_fd_sc_hd__a21o_1
X_12979_ _12981_/D _15899_/B _20134_/B _12981_/B _12981_/C vssd1 vssd1 vccd1 vccd1
+ _12982_/A sky130_fd_sc_hd__a32o_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17506_ _17502_/X _17910_/D _17853_/A vssd1 vssd1 vccd1 vccd1 _17508_/A sky130_fd_sc_hd__o21ai_1
XFILLER_17_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14718_ _15114_/C _15114_/D _14727_/A _14494_/D _14623_/X vssd1 vssd1 vccd1 vccd1
+ _14731_/A sky130_fd_sc_hd__a41o_1
X_18486_ _18706_/A _18691_/A _18691_/B vssd1 vssd1 vccd1 vccd1 _18487_/B sky130_fd_sc_hd__and3_1
XFILLER_61_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15698_ _15698_/A _15698_/B _15698_/C vssd1 vssd1 vccd1 vccd1 _15748_/A sky130_fd_sc_hd__nand3_2
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22466__A _22512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17437_ _17442_/A _17440_/A _17277_/Y _17431_/D _17436_/X vssd1 vssd1 vccd1 vccd1
+ _17437_/X sky130_fd_sc_hd__o311a_1
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14649_ _14638_/Y _14649_/B _14649_/C vssd1 vssd1 vccd1 vccd1 _14656_/C sky130_fd_sc_hd__nand3b_1
XFILLER_21_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17368_ _22896_/Q _17220_/B _17367_/Y _17223_/Y vssd1 vssd1 vccd1 vccd1 _17719_/C
+ sky130_fd_sc_hd__o22ai_4
XFILLER_146_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17126__A3 _17122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19197__D _19197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19107_ _19257_/A _19257_/B _19257_/C vssd1 vssd1 vccd1 vccd1 _19116_/A sky130_fd_sc_hd__nand3_2
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16319_ _16319_/A _16319_/B _16319_/C _16319_/D vssd1 vssd1 vccd1 vccd1 _16320_/B
+ sky130_fd_sc_hd__nand4_4
X_17299_ _17299_/A _17299_/B _17299_/C vssd1 vssd1 vccd1 vccd1 _17307_/C sky130_fd_sc_hd__nand3_1
XFILLER_173_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19038_ _19035_/X _19037_/X _19004_/Y _19010_/X vssd1 vssd1 vccd1 vccd1 _19095_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_134_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput101 _14420_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput112 _14348_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[8] sky130_fd_sc_hd__buf_2
Xoutput123 _22671_/Q vssd1 vssd1 vccd1 vccd1 y[7] sky130_fd_sc_hd__buf_2
XFILLER_115_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15808__A _15808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21000_ _21076_/A _21076_/B vssd1 vssd1 vccd1 vccd1 _21004_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19036__B1 _19012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19941__C _19981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22951_ _22951_/CLK _22951_/D vssd1 vssd1 vccd1 vccd1 _22951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11493__D _16078_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22591__A0 _11395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21902_ _21933_/A _21902_/B vssd1 vssd1 vccd1 vccd1 _21902_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11882__A1 _16564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22882_ _22916_/CLK input76/X vssd1 vssd1 vccd1 vccd1 _22882_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19339__A1 _19326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16270__B1 _16269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_716 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21833_ _21922_/A _21831_/B _21922_/B _21832_/X vssd1 vssd1 vccd1 vccd1 _22934_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18854__A _18854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21764_ _21846_/A _21765_/A _21846_/C _21846_/D vssd1 vssd1 vccd1 vccd1 _21789_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__21697__A2 _21415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_676 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20715_ _20630_/A _20602_/Y _20634_/C _20710_/Y _20714_/Y vssd1 vssd1 vccd1 vccd1
+ _20778_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_169_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21695_ _21695_/A _21917_/B _21695_/C vssd1 vssd1 vccd1 vccd1 _21815_/B sky130_fd_sc_hd__nand3_2
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20646_ _20870_/C vssd1 vssd1 vccd1 vccd1 _20928_/C sky130_fd_sc_hd__buf_2
XANTENNA__11937__A2 _11705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11949__C _19197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20577_ _20587_/B _20577_/B vssd1 vssd1 vccd1 vccd1 _20577_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11311__A _11404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22316_ _22316_/A _22316_/B vssd1 vssd1 vccd1 vccd1 _22318_/A sky130_fd_sc_hd__or2_1
XANTENNA__14336__B1 _14313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15718__A _15718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22247_ _22336_/A _22212_/Y _22245_/X _22246_/Y vssd1 vssd1 vccd1 vccd1 _22250_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_133_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12000_ _12135_/B _12154_/C _12135_/A vssd1 vssd1 vccd1 vccd1 _12001_/B sky130_fd_sc_hd__nand3_2
XFILLER_133_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22178_ _22238_/B _22178_/B vssd1 vssd1 vccd1 vccd1 _22193_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21129_ _21129_/A vssd1 vssd1 vccd1 vccd1 _22923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17652__B _17652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13951_ _13948_/X _13949_/X _13950_/X vssd1 vssd1 vccd1 vccd1 _13951_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20188__A2 _13045_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12902_ _20130_/A vssd1 vssd1 vccd1 vccd1 _20133_/A sky130_fd_sc_hd__clkbuf_4
X_16670_ _16670_/A vssd1 vssd1 vccd1 vccd1 _17227_/A sky130_fd_sc_hd__buf_2
XFILLER_19_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13882_ _13820_/X _13821_/Y _13823_/Y vssd1 vssd1 vccd1 vccd1 _14721_/B sky130_fd_sc_hd__a21oi_4
XFILLER_98_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16800__A2 _16799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15621_ _15792_/B _16737_/A _15616_/X _16397_/A vssd1 vssd1 vccd1 vccd1 _15621_/X
+ sky130_fd_sc_hd__o22a_1
X_12833_ _12824_/A _16320_/A _12519_/B _22698_/Q vssd1 vssd1 vccd1 vccd1 _20213_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18340_ _18340_/A _18340_/B vssd1 vssd1 vccd1 vccd1 _18340_/Y sky130_fd_sc_hd__nand2_2
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _16477_/B vssd1 vssd1 vccd1 vccd1 _19358_/B sky130_fd_sc_hd__clkbuf_4
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12651_/A _12651_/B _12651_/C _12763_/X vssd1 vssd1 vccd1 vccd1 _12764_/Y
+ sky130_fd_sc_hd__a31oi_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18483__B _18483_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _22961_/Q vssd1 vssd1 vccd1 vccd1 _15481_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14503_ _14503_/A vssd1 vssd1 vccd1 vccd1 _14503_/X sky130_fd_sc_hd__buf_2
XFILLER_188_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15483_ _22964_/Q vssd1 vssd1 vccd1 vccd1 _15486_/B sky130_fd_sc_hd__inv_2
X_18271_ _12241_/C _12241_/A _12241_/B vssd1 vssd1 vccd1 vccd1 _18271_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21621__C _21621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_624 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12592_/A _12592_/B _20584_/C _12588_/Y _16937_/B vssd1 vssd1 vccd1 vccd1
+ _12737_/A sky130_fd_sc_hd__o2111ai_4
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17222_ _17222_/A _17222_/B vssd1 vssd1 vccd1 vccd1 _17222_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14434_ _22964_/Q vssd1 vssd1 vccd1 vccd1 _14439_/A sky130_fd_sc_hd__clkbuf_2
X_11646_ _11551_/B _11551_/C _11645_/Y _11536_/A vssd1 vssd1 vccd1 vccd1 _11646_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_156_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput14 wb_adr_i[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__22101__A3 _21725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17153_ _17138_/X _17142_/X _17145_/Y _16937_/B _19504_/B vssd1 vssd1 vccd1 vccd1
+ _17155_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__16316__A1 _15988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 wb_adr_i[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_2
X_14365_ _22732_/Q vssd1 vssd1 vccd1 vccd1 _21307_/B sky130_fd_sc_hd__clkbuf_2
Xinput36 wb_dat_i[10] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__14532__D_N _14273_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20112__A2 _16039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ _11840_/A _11577_/B vssd1 vssd1 vccd1 vccd1 _11696_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12317__A _22818_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput47 wb_dat_i[20] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16104_ _16113_/C _16150_/B vssd1 vssd1 vccd1 vccd1 _16104_/Y sky130_fd_sc_hd__nand2_1
X_13316_ _13316_/A vssd1 vssd1 vccd1 vccd1 _13316_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput58 wb_dat_i[30] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17084_ _11636_/X _17874_/A _17875_/A _16737_/X _17083_/X vssd1 vssd1 vccd1 vccd1
+ _17084_/X sky130_fd_sc_hd__o32a_1
Xinput69 x[0] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14296_ input3/X input2/X input5/X input4/X vssd1 vssd1 vccd1 vccd1 _14300_/A sky130_fd_sc_hd__or4_1
XFILLER_183_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16035_ _16035_/A _16035_/B _16035_/C vssd1 vssd1 vccd1 vccd1 _16657_/C sky130_fd_sc_hd__nand3_4
X_13247_ _13421_/A vssd1 vssd1 vccd1 vccd1 _21724_/C sky130_fd_sc_hd__buf_2
XANTENNA__15628__A _20471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17277__C1 _20781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16450__C _16450_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15347__B _16450_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ _13120_/A _13120_/B _13105_/Y _13216_/A vssd1 vssd1 vccd1 vccd1 _13181_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_96_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13148__A _22844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _11770_/X _11980_/B _11771_/X vssd1 vssd1 vccd1 vccd1 _18512_/B sky130_fd_sc_hd__a21oi_4
XFILLER_112_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17986_ _18030_/A _18030_/B _18030_/C _18030_/D vssd1 vssd1 vccd1 vccd1 _17987_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__12052__A _12052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19725_ _19725_/A _19725_/B _19725_/C vssd1 vssd1 vccd1 vccd1 _19726_/A sky130_fd_sc_hd__nand3_1
X_16937_ _19694_/B _16937_/B _17128_/B _19496_/A vssd1 vssd1 vccd1 vccd1 _16937_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_133_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20179__A2 _20843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__A _18629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19656_ _19740_/A _19656_/B vssd1 vssd1 vccd1 vccd1 _19656_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16868_ _16873_/C _16873_/D vssd1 vssd1 vccd1 vccd1 _16869_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17281__C _20678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18607_ _18960_/B _18960_/C vssd1 vssd1 vccd1 vccd1 _18607_/Y sky130_fd_sc_hd__nand2_1
X_15819_ _15886_/A _15819_/B _15819_/C vssd1 vssd1 vccd1 vccd1 _15828_/A sky130_fd_sc_hd__nand3_1
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19587_ _19587_/A _19587_/B _19587_/C _19587_/D vssd1 vssd1 vccd1 vccd1 _19588_/A
+ sky130_fd_sc_hd__nand4_1
X_16799_ _17379_/A vssd1 vssd1 vccd1 vccd1 _16799_/X sky130_fd_sc_hd__buf_4
XFILLER_18_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18538_ _16921_/X _18371_/A _18536_/Y _18537_/X _18531_/A vssd1 vssd1 vccd1 vccd1
+ _18538_/X sky130_fd_sc_hd__o221a_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18544__A2 _11980_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18469_ _18770_/C _18461_/B _18474_/A vssd1 vssd1 vccd1 vccd1 _18469_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__15810__B _15810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22676__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20500_ _20500_/A _20500_/B _20500_/C vssd1 vssd1 vccd1 vccd1 _20501_/A sky130_fd_sc_hd__nand3_1
XFILLER_193_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21480_ _21480_/A _21480_/B _22229_/C vssd1 vssd1 vccd1 vccd1 _21481_/B sky130_fd_sc_hd__and3_1
XFILLER_148_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20639__B1 _20734_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20431_ _20423_/C _20431_/B _20431_/C vssd1 vssd1 vccd1 vccd1 _20549_/C sky130_fd_sc_hd__nand3b_2
XFILLER_147_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20362_ _20366_/B _20366_/C _20366_/A vssd1 vssd1 vccd1 vccd1 _20362_/Y sky130_fd_sc_hd__a21oi_2
X_22101_ _21683_/A _21725_/A _21725_/B _22102_/A _22102_/B vssd1 vssd1 vccd1 vccd1
+ _22129_/A sky130_fd_sc_hd__a32o_1
XANTENNA__14442__A _22662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20293_ _20293_/A _20293_/B vssd1 vssd1 vccd1 vccd1 _20319_/B sky130_fd_sc_hd__nor2_2
XFILLER_115_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22032_ _22031_/A _21522_/D _22031_/C _22031_/B vssd1 vssd1 vccd1 vccd1 _22034_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18849__A _19504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13058__A _22735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15878__A1_N _16209_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16369__A _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22934_ _22937_/CLK _22934_/D vssd1 vssd1 vccd1 vccd1 _22934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_768 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22865_ _22944_/CLK _22877_/Q vssd1 vssd1 vccd1 vccd1 _22865_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15423__D _15774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21816_ _21837_/A vssd1 vssd1 vccd1 vccd1 _21816_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22796_ _22799_/CLK _22796_/D vssd1 vssd1 vccd1 vccd1 _22796_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_24_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21747_ _21874_/C _21596_/B _21591_/Y vssd1 vssd1 vccd1 vccd1 _21753_/B sky130_fd_sc_hd__a21o_1
XFILLER_185_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11500_ _18131_/B _18131_/C _18507_/C vssd1 vssd1 vccd1 vccd1 _11500_/Y sky130_fd_sc_hd__nand3_1
XFILLER_40_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22619__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14557__B1 _14552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12480_ _12456_/Y _12463_/Y _12478_/Y _12479_/X vssd1 vssd1 vccd1 vccd1 _12480_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_184_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21678_ _21664_/A _21674_/Y _21677_/X vssd1 vssd1 vccd1 vccd1 _21680_/A sky130_fd_sc_hd__a21o_1
XFILLER_156_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18299__A1 _15538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11431_ _11431_/A _11431_/B vssd1 vssd1 vccd1 vccd1 _18663_/A sky130_fd_sc_hd__nand2_4
XANTENNA__17928__A _17928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12032__A1 _11762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20629_ _20629_/A _20629_/B _20629_/C _20702_/B vssd1 vssd1 vccd1 vccd1 _20634_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14150_ _14147_/A _14147_/B _14148_/Y _14149_/X vssd1 vssd1 vccd1 vccd1 _14151_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11362_ _22787_/Q _22786_/Q _22784_/Q _11374_/A vssd1 vssd1 vccd1 vccd1 _18116_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_125_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21842__A2 _21341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16551__B _20092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ _13101_/A _13101_/B vssd1 vssd1 vccd1 vccd1 _21343_/A sky130_fd_sc_hd__nand2_1
XFILLER_192_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14081_ _14082_/A _14083_/A _14149_/B vssd1 vssd1 vccd1 vccd1 _14147_/C sky130_fd_sc_hd__a21o_1
X_11293_ _22955_/Q vssd1 vssd1 vccd1 vccd1 _11404_/D sky130_fd_sc_hd__buf_4
XANTENNA__21169__B _22852_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13032_ _13028_/Y _13029_/Y _13031_/Y vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__a21o_1
XANTENNA_input52_A wb_dat_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14071__B _14686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15809__B1 _14432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17840_ _17840_/A vssd1 vssd1 vccd1 vccd1 _18030_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12099__A1 _12117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21185__A _21185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17771_ _17785_/A vssd1 vssd1 vccd1 vccd1 _17777_/C sky130_fd_sc_hd__inv_2
X_14983_ _14923_/B _14923_/A _14981_/X _14982_/Y vssd1 vssd1 vccd1 vccd1 _15047_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_102_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13835__A2 _13833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19510_ _19511_/B _19580_/A _19511_/A vssd1 vssd1 vccd1 vccd1 _19510_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18197__C _18197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16722_ _16312_/X _16714_/X _16721_/X vssd1 vssd1 vccd1 vccd1 _16743_/B sky130_fd_sc_hd__o21ai_2
X_13934_ _13926_/Y _13927_/X _13931_/X _13933_/X vssd1 vssd1 vccd1 vccd1 _13937_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19441_ _19293_/X _19294_/X _19301_/Y _19440_/X vssd1 vssd1 vccd1 vccd1 _19442_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ _16653_/A _16653_/B _16653_/C vssd1 vssd1 vccd1 vccd1 _17076_/B sky130_fd_sc_hd__nand3_2
X_13865_ _13865_/A _13873_/A _14808_/C vssd1 vssd1 vccd1 vccd1 _13866_/C sky130_fd_sc_hd__nand3_1
XFILLER_16_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15604_ _22700_/Q vssd1 vssd1 vccd1 vccd1 _16319_/D sky130_fd_sc_hd__inv_2
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19372_ _18158_/X _18995_/B _19171_/Y _19174_/Y vssd1 vssd1 vccd1 vccd1 _19372_/X
+ sky130_fd_sc_hd__o211a_1
X_12816_ _20089_/A _20089_/B _22818_/Q vssd1 vssd1 vccd1 vccd1 _12817_/B sky130_fd_sc_hd__and3_1
XFILLER_188_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15993__C1 _20452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16584_ _16584_/A vssd1 vssd1 vccd1 vccd1 _16585_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_16_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13796_ _13963_/A _13833_/B _13833_/C _13821_/B vssd1 vssd1 vccd1 vccd1 _14506_/C
+ sky130_fd_sc_hd__a211o_2
XANTENNA__14260__A2 _14181_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18323_ _11770_/X _18313_/Y _18679_/C _18678_/C vssd1 vssd1 vccd1 vccd1 _18495_/A
+ sky130_fd_sc_hd__o211ai_4
X_15535_ _16481_/D vssd1 vssd1 vccd1 vccd1 _16241_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__15630__B _16431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12732_/Y _12744_/Y _12745_/Y _12746_/X vssd1 vssd1 vccd1 vccd1 _12896_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__17734__B1 _17928_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13431__A _22846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _18772_/B _18772_/C _18250_/B vssd1 vssd1 vccd1 vccd1 _18598_/B sky130_fd_sc_hd__a21oi_1
XFILLER_129_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15466_ _15557_/A _15466_/B _15466_/C vssd1 vssd1 vccd1 vccd1 _15466_/Y sky130_fd_sc_hd__nand3_2
X_12678_ _16256_/D vssd1 vssd1 vccd1 vccd1 _16257_/D sky130_fd_sc_hd__buf_2
XFILLER_169_990 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17205_ _17205_/A _17205_/B _17205_/C vssd1 vssd1 vccd1 vccd1 _17206_/B sky130_fd_sc_hd__nand3_1
X_11629_ _11625_/X _11626_/X _17312_/A _11614_/Y _11623_/X vssd1 vssd1 vccd1 vccd1
+ _11647_/D sky130_fd_sc_hd__o2111ai_4
XANTENNA__12023__A1 _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14417_ _22714_/Q _14403_/X _14410_/X _22746_/Q _14416_/X vssd1 vssd1 vccd1 vccd1
+ _14417_/X sky130_fd_sc_hd__a221o_1
XANTENNA__19487__B1 _19340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18185_ _18278_/B _18278_/A _18279_/A vssd1 vssd1 vccd1 vccd1 _18395_/C sky130_fd_sc_hd__nand3b_1
XANTENNA__17838__A _21011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13220__B1 _21757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15397_ _15396_/Y _15344_/X _15426_/B vssd1 vssd1 vccd1 vccd1 _15397_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_11_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20097__A1 _12577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17136_ _12735_/X _16758_/A _16946_/X _16948_/X vssd1 vssd1 vccd1 vccd1 _17136_/X
+ sky130_fd_sc_hd__o22a_1
X_14348_ _12343_/B _14344_/X _14337_/X _13301_/X _14347_/X vssd1 vssd1 vccd1 vccd1
+ _14348_/X sky130_fd_sc_hd__a221o_1
XFILLER_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17501__A3 _17959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15358__A _15377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17067_ _17222_/B _22895_/Q _17222_/A vssd1 vssd1 vccd1 vccd1 _17071_/A sky130_fd_sc_hd__nand3_1
X_14279_ _14279_/A _14279_/B _14279_/C _14279_/D vssd1 vssd1 vccd1 vccd1 _14280_/C
+ sky130_fd_sc_hd__nand4_1
X_16018_ _15812_/C _15812_/D _16017_/X vssd1 vssd1 vccd1 vccd1 _16134_/B sky130_fd_sc_hd__a21oi_2
XFILLER_170_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19772__B _19772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21597__A1 _13662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17969_ _17970_/B _22903_/Q vssd1 vssd1 vccd1 vccd1 _17969_/Y sky130_fd_sc_hd__nand2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_510 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19708_ _19708_/A _19708_/B _19789_/A vssd1 vssd1 vccd1 vccd1 _19789_/B sky130_fd_sc_hd__nand3_1
X_20980_ _20980_/A _20980_/B vssd1 vssd1 vccd1 vccd1 _20982_/C sky130_fd_sc_hd__xnor2_1
XFILLER_84_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19639_ _19538_/B _19538_/C _19538_/A vssd1 vssd1 vccd1 vccd1 _19649_/B sky130_fd_sc_hd__a21bo_1
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16240__A3 _15486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15821__A _18648_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22650_ _22812_/Q input55/X _22652_/S vssd1 vssd1 vccd1 vccd1 _22651_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19714__A1 _17442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21601_ _13633_/A _21594_/Y _21587_/Y _21589_/Y vssd1 vssd1 vccd1 vccd1 _21604_/B
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__19714__B2 _19838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19012__B _19351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22581_ _22581_/A vssd1 vssd1 vccd1 vccd1 _22781_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14437__A _22965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13979__C _14191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21532_ _21531_/A _21531_/C _21531_/B vssd1 vssd1 vccd1 vccd1 _21545_/A sky130_fd_sc_hd__a21o_1
XFILLER_138_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17748__A _17833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21463_ _21463_/A vssd1 vssd1 vccd1 vccd1 _21666_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20414_ _20843_/A _20429_/B _20281_/B vssd1 vssd1 vccd1 vccd1 _20414_/X sky130_fd_sc_hd__o21a_1
XFILLER_105_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21394_ _21404_/A _21404_/B _21403_/A vssd1 vssd1 vccd1 vccd1 _21394_/Y sky130_fd_sc_hd__nand3_1
XFILLER_179_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11773__B1 _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20345_ _20343_/A _20342_/A _20339_/Y vssd1 vssd1 vccd1 vccd1 _20347_/A sky130_fd_sc_hd__o21ai_1
XFILLER_88_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20276_ _12500_/X _12501_/X _20275_/Y _20390_/B _20155_/A vssd1 vssd1 vccd1 vccd1
+ _20284_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_955 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22015_ _22155_/A _22145_/A _22086_/A _22086_/B vssd1 vssd1 vccd1 vccd1 _22016_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15267__A1 _14990_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12123__C _12123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15806__A3 _16106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__A3 _16058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17633__D _19774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_1_bq_clk_i clkbuf_1_1_1_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22841__CLK _22937_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12420__A _15335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ _11980_/A _11980_/B _11980_/C vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__and3_1
XFILLER_112_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21733__A _21733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22917_ _22922_/CLK _22917_/D vssd1 vssd1 vccd1 vccd1 _22917_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__17964__B1 _17502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_844 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13650_ _13650_/A _13650_/B _21195_/B _21195_/C vssd1 vssd1 vccd1 vccd1 _13650_/X
+ sky130_fd_sc_hd__and4_1
X_22848_ _22943_/CLK hold19/X vssd1 vssd1 vccd1 vccd1 _22848_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12601_/A _12601_/B _12601_/C vssd1 vssd1 vccd1 vccd1 _12601_/Y sky130_fd_sc_hd__nand3_4
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _13581_/A vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22779_ _22813_/CLK _22779_/D vssd1 vssd1 vccd1 vccd1 _22779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15990__A2 _16324_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12793__C _22825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15320_ _15320_/A vssd1 vssd1 vccd1 vccd1 _20611_/A sky130_fd_sc_hd__buf_2
X_12532_ _12532_/A vssd1 vssd1 vccd1 vccd1 _20134_/A sky130_fd_sc_hd__buf_2
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_bq_clk_i clkbuf_4_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _22929_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19469__B1 _18514_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15251_ _15180_/B _15233_/A _15180_/A _15205_/C _14551_/A vssd1 vssd1 vccd1 vccd1
+ _15262_/A sky130_fd_sc_hd__a41o_1
X_12463_ _12441_/Y _12460_/Y _12462_/Y vssd1 vssd1 vccd1 vccd1 _12463_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_32_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16562__A _16751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11414_ _11756_/A vssd1 vssd1 vccd1 vccd1 _11415_/A sky130_fd_sc_hd__clkbuf_4
X_14202_ _14259_/A _14259_/B _14131_/X _14201_/X _14157_/A vssd1 vssd1 vccd1 vccd1
+ _14261_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_137_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15182_ _15182_/A vssd1 vssd1 vccd1 vccd1 _15240_/A sky130_fd_sc_hd__clkbuf_2
X_12394_ _12396_/A _12324_/X _12396_/C vssd1 vssd1 vccd1 vccd1 _12467_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20618__A3 _20917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14133_ _14237_/A _14237_/B _14237_/C vssd1 vssd1 vccd1 vccd1 _14238_/B sky130_fd_sc_hd__nand3_2
X_11345_ _12090_/A vssd1 vssd1 vccd1 vccd1 _11345_/X sky130_fd_sc_hd__buf_2
X_19990_ _19988_/X _20037_/B vssd1 vssd1 vccd1 vccd1 _19992_/B sky130_fd_sc_hd__and2b_1
XFILLER_125_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18692__A1 _18890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18941_ _18941_/A _18941_/B _18941_/C vssd1 vssd1 vccd1 vccd1 _18952_/A sky130_fd_sc_hd__nand3_1
XFILLER_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14064_ _14126_/A vssd1 vssd1 vccd1 vccd1 _14510_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11276_ _22787_/Q vssd1 vssd1 vccd1 vccd1 _11277_/A sky130_fd_sc_hd__inv_2
XFILLER_140_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12314__B _16256_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13015_ _13037_/B _13037_/A vssd1 vssd1 vccd1 vccd1 _13038_/A sky130_fd_sc_hd__or2_1
X_18872_ _19091_/B _18920_/B _18871_/Y vssd1 vssd1 vccd1 vccd1 _18908_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__16455__B1 _15450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17823_ _17886_/A _17821_/C _17928_/D _19839_/B vssd1 vssd1 vccd1 vccd1 _17824_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_66_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22528__A0 _13815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20250__C _20250_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12968__C _20697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17754_ _17755_/A _17755_/B _17746_/X _17753_/Y vssd1 vssd1 vccd1 vccd1 _17760_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_181_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14966_ _14966_/A _14966_/B _14966_/C vssd1 vssd1 vccd1 vccd1 _14968_/A sky130_fd_sc_hd__and3_1
XFILLER_48_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12330__A _22818_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19944__A1 _19981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16207__B1 _16034_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16705_ _16606_/X _16704_/Y _16620_/C _16620_/A vssd1 vssd1 vccd1 vccd1 _16705_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_63_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13917_ _13879_/X _13886_/Y _14021_/C _13916_/Y vssd1 vssd1 vccd1 vccd1 _13917_/Y
+ sky130_fd_sc_hd__o211ai_2
X_17685_ _17627_/A _17581_/B _17628_/A _17580_/Y vssd1 vssd1 vccd1 vccd1 _17688_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__16737__A _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14897_ _14966_/A _14965_/A _14965_/B vssd1 vssd1 vccd1 vccd1 _14899_/A sky130_fd_sc_hd__a21oi_1
X_19424_ _19424_/A _19424_/B vssd1 vssd1 vccd1 vccd1 _19427_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16636_ _16636_/A _16636_/B vssd1 vssd1 vccd1 vccd1 _16636_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13848_ _13848_/A vssd1 vssd1 vccd1 vccd1 _14061_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_90_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19355_ _16940_/X _18718_/X _19357_/B vssd1 vssd1 vccd1 vccd1 _19355_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16567_ _16324_/B _16324_/C _14369_/X vssd1 vssd1 vccd1 vccd1 _16568_/A sky130_fd_sc_hd__a21oi_2
XFILLER_149_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20306__A2 _20195_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ _22873_/Q vssd1 vssd1 vccd1 vccd1 _14613_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19172__A2 _19167_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18306_ _18572_/A _18572_/B _18572_/C vssd1 vssd1 vccd1 vccd1 _18307_/A sky130_fd_sc_hd__nand3_1
X_15518_ _15510_/B _15510_/C _15516_/Y _15517_/Y vssd1 vssd1 vccd1 vccd1 _15738_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_176_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19286_ _19286_/A _19286_/B vssd1 vssd1 vccd1 vccd1 _19288_/B sky130_fd_sc_hd__nand2_1
XFILLER_175_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16498_ _16498_/A _17646_/A _16498_/C _16498_/D vssd1 vssd1 vccd1 vccd1 _16498_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_148_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18237_ _11832_/Y _11834_/Y _11838_/Y _11927_/Y vssd1 vssd1 vccd1 vccd1 _18240_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_175_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15449_ _12929_/A _16274_/A _12117_/A _15455_/A vssd1 vssd1 vccd1 vccd1 _15449_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_50_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18168_ _19199_/A vssd1 vssd1 vccd1 vccd1 _19504_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_117_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21806__A2 _13630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17119_ _19012_/C _21019_/A _21019_/B vssd1 vssd1 vccd1 vccd1 _17120_/B sky130_fd_sc_hd__and3_1
XFILLER_190_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18683__A1 _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18099_ _18099_/A vssd1 vssd1 vccd1 vccd1 _18841_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16694__B1 _22890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20130_ _20130_/A _20130_/B _20130_/C vssd1 vssd1 vccd1 vccd1 _20242_/A sky130_fd_sc_hd__nand3_1
XFILLER_89_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11507__B1 _11504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20061_ _20034_/B _20058_/Y _20059_/Y _20060_/Y vssd1 vssd1 vccd1 vccd1 _20061_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_98_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22864__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18986__A2 _19160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11522__A3 _15624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22519__A0 _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12240__A _12240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18199__B1 _19047_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20963_ _20963_/A _20963_/B vssd1 vssd1 vccd1 vccd1 _22918_/D sky130_fd_sc_hd__xnor2_2
XANTENNA__16647__A _17039_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22702_ _22735_/CLK _22702_/D vssd1 vssd1 vccd1 vccd1 _22702_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20894_ _20894_/A _20894_/B _20894_/C vssd1 vssd1 vccd1 vccd1 _20894_/Y sky130_fd_sc_hd__nand3_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22633_ _22804_/Q input47/X _22641_/S vssd1 vssd1 vccd1 vccd1 _22634_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15972__A2 _11988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19163__A2 _19517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13071__A _22842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22564_ _22564_/A vssd1 vssd1 vccd1 vccd1 _22773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18910__A2 _19334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21515_ _21666_/A _21514_/C _21666_/B vssd1 vssd1 vccd1 vccd1 _21515_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22495_ _22743_/Q input50/X _22497_/S vssd1 vssd1 vccd1 vccd1 _22496_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21446_ _21393_/B _21393_/C _21393_/A vssd1 vssd1 vccd1 vccd1 _21538_/A sky130_fd_sc_hd__a21boi_1
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21377_ _21376_/X _13343_/X _13366_/Y _21179_/B _21374_/Y vssd1 vssd1 vccd1 vccd1
+ _21378_/B sky130_fd_sc_hd__o311a_2
XFILLER_123_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16741__B1_N _16842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20328_ _20446_/A _20446_/B _20328_/C _20328_/D vssd1 vssd1 vccd1 vccd1 _20335_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_162_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21447__B _21629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20259_ _20252_/Y _20261_/A _20263_/B vssd1 vssd1 vccd1 vccd1 _20260_/A sky130_fd_sc_hd__o21bai_2
XFILLER_135_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14820_ _14822_/C _14902_/A _14821_/A _14821_/B vssd1 vssd1 vccd1 vccd1 _14825_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_92_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_800 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input15_A wb_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12474__A1 _12470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ _14751_/A _14751_/B vssd1 vssd1 vccd1 vccd1 _14839_/B sky130_fd_sc_hd__or2_1
XFILLER_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ _11963_/A _12219_/B vssd1 vssd1 vccd1 vccd1 _12054_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17398__D1 _19768_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20536__A2 _16179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13702_ _13733_/B vssd1 vssd1 vccd1 vccd1 _13849_/C sky130_fd_sc_hd__buf_2
X_17470_ _17470_/A _17470_/B vssd1 vssd1 vccd1 vccd1 _17474_/A sky130_fd_sc_hd__nand2_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _14998_/A _14568_/A _14467_/X _14576_/X _14942_/B vssd1 vssd1 vccd1 vccd1
+ _14682_/X sky130_fd_sc_hd__o32a_1
XFILLER_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11894_ _11894_/A _11894_/B _11894_/C vssd1 vssd1 vccd1 vccd1 _11896_/A sky130_fd_sc_hd__nand3_1
XFILLER_189_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16421_ _16422_/A _16657_/C _16421_/C _16421_/D vssd1 vssd1 vccd1 vccd1 _16424_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__15180__B _15180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13633_ _13633_/A _13633_/B _13633_/C vssd1 vssd1 vccd1 vccd1 _13657_/C sky130_fd_sc_hd__or3_1
XFILLER_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19140_ _19141_/B _19141_/C _22915_/Q vssd1 vssd1 vccd1 vccd1 _19290_/A sky130_fd_sc_hd__a21bo_2
XFILLER_160_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16352_ _16103_/D _21011_/C _17462_/A _16316_/Y _16351_/X vssd1 vssd1 vccd1 vccd1
+ _16352_/Y sky130_fd_sc_hd__a311oi_4
XANTENNA__19587__B _19587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17165__A1 _19694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13564_ _13563_/A _13563_/B _13563_/C vssd1 vssd1 vccd1 vccd1 _13565_/C sky130_fd_sc_hd__a21o_1
XFILLER_185_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15303_ _11705_/X _11704_/X _12500_/X _12501_/X _11707_/A vssd1 vssd1 vccd1 vccd1
+ _15304_/B sky130_fd_sc_hd__o221a_1
XANTENNA__17388__A _17388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19071_ _19074_/A _19074_/B _19044_/X _19046_/X vssd1 vssd1 vccd1 vccd1 _19148_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_12515_ _12515_/A _22824_/Q vssd1 vssd1 vccd1 vccd1 _20123_/A sky130_fd_sc_hd__nand2_1
X_16283_ _16283_/A _16283_/B _16540_/A _16288_/C vssd1 vssd1 vccd1 vccd1 _16606_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_40_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13495_ _13495_/A _13495_/B _13495_/C vssd1 vssd1 vccd1 vccd1 _13498_/B sky130_fd_sc_hd__nand3_1
XFILLER_157_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15715__A2 _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18022_ _17946_/A _17996_/A _17994_/B vssd1 vssd1 vccd1 vccd1 _18036_/A sky130_fd_sc_hd__o21bai_1
XFILLER_157_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15234_ _15209_/A _15209_/B _15231_/B vssd1 vssd1 vccd1 vccd1 _15247_/A sky130_fd_sc_hd__o21a_1
X_12446_ _12436_/Y _12441_/Y _12445_/Y vssd1 vssd1 vccd1 vccd1 _12454_/A sky130_fd_sc_hd__o21ai_1
XFILLER_139_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1020 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16125__C1 _16124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15165_ _15162_/Y _15163_/X _15129_/A _15145_/Y vssd1 vssd1 vccd1 vccd1 _15168_/C
+ sky130_fd_sc_hd__a211oi_1
X_12377_ _12377_/A vssd1 vssd1 vccd1 vccd1 _12378_/B sky130_fd_sc_hd__buf_4
XFILLER_176_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22887__CLK _22952_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15339__C _15339_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14116_ _14200_/A vssd1 vssd1 vccd1 vccd1 _14785_/B sky130_fd_sc_hd__buf_2
X_11328_ _11306_/A _11385_/C _11374_/A _11619_/B _11860_/C vssd1 vssd1 vccd1 vccd1
+ _11371_/A sky130_fd_sc_hd__o311ai_4
X_19973_ _19973_/A _19975_/A vssd1 vssd1 vccd1 vccd1 _19974_/A sky130_fd_sc_hd__nor2_1
XFILLER_141_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15096_ _15095_/A _15093_/A _15095_/C vssd1 vssd1 vccd1 vccd1 _15097_/B sky130_fd_sc_hd__a21o_1
XFILLER_153_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18924_ _18977_/A vssd1 vssd1 vccd1 vccd1 _18931_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14047_ _14098_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14096_/C sky130_fd_sc_hd__xor2_2
XFILLER_80_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18855_ _18855_/A vssd1 vssd1 vccd1 vccd1 _18856_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15355__B _15355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15636__D1 _20678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17806_ _20975_/B _19901_/D _17872_/C _17806_/D vssd1 vssd1 vccd1 vccd1 _17895_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_83_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17640__A2 _17440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18786_ _22913_/Q vssd1 vssd1 vccd1 vccd1 _18788_/A sky130_fd_sc_hd__inv_2
X_15998_ _15997_/X _16005_/A _15900_/B _15983_/Y vssd1 vssd1 vccd1 vccd1 _16000_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__14454__A2 _15435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18666__B _18666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17737_ _18305_/C vssd1 vssd1 vccd1 vccd1 _17929_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ _15006_/B _15058_/A _15058_/B _14889_/A _15010_/C vssd1 vssd1 vccd1 vccd1
+ _14951_/C sky130_fd_sc_hd__a32o_1
XFILLER_78_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15371__A _17423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17668_ _17666_/X _17667_/Y _17665_/C vssd1 vssd1 vccd1 vccd1 _17687_/A sky130_fd_sc_hd__o21bai_2
XFILLER_91_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19407_ _19407_/A vssd1 vssd1 vccd1 vccd1 _19407_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16619_ _16624_/A _16624_/B _16619_/C vssd1 vssd1 vccd1 vccd1 _16620_/C sky130_fd_sc_hd__nand3_2
XANTENNA__12217__A1 _12204_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16617__D _16617_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17599_ _17600_/B _17600_/C _17600_/A vssd1 vssd1 vccd1 vccd1 _17781_/A sky130_fd_sc_hd__o21ai_1
XFILLER_195_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11404__A _11404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19338_ _19340_/A _19340_/B _19332_/Y _19337_/Y vssd1 vssd1 vccd1 vccd1 _19338_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__21488__B1 _21874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19269_ _19122_/B _19122_/C _19122_/A vssd1 vssd1 vccd1 vccd1 _19269_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14509__A3 _13815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21300_ _21266_/B _21266_/A _21265_/Y vssd1 vssd1 vccd1 vccd1 _21406_/A sky130_fd_sc_hd__a21o_1
XFILLER_176_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22280_ _22213_/Y _22216_/Y _22259_/X vssd1 vssd1 vccd1 vccd1 _22280_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_163_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21231_ _21231_/A vssd1 vssd1 vccd1 vccd1 _21247_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18656__A1 _15358_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11777__C _19496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16930__A _16930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21162_ _21162_/A _21162_/B vssd1 vssd1 vccd1 vccd1 _21162_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20452__A _20452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20113_ _20119_/A _20119_/B _20111_/X _20112_/X vssd1 vssd1 vccd1 vccd1 _20115_/B
+ sky130_fd_sc_hd__o2bb2ai_4
XANTENNA__15546__A _15546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21093_ _21093_/A _21092_/A vssd1 vssd1 vccd1 vccd1 _21094_/B sky130_fd_sc_hd__or2b_1
XFILLER_172_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20044_ _20022_/A _20043_/Y _20042_/C vssd1 vssd1 vccd1 vccd1 _20044_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_105_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input7_A wb_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19620__A3 _20012_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21283__A _21422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21995_ _21987_/Y _21989_/Y _22075_/B _22072_/A _22029_/A vssd1 vssd1 vccd1 vccd1
+ _21996_/D sky130_fd_sc_hd__o2111ai_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19384__A2 _19340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ _20946_/A _20946_/B vssd1 vssd1 vccd1 vccd1 _20949_/C sky130_fd_sc_hd__nor2_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ _20877_/A _20877_/B vssd1 vssd1 vccd1 vccd1 _20879_/A sky130_fd_sc_hd__xor2_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22616_ _22616_/A vssd1 vssd1 vccd1 vccd1 _22796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11967__B1 _11965_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22547_ _22766_/Q input40/X _22547_/S vssd1 vssd1 vccd1 vccd1 _22548_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18895__A1 _11636_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18895__B2 _15888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ _12300_/A _12300_/B _12387_/A vssd1 vssd1 vccd1 vccd1 _12437_/A sky130_fd_sc_hd__nand3_2
XFILLER_154_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ _13271_/A _13633_/B _13633_/C _13272_/Y _13275_/X vssd1 vssd1 vccd1 vccd1
+ _13281_/B sky130_fd_sc_hd__o32ai_1
XANTENNA__11968__B _11968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22478_ _21169_/A input41/X _22486_/S vssd1 vssd1 vccd1 vccd1 _22479_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ _12231_/A _12231_/B _12231_/C vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__nand3_1
XANTENNA__18647__A1 _11819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21429_ _21297_/Y _21420_/X _21423_/Y vssd1 vssd1 vccd1 vccd1 _21565_/B sky130_fd_sc_hd__o21ai_1
XFILLER_170_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18111__A3 _12098_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ _12162_/A _15774_/B _19490_/C _19490_/D vssd1 vssd1 vccd1 vccd1 _12162_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12931__A2 _12968_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18373__A2_N _18387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16970_ _16978_/A _16978_/B _16968_/X _16969_/X vssd1 vssd1 vccd1 vccd1 _16970_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_123_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12093_ _12135_/A vssd1 vssd1 vccd1 vccd1 _19358_/C sky130_fd_sc_hd__buf_2
XFILLER_104_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15921_ _15921_/A _16157_/D _17652_/B _16414_/A vssd1 vssd1 vccd1 vccd1 _15921_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__20206__B2 _20101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19072__A1 _11380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15175__B _15175_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18640_ _18634_/Y _18638_/X _18933_/C vssd1 vssd1 vccd1 vccd1 _18646_/A sky130_fd_sc_hd__o21bai_2
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18280__C1 _19358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15852_ _15828_/X _15826_/Y _15836_/X vssd1 vssd1 vccd1 vccd1 _15853_/A sky130_fd_sc_hd__a21oi_2
XFILLER_92_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18486__B _18691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _14805_/A _14895_/B _14805_/C _14805_/D vssd1 vssd1 vccd1 vccd1 _14806_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _18402_/A _18571_/B _18571_/C _18571_/D vssd1 vssd1 vccd1 vccd1 _18571_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _15783_/A _15783_/B _15783_/C vssd1 vssd1 vccd1 vccd1 _15915_/B sky130_fd_sc_hd__nand3_2
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20509__A2 _16779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ _12990_/A _13031_/A _12994_/X vssd1 vssd1 vccd1 vccd1 _13037_/B sky130_fd_sc_hd__a21o_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17821__D _17833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17522_ _17585_/A vssd1 vssd1 vccd1 vccd1 _17701_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _14737_/A _14737_/B _14738_/B vssd1 vssd1 vccd1 vccd1 _14734_/Y sky130_fd_sc_hd__a21boi_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _18292_/A _11731_/A _11935_/B _11936_/Y _11938_/Y vssd1 vssd1 vccd1 vccd1
+ _11947_/C sky130_fd_sc_hd__o221ai_4
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17453_ _17304_/B _17307_/B _17307_/C vssd1 vssd1 vccd1 vccd1 _17454_/C sky130_fd_sc_hd__a21boi_1
XFILLER_72_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14665_ _14665_/A _14843_/C vssd1 vssd1 vccd1 vccd1 _22674_/D sky130_fd_sc_hd__xor2_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _11378_/X _11299_/X _11420_/C _11349_/X _18259_/A vssd1 vssd1 vccd1 vccd1
+ _11877_/Y sky130_fd_sc_hd__a311oi_4
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16404_ _16433_/A _16433_/B _16433_/C vssd1 vssd1 vccd1 vccd1 _16406_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__18933__C _18933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13616_ _13616_/A _13616_/B _13616_/C vssd1 vssd1 vccd1 vccd1 _13617_/C sky130_fd_sc_hd__nand3_1
XFILLER_158_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17384_ _19496_/A vssd1 vssd1 vccd1 vccd1 _17525_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__18335__B1 _11774_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14596_ _13748_/X _14562_/X _14942_/C _14729_/A _14591_/X vssd1 vssd1 vccd1 vccd1
+ _14712_/B sky130_fd_sc_hd__o311a_1
XANTENNA__11958__B1 _18292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19123_ _18812_/Y _19113_/X _18830_/B vssd1 vssd1 vccd1 vccd1 _19123_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16335_ _16310_/Y _16315_/X _16354_/A vssd1 vssd1 vccd1 vccd1 _16342_/A sky130_fd_sc_hd__o21ai_2
XFILLER_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13547_ _13550_/A _13469_/A _13550_/B vssd1 vssd1 vccd1 vccd1 _13551_/A sky130_fd_sc_hd__a21o_1
XFILLER_158_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20693__A1 _13022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19054_ _18611_/Y _19051_/X _19052_/Y _19053_/X vssd1 vssd1 vccd1 vccd1 _19231_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16266_ _16266_/A vssd1 vssd1 vccd1 vccd1 _16266_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13478_ _13501_/A _13550_/C _13477_/X vssd1 vssd1 vccd1 vccd1 _13478_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18005_ _18055_/A _18055_/B _22905_/Q vssd1 vssd1 vccd1 vccd1 _18053_/C sky130_fd_sc_hd__nand3_1
XFILLER_161_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15217_ _15217_/A _15217_/B _15217_/C vssd1 vssd1 vccd1 vccd1 _15217_/X sky130_fd_sc_hd__and3_1
XFILLER_161_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12429_ _12314_/Y _12329_/X _12428_/Y _12334_/X vssd1 vssd1 vccd1 vccd1 _12429_/X
+ sky130_fd_sc_hd__o211a_1
X_16197_ _16183_/Y _16187_/Y _16195_/Y _16196_/Y vssd1 vssd1 vccd1 vccd1 _16202_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_160_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16649__B1 _16650_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15148_ _15148_/A vssd1 vssd1 vccd1 vccd1 _15152_/B sky130_fd_sc_hd__inv_2
XFILLER_141_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19956_ _19860_/Y _19863_/Y _19916_/A vssd1 vssd1 vccd1 vccd1 _19956_/X sky130_fd_sc_hd__o21a_1
XFILLER_141_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15079_ _13851_/A _13851_/B _15182_/A vssd1 vssd1 vccd1 vccd1 _15085_/A sky130_fd_sc_hd__a21o_1
XANTENNA__14270__A _14270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14675__A2 _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18907_ _18907_/A _18907_/B _18907_/C vssd1 vssd1 vccd1 vccd1 _18908_/C sky130_fd_sc_hd__nand3_2
X_19887_ _19890_/A _19887_/B _19887_/C vssd1 vssd1 vccd1 vccd1 _19889_/A sky130_fd_sc_hd__and3_1
XFILLER_122_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13883__B1 _14721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18838_ _18725_/A _18741_/D _18836_/Y _18837_/X vssd1 vssd1 vccd1 vccd1 _18914_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22902__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18769_ _18770_/A _18779_/B _18770_/C vssd1 vssd1 vccd1 vccd1 _18769_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20800_ _20799_/A _20799_/B _20869_/A _20799_/D vssd1 vssd1 vccd1 vccd1 _20803_/C
+ sky130_fd_sc_hd__a22o_1
X_21780_ _21779_/X _21647_/Y _21624_/Y _21618_/Y vssd1 vssd1 vccd1 vccd1 _21781_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20731_ _20731_/A _20778_/A vssd1 vssd1 vccd1 vccd1 _20737_/B sky130_fd_sc_hd__nand2_1
XANTENNA__15388__B1 _15389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16925__A _18666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14150__A1_N _14147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20662_ _20548_/X _20551_/Y _20554_/Y vssd1 vssd1 vccd1 vccd1 _20827_/A sky130_fd_sc_hd__a21oi_1
XFILLER_195_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18326__B1 _19496_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22401_ _22401_/A vssd1 vssd1 vccd1 vccd1 _22701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20593_ _20593_/A _20593_/B _20593_/C _20593_/D vssd1 vssd1 vccd1 vccd1 _20682_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_177_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14445__A _16400_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22332_ _22310_/A _22313_/A _22329_/Y _22330_/Y vssd1 vssd1 vccd1 vccd1 _22333_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_52_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22662__A _22662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16352__A2 _21011_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14363__A1 _18128_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22263_ _22304_/B _22263_/B _22263_/C vssd1 vssd1 vccd1 vccd1 _22302_/A sky130_fd_sc_hd__and3_1
XFILLER_191_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14363__B2 _14362_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19674__C _22919_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20436__A1 _20553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21214_ _21214_/A vssd1 vssd1 vccd1 vccd1 _21724_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22194_ _22194_/A _22194_/B vssd1 vssd1 vccd1 vccd1 _22195_/B sky130_fd_sc_hd__xnor2_1
XFILLER_183_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12059__A_N _11899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21145_ _21138_/X _21115_/Y _21079_/Y _21066_/X vssd1 vssd1 vccd1 vccd1 _21157_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21076_ _21076_/A _21076_/B _21076_/C _21076_/D vssd1 vssd1 vccd1 vccd1 _21076_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13874__B1 _14122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20027_ _20025_/X _20026_/Y _20005_/A vssd1 vssd1 vccd1 vccd1 _20029_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__21725__B _21725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18801__B2 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15615__A1 _18706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15615__B2 _18875_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16819__B _20928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _12008_/A vssd1 vssd1 vccd1 vccd1 _11800_/X sky130_fd_sc_hd__buf_4
XFILLER_55_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17368__A1 _22896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11970__C _18875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _22827_/Q vssd1 vssd1 vccd1 vccd1 _20452_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21978_ _22036_/B _22036_/C _21977_/A vssd1 vssd1 vccd1 vccd1 _21978_/X sky130_fd_sc_hd__a21o_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15379__B1 _15918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ _11731_/A vssd1 vssd1 vccd1 vccd1 _17427_/A sky130_fd_sc_hd__clkbuf_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ _20864_/B _20865_/Y _20866_/B vssd1 vssd1 vccd1 vccd1 _20930_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__16835__A _17436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20911__A2 _17440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14450_ _14443_/X _11334_/X _14448_/X vssd1 vssd1 vccd1 vccd1 _22665_/D sky130_fd_sc_hd__a21o_1
XANTENNA__19211__A _19211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _18648_/B vssd1 vssd1 vccd1 vccd1 _19322_/A sky130_fd_sc_hd__clkbuf_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16591__A2 _16879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16554__B _17530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13401_ _13401_/A vssd1 vssd1 vccd1 vccd1 _13664_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_168_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18868__A1 _12114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ _11593_/A vssd1 vssd1 vccd1 vccd1 _15904_/A sky130_fd_sc_hd__buf_2
X_14381_ _14411_/A vssd1 vssd1 vccd1 vccd1 _14381_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16120_ _16115_/X _16082_/B _16082_/A _16126_/A vssd1 vssd1 vccd1 vccd1 _16120_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13332_ _21362_/A _21990_/A _13332_/C _21739_/B vssd1 vssd1 vccd1 vccd1 _13337_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_183_844 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16051_ _20745_/C _16130_/A _16051_/C _16103_/D vssd1 vssd1 vccd1 vccd1 _16051_/X
+ sky130_fd_sc_hd__and4_1
X_13263_ _13237_/X _13272_/A _13438_/B vssd1 vssd1 vccd1 vccd1 _13481_/A sky130_fd_sc_hd__o21ai_2
XFILLER_182_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15002_ _15002_/A _15002_/B vssd1 vssd1 vccd1 vccd1 _15015_/A sky130_fd_sc_hd__nand2_1
XFILLER_182_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12214_ _16473_/A vssd1 vssd1 vccd1 vccd1 _18445_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_135_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13194_ _13376_/A vssd1 vssd1 vccd1 vccd1 _13521_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_194_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20092__A _20092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19810_ _19808_/A _19808_/B _19809_/A vssd1 vssd1 vccd1 vccd1 _19833_/A sky130_fd_sc_hd__a21o_1
XANTENNA__15303__B1 _12500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ _18677_/C vssd1 vssd1 vccd1 vccd1 _18116_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_2_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1097 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19741_ _19746_/A _19746_/C vssd1 vssd1 vccd1 vccd1 _19741_/X sky130_fd_sc_hd__and2_1
XFILLER_173_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16953_ _12727_/A _17137_/A _16494_/A _16956_/A vssd1 vssd1 vccd1 vccd1 _16954_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_150_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12076_ _11914_/Y _11606_/X _11923_/A _11918_/Y _11923_/B vssd1 vssd1 vccd1 vccd1
+ _12076_/X sky130_fd_sc_hd__o2111a_1
XFILLER_104_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22925__CLK _22948_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15904_ _15904_/A vssd1 vssd1 vccd1 vccd1 _15904_/X sky130_fd_sc_hd__buf_4
X_19672_ _19293_/X _19294_/X _19569_/A _19669_/Y _19761_/D vssd1 vssd1 vccd1 vccd1
+ _19674_/B sky130_fd_sc_hd__o221ai_4
XFILLER_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16884_ _16879_/B _17840_/A _16879_/A _16880_/X vssd1 vssd1 vccd1 vccd1 _16884_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_37_416 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18623_ _18623_/A _18623_/B _18623_/C vssd1 vssd1 vccd1 vccd1 _18624_/A sky130_fd_sc_hd__nand3_1
XFILLER_2_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13880__A3 _14808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _15921_/A _16613_/C _17652_/B _16414_/A vssd1 vssd1 vccd1 vccd1 _16414_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA__15633__B _15633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18554_ _18554_/A _18554_/B vssd1 vssd1 vccd1 vccd1 _18555_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _15766_/A _15859_/C _15859_/D vssd1 vssd1 vccd1 vccd1 _15766_/X sky130_fd_sc_hd__and3_1
XFILLER_46_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ _12522_/A _12522_/B _12968_/A _20697_/A _12930_/A vssd1 vssd1 vccd1 vccd1
+ _12981_/C sky130_fd_sc_hd__a2111o_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17505_ _17800_/D vssd1 vssd1 vccd1 vccd1 _17910_/D sky130_fd_sc_hd__clkbuf_2
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14717_ _14714_/C _14717_/B _14717_/C vssd1 vssd1 vccd1 vccd1 _14737_/B sky130_fd_sc_hd__nand3b_2
X_18485_ _18340_/B _18482_/Y _18488_/A vssd1 vssd1 vccd1 vccd1 _18487_/A sky130_fd_sc_hd__o21ai_1
X_11929_ _11837_/B _11831_/C _12084_/A vssd1 vssd1 vccd1 vccd1 _12245_/A sky130_fd_sc_hd__a21boi_1
X_15697_ _18666_/B _15774_/D _15457_/A _15696_/Y vssd1 vssd1 vccd1 vccd1 _15698_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16745__A _16745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17436_ _17436_/A _21011_/C _17462_/A vssd1 vssd1 vccd1 vccd1 _17436_/X sky130_fd_sc_hd__and3_1
X_14648_ _14750_/B _14651_/B vssd1 vssd1 vccd1 vccd1 _14649_/C sky130_fd_sc_hd__and2_1
XFILLER_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11889__A _16103_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17367_ _17220_/A _17219_/A _17219_/B _17071_/A vssd1 vssd1 vccd1 vccd1 _17367_/Y
+ sky130_fd_sc_hd__o31ai_2
X_14579_ _14468_/B _14685_/A _14576_/X _14942_/B _14568_/Y vssd1 vssd1 vccd1 vccd1
+ _14602_/C sky130_fd_sc_hd__o221ai_2
X_19106_ _19106_/A _19106_/B _19106_/C _19106_/D vssd1 vssd1 vccd1 vccd1 _19257_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_118_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16318_ _16318_/A vssd1 vssd1 vccd1 vccd1 _16435_/B sky130_fd_sc_hd__buf_4
X_17298_ _17298_/A _17298_/B _17298_/C vssd1 vssd1 vccd1 vccd1 _17299_/B sky130_fd_sc_hd__nand3_1
XFILLER_158_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19037_ _19037_/A _19037_/B _19037_/C vssd1 vssd1 vccd1 vccd1 _19037_/X sky130_fd_sc_hd__and3_1
XANTENNA__14345__A1 _18115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15542__B1 _12968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16249_ _16248_/X _16179_/A _15589_/X _16474_/A _16221_/Y vssd1 vssd1 vccd1 vccd1
+ _16250_/C sky130_fd_sc_hd__o221ai_2
XANTENNA__14345__B2 _13736_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput102 _14422_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput113 _14350_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[9] sky130_fd_sc_hd__buf_2
Xoutput124 _22949_/Q vssd1 vssd1 vccd1 vccd1 y[8] sky130_fd_sc_hd__buf_2
XFILLER_127_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_bq_clk_i clkbuf_3_6_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _22922_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_82_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19939_ _19939_/A vssd1 vssd1 vccd1 vccd1 _19939_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20730__A _20818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22950_ _22951_/CLK _22950_/D vssd1 vssd1 vccd1 vccd1 _22950_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18200__A _18200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22591__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21901_ _21901_/A _21996_/A _21933_/B vssd1 vssd1 vccd1 vccd1 _21901_/Y sky130_fd_sc_hd__nand3_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11882__A2 _19202_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22881_ _22916_/CLK input75/X vssd1 vssd1 vccd1 vccd1 _22881_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19339__A2 _19512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21832_ _21832_/A _21832_/B _21832_/C vssd1 vssd1 vccd1 vccd1 _21832_/X sky130_fd_sc_hd__and3_1
XANTENNA__11790__C _11790_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18547__B1 _18546_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21763_ _21763_/A _21763_/B vssd1 vssd1 vccd1 vccd1 _21846_/D sky130_fd_sc_hd__nand2_1
XANTENNA__20354__B1 _20358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20714_ _20711_/Y _20712_/Y _20720_/A vssd1 vssd1 vccd1 vccd1 _20714_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_168_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21694_ _21837_/A _21837_/B vssd1 vssd1 vccd1 vccd1 _21695_/C sky130_fd_sc_hd__and2_1
XFILLER_52_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_839 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20645_ _20645_/A _20645_/B _20645_/C vssd1 vssd1 vccd1 vccd1 _20650_/B sky130_fd_sc_hd__nand3_2
XFILLER_149_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21854__B1 _21853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20576_ _20582_/A _20576_/B _20582_/C vssd1 vssd1 vccd1 vccd1 _20577_/B sky130_fd_sc_hd__nand3_2
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11949__D _11949_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14336__A1 _12387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22315_ _22314_/A _22314_/B _22314_/C vssd1 vssd1 vccd1 vccd1 _22316_/B sky130_fd_sc_hd__o21a_1
XFILLER_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22246_ _22216_/B _22202_/A _22244_/Y vssd1 vssd1 vccd1 vccd1 _22246_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22948__CLK _22948_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17286__B1 _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22177_ _22176_/A _22265_/B _22176_/C _22238_/A vssd1 vssd1 vccd1 vccd1 _22178_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_87_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21128_ _21128_/A _21128_/B vssd1 vssd1 vccd1 vccd1 _21129_/A sky130_fd_sc_hd__or2_1
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13950_ _14502_/A vssd1 vssd1 vccd1 vccd1 _13950_/X sky130_fd_sc_hd__clkbuf_2
X_21059_ _21006_/B _21062_/B _21057_/Y _21058_/Y vssd1 vssd1 vccd1 vccd1 _21068_/A
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__18110__A _18810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22582__A1 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12901_ _13007_/B _13007_/C _12750_/B vssd1 vssd1 vccd1 vccd1 _12966_/A sky130_fd_sc_hd__a21bo_1
XFILLER_143_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13881_ _13881_/A _13881_/B vssd1 vssd1 vccd1 vccd1 _13881_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15620_ _15646_/A _16332_/A vssd1 vssd1 vccd1 vccd1 _16397_/A sky130_fd_sc_hd__nor2_2
XFILLER_59_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12832_ _15617_/A _12827_/X _20357_/B _20092_/A vssd1 vssd1 vccd1 vccd1 _12832_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_15_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_622 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15551_ _16477_/A vssd1 vssd1 vccd1 vccd1 _19358_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12763_ _12891_/A _12763_/B vssd1 vssd1 vccd1 vccd1 _12763_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11625__A2 _11395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18483__C _18691_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14502_/A vssd1 vssd1 vccd1 vccd1 _14818_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18270_ _18251_/A _18257_/B _12256_/A _18251_/Y vssd1 vssd1 vccd1 vccd1 _18430_/A
+ sky130_fd_sc_hd__o211ai_4
X_11714_ _11714_/A vssd1 vssd1 vccd1 vccd1 _15536_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _15482_/A _15482_/B _15482_/C _15482_/D vssd1 vssd1 vccd1 vccd1 _15522_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _17246_/A vssd1 vssd1 vccd1 vccd1 _16937_/B sky130_fd_sc_hd__clkbuf_4
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17221_ _22895_/Q vssd1 vssd1 vccd1 vccd1 _17221_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _22965_/Q _22966_/Q vssd1 vssd1 vccd1 vccd1 _16481_/C sky130_fd_sc_hd__nor2_2
XANTENNA__22098__B1 _21269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11645_ _11645_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _11645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11502__A _11502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17152_ _16060_/A _16758_/X _17149_/A vssd1 vssd1 vccd1 vccd1 _17155_/A sky130_fd_sc_hd__o21ai_1
X_14364_ _16322_/B _14344_/X _14351_/X _14359_/X _14363_/X vssd1 vssd1 vccd1 vccd1
+ _14364_/X sky130_fd_sc_hd__a221o_1
Xinput15 wb_adr_i[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput26 wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_2
X_11576_ _11839_/A _11576_/B vssd1 vssd1 vccd1 vccd1 _11577_/B sky130_fd_sc_hd__nand2_1
XFILLER_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 wb_dat_i[11] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_4
X_16103_ _20390_/C _16150_/A _16103_/C _16103_/D vssd1 vssd1 vccd1 vccd1 _16150_/B
+ sky130_fd_sc_hd__nand4_2
Xinput48 wb_dat_i[21] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput59 wb_dat_i[31] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_2
XANTENNA__14327__A1 _11306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13315_ _13354_/A vssd1 vssd1 vccd1 vccd1 _13315_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15524__B1 _12929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17083_ _17083_/A vssd1 vssd1 vccd1 vccd1 _17083_/X sky130_fd_sc_hd__buf_4
XFILLER_122_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14327__B2 _13761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14295_ input23/X vssd1 vssd1 vccd1 vccd1 _22586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16034_ _16034_/A _16210_/A _16034_/C vssd1 vssd1 vccd1 vccd1 _16035_/B sky130_fd_sc_hd__nand3_1
XFILLER_182_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13246_ _13273_/B _13421_/A _13273_/A vssd1 vssd1 vccd1 vccd1 _13272_/A sky130_fd_sc_hd__nand3_2
XFILLER_124_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17277__B1 _11672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13177_ _13344_/A _13345_/A _13633_/A vssd1 vssd1 vccd1 vccd1 _13216_/A sky130_fd_sc_hd__a21o_1
XANTENNA__15347__C _16313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12128_ _18141_/A vssd1 vssd1 vccd1 vccd1 _12128_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17985_ _19419_/B vssd1 vssd1 vccd1 vccd1 _18030_/A sky130_fd_sc_hd__buf_2
XFILLER_123_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19724_ _19724_/A _19724_/B vssd1 vssd1 vccd1 vccd1 _19725_/A sky130_fd_sc_hd__nand2_1
X_16936_ _17631_/A vssd1 vssd1 vccd1 vccd1 _19496_/A sky130_fd_sc_hd__buf_2
X_12059_ _11899_/A _12059_/B _12247_/B vssd1 vssd1 vccd1 vccd1 _12061_/B sky130_fd_sc_hd__nand3b_1
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16237__D1 _15991_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19655_ _19653_/Y _19658_/A _19545_/Y _19555_/C vssd1 vssd1 vccd1 vccd1 _19814_/A
+ sky130_fd_sc_hd__o211a_1
X_16867_ _16867_/A _16867_/B _16867_/C vssd1 vssd1 vccd1 vccd1 _16873_/D sky130_fd_sc_hd__nand3_1
XFILLER_37_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15363__B _16322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16252__A1 _15545_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17281__D _18839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18606_ _18606_/A _18606_/B vssd1 vssd1 vccd1 vccd1 _22892_/D sky130_fd_sc_hd__xnor2_1
X_15818_ _15727_/A _15727_/B _15825_/B _15825_/C vssd1 vssd1 vccd1 vccd1 _15819_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_80_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19586_ _19602_/A _19602_/B _18156_/X _17819_/A vssd1 vssd1 vccd1 vccd1 _19607_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16798_ _15840_/A _15903_/X _20255_/A _16792_/A vssd1 vssd1 vccd1 vccd1 _16798_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18674__B _18698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18537_ _12157_/X _12158_/X _11561_/X _11563_/X vssd1 vssd1 vccd1 vccd1 _18537_/X
+ sky130_fd_sc_hd__a22o_2
X_15749_ _15479_/A _15448_/X _15517_/A _15517_/B vssd1 vssd1 vccd1 vccd1 _15756_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18544__A3 _12111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18468_ _18465_/X _18467_/Y _18462_/A vssd1 vssd1 vccd1 vccd1 _18474_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__15810__C _15810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17419_ _17413_/Y _17414_/X _17399_/Y _17410_/X vssd1 vssd1 vccd1 vccd1 _17420_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_21_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18399_ _18183_/Y _18395_/X _18396_/Y _18398_/Y vssd1 vssd1 vccd1 vccd1 _18399_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__18690__A _18690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20639__A1 _20449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20430_ _20281_/B _20429_/X _20420_/A _20413_/A vssd1 vssd1 vccd1 vccd1 _20431_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20361_ _20354_/X _20511_/B _20360_/X vssd1 vssd1 vccd1 vccd1 _20366_/A sky130_fd_sc_hd__o21ai_1
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22100_ _22098_/X _22100_/B _22100_/C vssd1 vssd1 vccd1 vccd1 _22102_/B sky130_fd_sc_hd__nand3b_1
XFILLER_161_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20292_ _20293_/A _20293_/B _20298_/A _20298_/B vssd1 vssd1 vccd1 vccd1 _20292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22031_ _22031_/A _22031_/B _22031_/C _22172_/A vssd1 vssd1 vccd1 vccd1 _22196_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15818__A1 _15727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21556__A _21556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_872 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16369__B _16627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22933_ _22933_/CLK _22933_/D vssd1 vssd1 vccd1 vccd1 _22933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22864_ _22943_/CLK _22876_/Q vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21815_ _21837_/A _21815_/B _21837_/C _21837_/D vssd1 vssd1 vccd1 vccd1 _21834_/C
+ sky130_fd_sc_hd__nand4_2
X_22795_ _22795_/CLK _22795_/D vssd1 vssd1 vccd1 vccd1 _22795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13802__A _22867_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21746_ _21610_/B _21740_/X _22057_/B _21742_/Y _22176_/A vssd1 vssd1 vccd1 vccd1
+ _21761_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_25_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13521__B _13521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14557__A1 _14843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21677_ _21677_/A _21677_/B vssd1 vssd1 vccd1 vccd1 _21677_/X sky130_fd_sc_hd__or2_1
XFILLER_40_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11322__A _22954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ _11608_/A _11430_/B _11430_/C vssd1 vssd1 vccd1 vccd1 _11431_/B sky130_fd_sc_hd__nand3_2
XANTENNA__18299__A2 _15541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12032__A2 _11762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20628_ _20629_/A _20629_/B _20629_/C _20702_/B vssd1 vssd1 vccd1 vccd1 _20634_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _11361_/A vssd1 vssd1 vccd1 vccd1 _15932_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_138_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20559_ _20559_/A _20559_/B vssd1 vssd1 vccd1 vccd1 _20564_/A sky130_fd_sc_hd__and2_1
XFILLER_164_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18105__A _19061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16551__C _20092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13100_ _13099_/B _14380_/A _13095_/X vssd1 vssd1 vccd1 vccd1 _13101_/B sky130_fd_sc_hd__a21bo_1
X_11292_ _22954_/Q _22953_/Q _22968_/Q vssd1 vssd1 vccd1 vccd1 _11325_/B sky130_fd_sc_hd__o21ai_4
X_14080_ _13948_/X _13949_/X _14618_/A vssd1 vssd1 vccd1 vccd1 _14149_/B sky130_fd_sc_hd__a21o_1
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13031_ _13031_/A _13031_/B vssd1 vssd1 vccd1 vccd1 _13031_/Y sky130_fd_sc_hd__nand2_1
XFILLER_152_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22229_ _22229_/A _22229_/B _22229_/C vssd1 vssd1 vccd1 vccd1 _22233_/A sky130_fd_sc_hd__and3_1
XFILLER_79_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11543__A1 _11541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15809__A1 _12772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15809__B2 _15808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input45_A wb_dat_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15464__A _16256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17770_ _17695_/A _17727_/X _17697_/C _17769_/Y vssd1 vssd1 vccd1 vccd1 _17785_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14982_ _14982_/A _14982_/B _14982_/C vssd1 vssd1 vccd1 vccd1 _14982_/Y sky130_fd_sc_hd__nand3_1
XFILLER_66_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16721_ _16312_/X _16714_/X _16720_/Y vssd1 vssd1 vccd1 vccd1 _16721_/X sky130_fd_sc_hd__a21o_1
X_13933_ _13948_/A _13949_/A _14624_/A vssd1 vssd1 vccd1 vccd1 _13933_/X sky130_fd_sc_hd__a21o_1
XANTENNA__18197__D _18288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16234__A1 _12719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19440_ _19446_/A _19561_/B vssd1 vssd1 vccd1 vccd1 _19440_/X sky130_fd_sc_hd__and2_1
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16652_ _16652_/A _16652_/B vssd1 vssd1 vccd1 vccd1 _16653_/C sky130_fd_sc_hd__nand2_1
XFILLER_47_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13864_ _14118_/B vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15603_ _22698_/Q _22699_/Q vssd1 vssd1 vccd1 vccd1 _16319_/B sky130_fd_sc_hd__nor2_2
X_19371_ _19371_/A _19379_/A vssd1 vssd1 vccd1 vccd1 _19376_/A sky130_fd_sc_hd__nand2_1
X_12815_ _12333_/B _20219_/A _12596_/A _15637_/A _12808_/Y vssd1 vssd1 vccd1 vccd1
+ _12818_/B sky130_fd_sc_hd__o221ai_1
X_16583_ _14369_/X _16324_/B _16571_/Y _16324_/C vssd1 vssd1 vccd1 vccd1 _16584_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_76_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15993__B1 _20452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13795_ _22868_/Q vssd1 vssd1 vccd1 vccd1 _13989_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18322_ _19322_/B _19322_/C _16078_/C _19194_/A _19329_/C vssd1 vssd1 vccd1 vccd1
+ _18322_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_43_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14260__A3 _14181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15534_ _22961_/Q _22962_/Q _22662_/B _22964_/Q vssd1 vssd1 vccd1 vccd1 _16481_/D
+ sky130_fd_sc_hd__nor4_2
XFILLER_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _12624_/A _12619_/A _12745_/C vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15630__C _15912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11614__A_N _11606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18253_ _18232_/X _18233_/Y _18224_/Y _18230_/Y vssd1 vssd1 vccd1 vccd1 _18772_/C
+ sky130_fd_sc_hd__o211ai_4
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15465_ _14438_/A _11560_/C _11667_/Y _11668_/Y vssd1 vssd1 vccd1 vccd1 _15465_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12677_ _16932_/C vssd1 vssd1 vccd1 vccd1 _12689_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_124_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17204_ _17205_/C _17205_/B _17205_/A vssd1 vssd1 vccd1 vccd1 _17206_/A sky130_fd_sc_hd__a21o_1
XFILLER_175_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14416_ _22810_/Q _14411_/X _14412_/X _14413_/X _22778_/Q vssd1 vssd1 vccd1 vccd1
+ _14416_/X sky130_fd_sc_hd__a32o_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18184_ _18184_/A _18184_/B vssd1 vssd1 vccd1 vccd1 _18395_/B sky130_fd_sc_hd__nand2_1
X_11628_ _18716_/A vssd1 vssd1 vccd1 vccd1 _17312_/A sky130_fd_sc_hd__buf_4
X_15396_ _19329_/D _18130_/C _15909_/A _17128_/B vssd1 vssd1 vccd1 vccd1 _15396_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12023__A2 _11809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17135_ _12207_/X _15919_/A _16932_/Y _17133_/Y _17288_/A vssd1 vssd1 vccd1 vccd1
+ _17270_/B sky130_fd_sc_hd__o221ai_4
XFILLER_128_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20097__A2 _12576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14347_ _11771_/X _14338_/X _14339_/X _14334_/X _13896_/A vssd1 vssd1 vccd1 vccd1
+ _14347_/X sky130_fd_sc_hd__a32o_1
X_11559_ _11659_/D vssd1 vssd1 vccd1 vccd1 _11560_/C sky130_fd_sc_hd__buf_2
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11782__A1 _18116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17066_ _16665_/X _17371_/A _17215_/D _17373_/A vssd1 vssd1 vccd1 vccd1 _17222_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ _14276_/D _14834_/C _14834_/A _14269_/A _14263_/C vssd1 vssd1 vccd1 vccd1
+ _14279_/D sky130_fd_sc_hd__a32o_1
XFILLER_170_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16017_ _16015_/X _13022_/D _16016_/X _13022_/A vssd1 vssd1 vccd1 vccd1 _16017_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_98_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13229_ _13229_/A vssd1 vssd1 vccd1 vccd1 _13423_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12063__A _12116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19772__C _19772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21597__A2 _21594_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18998__B1 _15427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21376__A _21964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22910__D _22910_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13309__D _13521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15374__A _15389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _17968_/A _17968_/B vssd1 vssd1 vccd1 vccd1 _18007_/D sky130_fd_sc_hd__nor2_1
XFILLER_112_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14484__B1 _13904_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19707_ _19704_/Y _19706_/X _19709_/C vssd1 vssd1 vccd1 vccd1 _19707_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16919_ _16919_/A _16919_/B _16919_/C vssd1 vssd1 vccd1 vccd1 _16930_/A sky130_fd_sc_hd__nand3_1
X_17899_ _17899_/A _17899_/B vssd1 vssd1 vccd1 vccd1 _18020_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11407__A _11727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19638_ _19488_/A _19636_/X _19637_/Y vssd1 vssd1 vccd1 vccd1 _19638_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19569_ _19569_/A _19669_/A _19669_/B _19750_/A vssd1 vssd1 vccd1 vccd1 _19571_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19714__A2 _19517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21600_ _21478_/X _21596_/A _21481_/B _21482_/Y vssd1 vssd1 vccd1 vccd1 _21604_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22580_ _22781_/Q input56/X _22580_/S vssd1 vssd1 vccd1 vccd1 _22581_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19012__C _19012_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21531_ _21531_/A _21531_/B _21531_/C vssd1 vssd1 vccd1 vccd1 _21531_/X sky130_fd_sc_hd__and3_1
XFILLER_166_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_736 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1080 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21462_ _21173_/Y _21449_/A _21372_/C _21372_/B vssd1 vssd1 vccd1 vccd1 _21463_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20413_ _20413_/A vssd1 vssd1 vccd1 vccd1 _20545_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15549__A _16964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21393_ _21393_/A _21393_/B _21393_/C vssd1 vssd1 vccd1 vccd1 _21403_/A sky130_fd_sc_hd__nand3_2
XFILLER_174_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20344_ _20083_/X _20339_/A _20457_/B _20457_/A vssd1 vssd1 vccd1 vccd1 _20344_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_88_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20275_ _20143_/A _20143_/B _20125_/A vssd1 vssd1 vccd1 vccd1 _20275_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_150_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22014_ _22014_/A _22014_/B vssd1 vssd1 vccd1 vccd1 _22086_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12722__B1 _12968_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13817__A3 _13815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13516__B _21591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17413__B1 _17412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__A _11790_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22916_ _22916_/CLK _22916_/D vssd1 vssd1 vccd1 vccd1 _22916_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_856 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22847_ _22915_/CLK hold21/X vssd1 vssd1 vccd1 vccd1 _22847_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14628__A _15008_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12424_/Y _15450_/A _20471_/C _16261_/B _12595_/Y vssd1 vssd1 vccd1 vccd1
+ _12601_/C sky130_fd_sc_hd__o2111ai_4
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13591_/A vssd1 vssd1 vccd1 vccd1 _21489_/A sky130_fd_sc_hd__buf_2
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22778_ _22810_/CLK _22778_/D vssd1 vssd1 vccd1 vccd1 _22778_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _22825_/Q vssd1 vssd1 vccd1 vccd1 _12789_/A sky130_fd_sc_hd__inv_2
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21729_ _21853_/A _21341_/A _21728_/Y vssd1 vssd1 vccd1 vccd1 _21730_/D sky130_fd_sc_hd__o21ai_4
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _15230_/A _15247_/X _15249_/Y vssd1 vssd1 vccd1 vccd1 _15252_/A sky130_fd_sc_hd__o21a_1
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12005__A2 _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12462_ _12734_/A _12420_/X _12424_/Y _15569_/A _12449_/Y vssd1 vssd1 vccd1 vccd1
+ _12462_/Y sky130_fd_sc_hd__o221ai_1
XANTENNA__19469__B2 _19308_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14201_ _14231_/A _14231_/B _14693_/D _14786_/B _14199_/A vssd1 vssd1 vccd1 vccd1
+ _14201_/X sky130_fd_sc_hd__a32o_1
XANTENNA__11987__A _15482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ _15482_/A _11988_/A _11464_/A vssd1 vssd1 vccd1 vccd1 _11756_/A sky130_fd_sc_hd__o21ai_1
X_15181_ _15181_/A _15181_/B vssd1 vssd1 vccd1 vccd1 _15200_/A sky130_fd_sc_hd__or2_1
X_12393_ _22822_/Q vssd1 vssd1 vccd1 vccd1 _20359_/B sky130_fd_sc_hd__inv_2
XFILLER_193_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _14131_/X _14191_/A _14126_/Y _14085_/Y vssd1 vssd1 vccd1 vccd1 _14237_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16152__B1 _12772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ _11420_/A _12148_/B _11471_/C vssd1 vssd1 vccd1 vccd1 _12090_/A sky130_fd_sc_hd__a21oi_2
XFILLER_192_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14702__A1 _14366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18940_ _18757_/X _18758_/Y _18765_/X _18754_/X vssd1 vssd1 vccd1 vccd1 _18941_/C
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_98_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14063_ _13861_/Y _13862_/X _14169_/A _14169_/B vssd1 vssd1 vccd1 vccd1 _14167_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _11995_/B vssd1 vssd1 vccd1 vccd1 _11783_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13014_ _13011_/C _13009_/Y _13000_/X _13039_/A vssd1 vssd1 vccd1 vccd1 _13040_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_18871_ _19091_/C _19091_/A _18863_/Y _18870_/Y vssd1 vssd1 vccd1 vccd1 _18871_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16455__A1 _15530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15258__A2 _15259_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22666__CLK _22959_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17822_ _17822_/A vssd1 vssd1 vccd1 vccd1 _19839_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16341__A_N _16354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22528__A1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12611__A _16515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17753_ _17753_/A _17753_/B vssd1 vssd1 vccd1 vccd1 _17753_/Y sky130_fd_sc_hd__nor2_1
X_14965_ _14965_/A _14965_/B vssd1 vssd1 vccd1 vccd1 _14966_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12968__D _12968_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17404__B1 _18814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16704_ _16704_/A _16704_/B vssd1 vssd1 vccd1 vccd1 _16704_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13916_ _14021_/A _14021_/B vssd1 vssd1 vccd1 vccd1 _13916_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17684_ _17628_/Y _17629_/Y _17682_/Y _17683_/X vssd1 vssd1 vccd1 vccd1 _17697_/B
+ sky130_fd_sc_hd__o22ai_2
X_14896_ _14810_/X _14808_/Y _14809_/Y vssd1 vssd1 vccd1 vccd1 _14965_/B sky130_fd_sc_hd__a21boi_1
XFILLER_74_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19423_ _12064_/X _18023_/A _19306_/X _19211_/A vssd1 vssd1 vccd1 vccd1 _19424_/B
+ sky130_fd_sc_hd__o31a_1
X_16635_ _16635_/A vssd1 vssd1 vccd1 vccd1 _16895_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _14013_/A _14013_/B _13975_/D _14126_/A _14110_/B vssd1 vssd1 vccd1 vccd1
+ _13848_/A sky130_fd_sc_hd__a32o_1
XFILLER_90_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16939__B1_N _16976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13442__A _13475_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19354_ _17381_/X _17380_/X _19496_/B _19496_/C _18197_/C vssd1 vssd1 vccd1 vccd1
+ _19357_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16566_ _16566_/A vssd1 vssd1 vccd1 vccd1 _17874_/A sky130_fd_sc_hd__buf_2
XFILLER_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13778_ _13948_/A _13949_/A _14502_/A _14503_/A _14042_/A vssd1 vssd1 vccd1 vccd1
+ _14043_/A sky130_fd_sc_hd__a2111o_2
XFILLER_31_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18305_ _18305_/A _18305_/B _18305_/C _18305_/D vssd1 vssd1 vccd1 vccd1 _18572_/B
+ sky130_fd_sc_hd__nand4_4
X_15517_ _15517_/A _15517_/B vssd1 vssd1 vccd1 vccd1 _15517_/Y sky130_fd_sc_hd__nand2_1
X_19285_ _19443_/A _19681_/C _19681_/A vssd1 vssd1 vccd1 vccd1 _19286_/B sky130_fd_sc_hd__o21ai_1
XFILLER_149_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12729_ _12988_/B _15890_/A _20096_/A _12583_/A _12583_/C vssd1 vssd1 vccd1 vccd1
+ _12916_/B sky130_fd_sc_hd__o311a_1
X_16497_ _15536_/X _16240_/X _16484_/X _16483_/A _16483_/B vssd1 vssd1 vccd1 vccd1
+ _17646_/A sky130_fd_sc_hd__a32oi_4
XFILLER_148_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18236_ _18239_/B _18236_/B _18272_/B vssd1 vssd1 vccd1 vccd1 _18236_/Y sky130_fd_sc_hd__nand3_1
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15448_ _18197_/C _19351_/C _12913_/A _16106_/D _19694_/A vssd1 vssd1 vccd1 vccd1
+ _15448_/X sky130_fd_sc_hd__a32o_2
XFILLER_90_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_706 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22464__A0 _13304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18167_ _18167_/A vssd1 vssd1 vccd1 vccd1 _19199_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14941__A1 _15056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15379_ _15389_/B _15389_/C _15918_/A _17111_/A vssd1 vssd1 vccd1 vccd1 _15665_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__14941__B2 _14953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17118_ _20781_/B vssd1 vssd1 vccd1 vccd1 _21019_/B sky130_fd_sc_hd__buf_2
X_18098_ _18098_/A _18098_/B _18098_/C vssd1 vssd1 vccd1 vccd1 _18279_/A sky130_fd_sc_hd__nand3_4
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16694__A1 _22889_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17049_ _17049_/A _17049_/B vssd1 vssd1 vccd1 vccd1 _17049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11507__A1 _11502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11507__B2 _11505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20060_ _22927_/Q vssd1 vssd1 vccd1 vccd1 _20060_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12180__A1 _12164_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22519__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18199__A1 _11502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ _20901_/A _20960_/X _20961_/Y vssd1 vssd1 vccd1 vccd1 _20963_/B sky130_fd_sc_hd__o21ai_1
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22701_ _22701_/CLK _22701_/D vssd1 vssd1 vccd1 vccd1 _22701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14448__A _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20893_ _20891_/A _20891_/B _20842_/X vssd1 vssd1 vccd1 vccd1 _20894_/A sky130_fd_sc_hd__a21o_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22632_ _22643_/A vssd1 vssd1 vccd1 vccd1 _22641_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13432__B2 _21848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18862__B _18862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22563_ _22773_/Q input48/X _22569_/S vssd1 vssd1 vccd1 vccd1 _22564_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21514_ _21666_/B _21666_/A _21514_/C vssd1 vssd1 vccd1 vccd1 _21514_/X sky130_fd_sc_hd__and3b_1
XFILLER_166_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22494_ _22494_/A vssd1 vssd1 vccd1 vccd1 _22742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21445_ _21445_/A _22231_/D _21445_/C vssd1 vssd1 vccd1 vccd1 _21547_/A sky130_fd_sc_hd__and3_1
XFILLER_135_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11746__A1 _11606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21376_ _21964_/A vssd1 vssd1 vccd1 vccd1 _21376_/X sky130_fd_sc_hd__buf_2
XFILLER_162_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20913__A _20913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20327_ _20247_/Y _20326_/Y _20249_/B _20324_/Y _15909_/A vssd1 vssd1 vccd1 vccd1
+ _20328_/D sky130_fd_sc_hd__o2111ai_4
XANTENNA__22689__CLK _22690_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14911__A _14911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20258_ _12671_/X _12735_/X _20242_/X _20142_/B vssd1 vssd1 vccd1 vccd1 _20263_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20189_ _20189_/A _20189_/B _20189_/C vssd1 vssd1 vccd1 vccd1 _20189_/Y sky130_fd_sc_hd__nand3_1
XFILLER_77_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12788__D _20502_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15742__A _19587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ _14750_/A _14750_/B vssd1 vssd1 vccd1 vccd1 _14751_/B sky130_fd_sc_hd__nand2_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ _11751_/X _11703_/X _11935_/X vssd1 vssd1 vccd1 vccd1 _12219_/B sky130_fd_sc_hd__o21ai_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12474__A2 _12669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _22767_/Q vssd1 vssd1 vccd1 vccd1 _13733_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11682__B1 _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14681_ _14934_/A _14948_/C _14998_/A _14467_/X vssd1 vssd1 vccd1 vccd1 _14681_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _11895_/C _11893_/B vssd1 vssd1 vccd1 vccd1 _11894_/C sky130_fd_sc_hd__nand2_1
XFILLER_60_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16420_ _16695_/C _16695_/D vssd1 vssd1 vccd1 vccd1 _16424_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13632_ _13520_/B _13593_/X _21874_/A _13595_/Y _21399_/A vssd1 vssd1 vccd1 vccd1
+ _13666_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_189_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16351_ _16351_/A vssd1 vssd1 vccd1 vccd1 _16351_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__21497__A1 _21383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13563_ _13563_/A _13563_/B _13563_/C vssd1 vssd1 vccd1 vccd1 _13565_/B sky130_fd_sc_hd__nand3_1
XFILLER_158_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19587__C _19587_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16573__A _20579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ _15302_/A _15302_/B vssd1 vssd1 vccd1 vccd1 _15454_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19070_ _18912_/B _18912_/A _19091_/C _19091_/A vssd1 vssd1 vccd1 vccd1 _19148_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_12514_ _22823_/Q vssd1 vssd1 vccd1 vccd1 _12515_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16282_ _16282_/A _16288_/A vssd1 vssd1 vccd1 vccd1 _16606_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13494_ _13494_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _13498_/A sky130_fd_sc_hd__nand2_1
X_18021_ _17897_/A _17897_/B _17897_/C _18020_/C _17996_/A vssd1 vssd1 vccd1 vccd1
+ _18038_/A sky130_fd_sc_hd__a2111oi_1
XFILLER_12_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ _15233_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _22684_/D sky130_fd_sc_hd__xnor2_1
XFILLER_139_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12445_ _15394_/A _15799_/A _15799_/B _20694_/A vssd1 vssd1 vccd1 vccd1 _12445_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_166_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11510__A _18512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15164_ _15129_/A _15145_/Y _15162_/Y _15163_/X vssd1 vssd1 vccd1 vccd1 _15181_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12376_ _12343_/B _12341_/A _12363_/Y _15608_/C vssd1 vssd1 vccd1 vccd1 _12379_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_158_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14115_ _14165_/B _14115_/B _14115_/C vssd1 vssd1 vccd1 vccd1 _14285_/C sky130_fd_sc_hd__and3_1
XFILLER_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11327_ _11496_/B vssd1 vssd1 vccd1 vccd1 _11619_/B sky130_fd_sc_hd__buf_2
X_19972_ _19972_/A _19972_/B vssd1 vssd1 vccd1 vccd1 _22904_/D sky130_fd_sc_hd__xor2_1
X_15095_ _15095_/A _15095_/B _15095_/C vssd1 vssd1 vccd1 vccd1 _15097_/A sky130_fd_sc_hd__nand3_1
XFILLER_181_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18923_ _18917_/Y _18918_/Y _18919_/Y _18922_/Y vssd1 vssd1 vccd1 vccd1 _18977_/A
+ sky130_fd_sc_hd__o211ai_1
X_14046_ _14561_/C _14044_/Y _14045_/X vssd1 vssd1 vccd1 vccd1 _14098_/B sky130_fd_sc_hd__o21ai_4
XFILLER_122_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18854_ _18854_/A _18861_/A _18861_/B vssd1 vssd1 vccd1 vccd1 _19091_/C sky130_fd_sc_hd__nand3_1
XFILLER_122_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17805_ _19901_/A vssd1 vssd1 vccd1 vccd1 _17872_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18785_ _19293_/A _19294_/A _19138_/D _18607_/Y vssd1 vssd1 vccd1 vccd1 _18969_/B
+ sky130_fd_sc_hd__o211a_1
X_15997_ _18984_/A _18984_/B _15997_/C vssd1 vssd1 vccd1 vccd1 _15997_/X sky130_fd_sc_hd__and3_2
XANTENNA__21709__C1 _22675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18666__C _18839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15651__A2 _15319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17736_ _17736_/A _17736_/B vssd1 vssd1 vccd1 vccd1 _17736_/X sky130_fd_sc_hd__xor2_1
X_14948_ _15069_/A _15010_/C _14948_/C _15115_/C vssd1 vssd1 vccd1 vccd1 _15002_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_54_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11673__B1 _18288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15371__B _17424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17667_ _17660_/A _17660_/B _17662_/B vssd1 vssd1 vccd1 vccd1 _17667_/Y sky130_fd_sc_hd__a21boi_1
X_14879_ _14880_/B _14877_/C _14880_/A vssd1 vssd1 vccd1 vccd1 _14879_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16600__A1 _16354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19406_ _19404_/Y _19251_/Y _19405_/X _19261_/Y vssd1 vssd1 vccd1 vccd1 _19410_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16618_ _16624_/C _16873_/B vssd1 vssd1 vccd1 vccd1 _16619_/C sky130_fd_sc_hd__nand2_1
XFILLER_196_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17598_ _17704_/A vssd1 vssd1 vccd1 vccd1 _17600_/C sky130_fd_sc_hd__inv_2
XANTENNA__12217__A2 _12207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19337_ _19521_/A _19512_/A _19334_/X _19336_/X vssd1 vssd1 vccd1 vccd1 _19337_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_16549_ _16624_/A _16608_/A vssd1 vssd1 vccd1 vccd1 _16605_/A sky130_fd_sc_hd__nand2_1
XFILLER_149_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19268_ _19296_/A _19434_/A _19434_/B vssd1 vssd1 vccd1 vccd1 _19268_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__16364__B1 _16369_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17561__C1 _21011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18219_ _18219_/A _18219_/B vssd1 vssd1 vccd1 vccd1 _18276_/A sky130_fd_sc_hd__nand2_1
X_19199_ _19199_/A _19199_/B _19199_/C vssd1 vssd1 vccd1 vccd1 _19200_/B sky130_fd_sc_hd__and3_1
XFILLER_102_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22831__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21230_ _21230_/A _21230_/B _21230_/C vssd1 vssd1 vccd1 vccd1 _21231_/A sky130_fd_sc_hd__nand3_1
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18656__A2 _19176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16930__B _17341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11777__D _11949_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21161_ _21165_/A _22947_/Q vssd1 vssd1 vccd1 vccd1 _21161_/X sky130_fd_sc_hd__and2_1
XFILLER_171_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18203__A _18203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20452__B _20452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20112_ _12928_/A _16039_/A _20110_/A _20110_/B _20096_/Y vssd1 vssd1 vccd1 vccd1
+ _20112_/X sky130_fd_sc_hd__o221a_1
XFILLER_160_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21092_ _21092_/A _21093_/A vssd1 vssd1 vccd1 vccd1 _21138_/A sky130_fd_sc_hd__or2b_1
XFILLER_113_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20043_ _20024_/A _20024_/B _20024_/C vssd1 vssd1 vccd1 vccd1 _20043_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12251__A _12251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17092__A1 _15888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15642__A2 _16720_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13653__A1 _21489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21994_ _21994_/A vssd1 vssd1 vccd1 vccd1 _22072_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16377__B _16377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ _20945_/A _20945_/B vssd1 vssd1 vccd1 vccd1 _20946_/B sky130_fd_sc_hd__nand2_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13082__A _22841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13513__C _13521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20876_ _20876_/A _20876_/B vssd1 vssd1 vccd1 vccd1 _20877_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11314__B _22955_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22615_ _22796_/Q input38/X _22619_/S vssd1 vssd1 vccd1 vccd1 _22616_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11967__B2 _11966_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22546_ _22546_/A vssd1 vssd1 vccd1 vccd1 _22765_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18895__A2 _18889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14905__A1 _15188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22477_ _22499_/A vssd1 vssd1 vccd1 vccd1 _22486_/S sky130_fd_sc_hd__clkbuf_2
X_12230_ _18228_/A _18228_/B _12230_/C vssd1 vssd1 vccd1 vccd1 _12231_/C sky130_fd_sc_hd__nand3_1
XFILLER_108_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16107__B1 _19000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21428_ _21700_/A _21701_/A _21426_/Y vssd1 vssd1 vccd1 vccd1 _21430_/A sky130_fd_sc_hd__o21ai_1
XFILLER_170_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12161_ _19016_/C vssd1 vssd1 vccd1 vccd1 _19490_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21359_ _21359_/A _21359_/B _21359_/C vssd1 vssd1 vccd1 vccd1 _21388_/A sky130_fd_sc_hd__nand3_1
XFILLER_190_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12092_ _12135_/B vssd1 vssd1 vccd1 vccd1 _19358_/D sky130_fd_sc_hd__buf_2
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22600__A0 _11430_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15920_ _15921_/A _16414_/A _15918_/X _15919_/X vssd1 vssd1 vccd1 vccd1 _15920_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19072__A2 _11380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12058__A2_N _11924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11352__C1 _11351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18280__B1 _19358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15851_ _15756_/X _15750_/Y _15845_/X _15846_/Y vssd1 vssd1 vccd1 vccd1 _15855_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_7_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _14802_/A _14802_/B _14802_/C vssd1 vssd1 vccd1 vccd1 _14822_/C sky130_fd_sc_hd__nand3_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18486__C _18691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18570_ _18570_/A vssd1 vssd1 vccd1 vccd1 _18575_/B sky130_fd_sc_hd__clkbuf_2
X_15782_ _15775_/B _15775_/C _15728_/X vssd1 vssd1 vccd1 vccd1 _15783_/C sky130_fd_sc_hd__a21o_1
XFILLER_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12994_ _12944_/X _12991_/X _12993_/X vssd1 vssd1 vccd1 vccd1 _12994_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17521_ _17523_/B _17523_/C _17523_/A vssd1 vssd1 vccd1 vccd1 _17585_/A sky130_fd_sc_hd__a21oi_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14733_ _14733_/A _14733_/B vssd1 vssd1 vccd1 vccd1 _14738_/B sky130_fd_sc_hd__nor2_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ _11945_/A _11945_/B vssd1 vssd1 vccd1 vccd1 _11947_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17452_ _17452_/A _17457_/C _17457_/D vssd1 vssd1 vccd1 vccd1 _17454_/B sky130_fd_sc_hd__nand3_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14664_ _14664_/A _14664_/B vssd1 vssd1 vccd1 vccd1 _14843_/C sky130_fd_sc_hd__xnor2_4
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _11371_/X _11393_/Y _11399_/Y vssd1 vssd1 vccd1 vccd1 _11883_/A sky130_fd_sc_hd__a21bo_1
XFILLER_33_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20818__A _20818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16403_ _16403_/A _16403_/B vssd1 vssd1 vccd1 vccd1 _16433_/C sky130_fd_sc_hd__nand2_1
XFILLER_177_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13615_ _13602_/Y _13605_/Y _13566_/X _13599_/Y vssd1 vssd1 vccd1 vccd1 _13616_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_60_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17383_ _15919_/X _17388_/A _17382_/Y vssd1 vssd1 vccd1 vccd1 _17383_/Y sky130_fd_sc_hd__o21ai_2
X_14595_ _15056_/B _14595_/B _15056_/A vssd1 vssd1 vccd1 vccd1 _14942_/C sky130_fd_sc_hd__nand3_2
XANTENNA__18335__A1 _11511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18335__B2 _18980_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22854__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19122_ _19122_/A _19122_/B _19122_/C vssd1 vssd1 vccd1 vccd1 _19122_/Y sky130_fd_sc_hd__nand3_1
X_16334_ _16316_/Y _16327_/Y _16333_/Y vssd1 vssd1 vccd1 vccd1 _16354_/A sky130_fd_sc_hd__o21ai_4
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13546_ _13546_/A _13546_/B vssd1 vssd1 vccd1 vccd1 _13550_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19053_ _15522_/X _15521_/X _15523_/X _18795_/A vssd1 vssd1 vccd1 vccd1 _19053_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14357__C1 _14356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16265_ _16265_/A _16265_/B vssd1 vssd1 vccd1 vccd1 _16272_/A sky130_fd_sc_hd__nand2_1
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20693__A2 _17007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13477_ _13470_/Y _13474_/X _13475_/Y _13476_/Y vssd1 vssd1 vccd1 vccd1 _13477_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18004_ _17960_/A _17960_/D _18045_/B _18048_/B _18048_/A vssd1 vssd1 vccd1 vccd1
+ _18055_/B sky130_fd_sc_hd__a32o_1
X_15216_ _15216_/A vssd1 vssd1 vccd1 vccd1 _15217_/C sky130_fd_sc_hd__inv_2
XFILLER_126_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12428_ _20359_/A _12428_/B _20359_/C vssd1 vssd1 vccd1 vccd1 _12428_/Y sky130_fd_sc_hd__nor3_2
X_16196_ _16195_/A _16195_/B _16195_/C vssd1 vssd1 vccd1 vccd1 _16196_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__20553__A _20553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15147_ _15186_/A _15149_/A _15121_/X _15123_/X _15146_/Y vssd1 vssd1 vccd1 vccd1
+ _15148_/A sky130_fd_sc_hd__a221oi_2
XFILLER_141_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12359_ _22821_/Q vssd1 vssd1 vccd1 vccd1 _12687_/B sky130_fd_sc_hd__buf_2
XANTENNA__18023__A _18023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_591 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19955_ _19955_/A _19955_/B vssd1 vssd1 vccd1 vccd1 _19959_/A sky130_fd_sc_hd__xnor2_1
XFILLER_99_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15078_ _15078_/A _15078_/B vssd1 vssd1 vccd1 vccd1 _15086_/A sky130_fd_sc_hd__nand2_1
XFILLER_142_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17862__A _22902_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18906_ _18904_/Y _18709_/C _18905_/Y _18722_/C vssd1 vssd1 vccd1 vccd1 _18907_/C
+ sky130_fd_sc_hd__a22oi_2
X_14029_ _14029_/A _14029_/B vssd1 vssd1 vccd1 vccd1 _14052_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12071__A _18830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19886_ _19976_/A _19893_/A vssd1 vssd1 vccd1 vccd1 _19887_/C sky130_fd_sc_hd__nand2_1
XFILLER_122_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13883__A1 _14722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18837_ _18722_/A _18722_/B _18721_/A _18723_/A vssd1 vssd1 vccd1 vccd1 _18837_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_1098 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_778 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16821__A1 _16014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15382__A _15389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18768_ _18768_/A _18768_/B _18768_/C vssd1 vssd1 vccd1 vccd1 _18779_/B sky130_fd_sc_hd__nand3_2
XFILLER_67_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17719_ _17719_/A _17719_/B _17719_/C vssd1 vssd1 vccd1 vccd1 _17720_/B sky130_fd_sc_hd__nor3_1
XANTENNA__13813__B1_N _13826_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18699_ _18699_/A _18699_/B vssd1 vssd1 vccd1 vccd1 _19329_/A sky130_fd_sc_hd__nand2_4
XANTENNA__11415__A _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15388__A1 _15389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20730_ _20818_/B _20730_/B vssd1 vssd1 vccd1 vccd1 _20778_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20728__A _20728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16925__B _17386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20661_ _20658_/Y _20551_/Y _20659_/Y _20660_/Y vssd1 vssd1 vccd1 vccd1 _20827_/C
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_189_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18326__A1 _11904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13630__A _13630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22400_ _14369_/X input39/X _22402_/S vssd1 vssd1 vccd1 vccd1 _22401_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16644__C _16644_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20592_ _20593_/C _17281_/B _16708_/X _12928_/A vssd1 vssd1 vccd1 vccd1 _20595_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__17534__C1 _15960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22331_ _22309_/A _22309_/B _22329_/Y _22330_/Y _22313_/A vssd1 vssd1 vccd1 vccd1
+ _22333_/A sky130_fd_sc_hd__o221a_1
XANTENNA__14348__C1 _14347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16352__A3 _17462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22662__B _22662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22262_ _22262_/A vssd1 vssd1 vccd1 vccd1 _22263_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_118_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15557__A _15557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21213_ _21213_/A vssd1 vssd1 vccd1 vccd1 _21724_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22193_ _22193_/A _22193_/B vssd1 vssd1 vccd1 vccd1 _22194_/B sky130_fd_sc_hd__xor2_1
XFILLER_117_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15312__A1 _11935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21144_ _21150_/A _21150_/B _21150_/C _21142_/A vssd1 vssd1 vccd1 vccd1 _21147_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_116_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_1_0_bq_clk_i_A clkbuf_3_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20592__A2_N _17281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22043__D1 _22176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21075_ _21076_/B _21076_/D vssd1 vssd1 vccd1 vccd1 _21075_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20026_ _20026_/A _20026_/B vssd1 vssd1 vccd1 vccd1 _20026_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__21294__A _22672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11885__B1 _11895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21725__C _22041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15615__A2 _16715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16819__C _20928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13805__A _22866_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21977_ _21977_/A _22036_/B _22036_/C vssd1 vssd1 vccd1 vccd1 _21977_/Y sky130_fd_sc_hd__nand3_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11970__D _18875_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22877__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _12112_/A vssd1 vssd1 vccd1 vccd1 _11731_/A sky130_fd_sc_hd__buf_2
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20928_ _20928_/A _20928_/B _20928_/C vssd1 vssd1 vccd1 vccd1 _20933_/A sky130_fd_sc_hd__and3_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21741__B _21741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15379__B2 _17111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20911__A3 _17460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _11656_/Y _11737_/A _11732_/A vssd1 vssd1 vccd1 vccd1 _18648_/B sky130_fd_sc_hd__a21boi_2
XFILLER_109_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20859_ _20860_/B _20860_/C _20689_/Y _20790_/Y vssd1 vssd1 vccd1 vccd1 _20866_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13400_ _13495_/A _13495_/B vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16554__C _16554_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20124__A1 _15504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14380_ _14380_/A vssd1 vssd1 vccd1 vccd1 _21169_/A sky130_fd_sc_hd__buf_2
XFILLER_23_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18868__A2 _18330_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11592_ _11592_/A vssd1 vssd1 vccd1 vccd1 _11647_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _13502_/D vssd1 vssd1 vccd1 vccd1 _21739_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22529_ _22529_/A vssd1 vssd1 vccd1 vccd1 _22757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_856 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16050_ _16613_/C _20745_/C _16130_/A _16051_/C vssd1 vssd1 vccd1 vccd1 _16050_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_157_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13262_ _13262_/A _13265_/A _13401_/A _13262_/D vssd1 vssd1 vccd1 vccd1 _13438_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA_input75_A x[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15001_ _15001_/A _15001_/B _15001_/C _15001_/D vssd1 vssd1 vccd1 vccd1 _15018_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_182_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12213_ _15440_/A vssd1 vssd1 vccd1 vccd1 _16473_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ _13144_/A _13097_/A _13158_/A vssd1 vssd1 vccd1 vccd1 _13376_/A sky130_fd_sc_hd__a21o_1
XANTENNA__17385__C _17385_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20092__B _20092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15303__A1 _11705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ _22794_/Q vssd1 vssd1 vccd1 vccd1 _18677_/C sky130_fd_sc_hd__clkinv_2
XANTENNA__16500__B1 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15303__B2 _12501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18778__A _18778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19740_ _19740_/A _19740_/B vssd1 vssd1 vccd1 vccd1 _19746_/C sky130_fd_sc_hd__nand2_1
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16952_ _15546_/A _17403_/A _12930_/A _18814_/A vssd1 vssd1 vccd1 vccd1 _16952_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_1_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12075_ _11924_/C _11924_/D _12070_/X _12074_/X vssd1 vssd1 vccd1 vccd1 _12075_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15903_ _20255_/C vssd1 vssd1 vccd1 vccd1 _15903_/X sky130_fd_sc_hd__clkbuf_4
X_19671_ _19880_/D vssd1 vssd1 vccd1 vccd1 _19761_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_103_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16883_ _16882_/X _16637_/Y _16638_/Y _16635_/A _16644_/C vssd1 vssd1 vccd1 vccd1
+ _16886_/B sky130_fd_sc_hd__a32oi_4
XFILLER_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16298__A _16450_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18622_ _18453_/X _18450_/B _18451_/B _18451_/A vssd1 vssd1 vccd1 vccd1 _18623_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_37_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _15834_/A vssd1 vssd1 vccd1 vccd1 _16414_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15633__C _16450_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _18553_/A _18553_/B _18553_/C vssd1 vssd1 vccd1 vccd1 _18554_/B sky130_fd_sc_hd__nand3_1
XFILLER_46_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _15682_/Y _15433_/A _15681_/C _15681_/D vssd1 vssd1 vccd1 vccd1 _15769_/B
+ sky130_fd_sc_hd__o211ai_1
X_12977_ _15776_/D vssd1 vssd1 vccd1 vccd1 _20134_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_79_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17504_ _17354_/Y _17503_/X _17361_/Y vssd1 vssd1 vccd1 vccd1 _17800_/D sky130_fd_sc_hd__a21oi_4
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11928_ _11832_/Y _11834_/Y _11838_/Y _11927_/Y vssd1 vssd1 vccd1 vccd1 _12087_/A
+ sky130_fd_sc_hd__o211a_1
X_14716_ _14716_/A _14716_/B _14716_/C vssd1 vssd1 vccd1 vccd1 _14717_/C sky130_fd_sc_hd__nand3_1
XFILLER_73_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15696_ _18848_/D _16912_/A _15997_/C _15696_/D vssd1 vssd1 vccd1 vccd1 _15696_/Y
+ sky130_fd_sc_hd__nand4_2
X_18484_ _18484_/A _18695_/A vssd1 vssd1 vccd1 vccd1 _18488_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16567__B1 _14369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12840__A2 _16708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ _17435_/A vssd1 vssd1 vccd1 vccd1 _17440_/A sky130_fd_sc_hd__buf_2
X_14647_ _14963_/C _14181_/C _14181_/A _14646_/Y vssd1 vssd1 vccd1 vccd1 _14651_/B
+ sky130_fd_sc_hd__a31o_1
X_11859_ _11859_/A vssd1 vssd1 vccd1 vccd1 _11859_/X sky130_fd_sc_hd__buf_4
XFILLER_61_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19505__B1 _17393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17366_ _17616_/C _17358_/Y _17365_/Y vssd1 vssd1 vccd1 vccd1 _17719_/A sky130_fd_sc_hd__o21ai_2
X_14578_ _14578_/A vssd1 vssd1 vccd1 vccd1 _14942_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_186_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19105_ _19106_/A _19106_/B _19103_/Y _19104_/X vssd1 vssd1 vccd1 vccd1 _19257_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_16317_ _15904_/X _15905_/X _20471_/A _20471_/B vssd1 vssd1 vccd1 vccd1 _16332_/B
+ sky130_fd_sc_hd__o211ai_4
X_13529_ _13213_/X _13050_/X _13520_/B _13520_/A vssd1 vssd1 vccd1 vccd1 _13529_/Y
+ sky130_fd_sc_hd__o22ai_1
X_17297_ _17262_/X _17266_/Y _17307_/B _17304_/B vssd1 vssd1 vccd1 vccd1 _17301_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12066__A _16106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16248_ _16940_/A vssd1 vssd1 vccd1 vccd1 _16248_/X sky130_fd_sc_hd__clkbuf_4
X_19036_ _18866_/Y _19013_/B _19012_/X vssd1 vssd1 vccd1 vccd1 _19037_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__15542__A1 _15538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22913__D _22913_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15377__A _15377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput103 _14424_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[29] sky130_fd_sc_hd__buf_2
Xoutput114 _22664_/Q vssd1 vssd1 vccd1 vccd1 y[0] sky130_fd_sc_hd__buf_2
X_16179_ _16179_/A vssd1 vssd1 vccd1 vccd1 _16179_/X sky130_fd_sc_hd__buf_4
Xoutput125 _22950_/Q vssd1 vssd1 vccd1 vccd1 y[9] sky130_fd_sc_hd__buf_2
XFILLER_142_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18688__A _18691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19938_ _19913_/A _19913_/B _19913_/C vssd1 vssd1 vccd1 vccd1 _19952_/B sky130_fd_sc_hd__o21ai_1
XFILLER_99_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20730__B _20730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19869_ _19836_/D _19836_/Y _19867_/X _19894_/A vssd1 vssd1 vccd1 vccd1 _19921_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18200__B _19351_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21900_ _21909_/A vssd1 vssd1 vccd1 vccd1 _22008_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22880_ _22916_/CLK input74/X vssd1 vssd1 vccd1 vccd1 _22880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21831_ _21922_/A _21831_/B vssd1 vssd1 vccd1 vccd1 _21832_/C sky130_fd_sc_hd__nand2_1
XFILLER_71_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16936__A _17631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15840__A _15840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21762_ _21762_/A _21762_/B vssd1 vssd1 vccd1 vccd1 _21846_/C sky130_fd_sc_hd__nand2_1
XFILLER_52_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20354__A1 _12988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20713_ _20718_/A _20713_/B vssd1 vssd1 vccd1 vccd1 _20720_/A sky130_fd_sc_hd__nor2_1
XFILLER_168_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21693_ _21688_/B _21693_/B _21693_/C vssd1 vssd1 vccd1 vccd1 _21837_/B sky130_fd_sc_hd__nand3b_1
XFILLER_178_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13360__A _13423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15781__A1 _20249_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20644_ _20638_/Y _20639_/X _20631_/Y _20737_/A vssd1 vssd1 vccd1 vccd1 _20645_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__20608__D _20917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20575_ _20734_/A _20575_/B _20637_/A _20870_/C vssd1 vssd1 vccd1 vccd1 _20575_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_149_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22314_ _22314_/A _22314_/B _22314_/C vssd1 vssd1 vccd1 vccd1 _22316_/A sky130_fd_sc_hd__nor3_1
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21289__A _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22245_ _22213_/Y _22216_/Y _22216_/B _22244_/Y vssd1 vssd1 vccd1 vccd1 _22245_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_133_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14191__A _14191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17286__A1 _11561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22176_ _22176_/A _22238_/A _22176_/C _22265_/B vssd1 vssd1 vccd1 vccd1 _22238_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__13519__B _13519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21127_ _21150_/A _21127_/B _21127_/C vssd1 vssd1 vccd1 vccd1 _21128_/B sky130_fd_sc_hd__and3_1
XANTENNA__19027__A2 _19023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13847__A1 _14013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21058_ _21095_/A vssd1 vssd1 vccd1 vccd1 _21058_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18110__B _18848_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12900_ _12900_/A _12900_/B _12900_/C vssd1 vssd1 vccd1 vccd1 _13011_/B sky130_fd_sc_hd__nand3_2
X_20009_ _20057_/A _20057_/B _20010_/A vssd1 vssd1 vccd1 vccd1 _20035_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__17007__A _17007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13880_ _13807_/A _13873_/A _14808_/C _13808_/Y vssd1 vssd1 vccd1 vccd1 _13920_/A
+ sky130_fd_sc_hd__a31o_1
X_12831_ _20213_/A vssd1 vssd1 vccd1 vccd1 _20092_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18538__A1 _16921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15550_ _19507_/B vssd1 vssd1 vccd1 vccd1 _19687_/B sky130_fd_sc_hd__clkbuf_4
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _13022_/A _12761_/X _12757_/B vssd1 vssd1 vccd1 vccd1 _12763_/B sky130_fd_sc_hd__o21ai_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_634 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14499_/Y _14607_/B _14492_/Y _14497_/Y vssd1 vssd1 vccd1 vccd1 _14501_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11718_/A _11713_/B vssd1 vssd1 vccd1 vccd1 _11714_/A sky130_fd_sc_hd__nand2_2
XFILLER_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15481_/A _22660_/B _22662_/B vssd1 vssd1 vccd1 vccd1 _15482_/D sky130_fd_sc_hd__nor3_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12693_ _15394_/A vssd1 vssd1 vccd1 vccd1 _17246_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14366__A _22764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17220_/A _17220_/B vssd1 vssd1 vccd1 vccd1 _17225_/A sky130_fd_sc_hd__xor2_1
X_14432_ _14432_/A vssd1 vssd1 vccd1 vccd1 _18259_/B sky130_fd_sc_hd__buf_4
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11644_ _11644_/A _11645_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _11644_/X sky130_fd_sc_hd__and3_1
XANTENNA__15772__A1 _15350_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15772__B2 _15389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17151_ _17168_/A vssd1 vssd1 vccd1 vccd1 _17180_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14363_ _18128_/C _14354_/X _14355_/X _14361_/X _14362_/X vssd1 vssd1 vccd1 vccd1
+ _14363_/X sky130_fd_sc_hd__a32o_1
XFILLER_168_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 wb_adr_i[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
X_11575_ _11899_/A _11899_/B vssd1 vssd1 vccd1 vccd1 _11576_/B sky130_fd_sc_hd__and2_1
XFILLER_183_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput27 wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16102_ _16103_/D _20452_/A _20452_/B _16150_/A _16103_/C vssd1 vssd1 vccd1 vccd1
+ _16113_/C sky130_fd_sc_hd__a32o_1
XFILLER_183_642 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ _13314_/A _13314_/B _13314_/C vssd1 vssd1 vccd1 vccd1 _13354_/A sky130_fd_sc_hd__nand3_1
Xinput38 wb_dat_i[12] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_2
X_17082_ _17081_/A _17591_/B _16098_/X _17007_/A vssd1 vssd1 vccd1 vccd1 _17082_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput49 wb_dat_i[22] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14294_ _14843_/A vssd1 vssd1 vccd1 vccd1 _22672_/D sky130_fd_sc_hd__inv_2
XANTENNA__15909__B _16192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16033_ _16034_/A _16210_/A _16034_/C vssd1 vssd1 vccd1 vccd1 _16035_/A sky130_fd_sc_hd__a21o_1
XFILLER_109_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ _13230_/X _13623_/A _21584_/C _13257_/B vssd1 vssd1 vccd1 vccd1 _13273_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_109_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17277__A1 _14431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13176_ _13176_/A vssd1 vssd1 vccd1 vccd1 _13633_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_97_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ _12127_/A _12130_/A _18338_/C vssd1 vssd1 vccd1 vccd1 _18141_/A sky130_fd_sc_hd__nand3_1
XFILLER_97_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19018__A2 _19015_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20820__A2 _20748_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17984_ _19419_/B _18030_/B _18030_/C _18030_/D vssd1 vssd1 vccd1 vccd1 _17987_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19723_ _19723_/A _19723_/B vssd1 vssd1 vccd1 vccd1 _19735_/B sky130_fd_sc_hd__nand2_1
X_16935_ _19587_/C vssd1 vssd1 vccd1 vccd1 _19694_/B sky130_fd_sc_hd__clkbuf_4
X_12058_ _12079_/C _11924_/X _11897_/Y _11900_/Y vssd1 vssd1 vccd1 vccd1 _12061_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_96_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16237__C1 _19047_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19654_ _19652_/A _19652_/B _19740_/A _19656_/B vssd1 vssd1 vccd1 vccd1 _19658_/A
+ sky130_fd_sc_hd__o211a_1
X_16866_ _16866_/A _16866_/B _16866_/C _16866_/D vssd1 vssd1 vccd1 vccd1 _16867_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__16788__B1 _12294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15363__C _15363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18605_ _18432_/A _18603_/Y _18604_/Y vssd1 vssd1 vccd1 vccd1 _18606_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__16252__A2 _15546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15817_ _15817_/A _15825_/A vssd1 vssd1 vccd1 vccd1 _15819_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19585_ _19602_/A _19602_/B _19602_/C _19585_/D vssd1 vssd1 vccd1 vccd1 _19607_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_19_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16797_ _16834_/A vssd1 vssd1 vccd1 vccd1 _16845_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18536_ _14430_/A _15297_/A _15559_/B _18328_/B _18328_/C vssd1 vssd1 vccd1 vccd1
+ _18536_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _15748_/A _15748_/B vssd1 vssd1 vccd1 vccd1 _15755_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_751 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ _18455_/Y _18296_/B _18466_/Y _18289_/Y vssd1 vssd1 vccd1 vccd1 _18467_/Y
+ sky130_fd_sc_hd__o211ai_4
X_15679_ _15859_/C _15679_/B vssd1 vssd1 vccd1 vccd1 _15680_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17418_ _17399_/Y _17410_/A _17550_/A _17550_/B vssd1 vssd1 vccd1 vccd1 _17420_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18398_ _18407_/A _18407_/B _18397_/Y vssd1 vssd1 vccd1 vccd1 _18398_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_21_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18690__B _18690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13774__B1 _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20639__A2 _20178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17349_ _17341_/X _17338_/X _17330_/Y _17337_/X vssd1 vssd1 vccd1 vccd1 _17350_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_14_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20360_ _20368_/A _20370_/D _20359_/X vssd1 vssd1 vccd1 vccd1 _20360_/X sky130_fd_sc_hd__a21o_1
XFILLER_162_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19019_ _17421_/A _17422_/A _18512_/B _18512_/C vssd1 vssd1 vccd1 vccd1 _19020_/B
+ sky130_fd_sc_hd__a211o_1
X_20291_ _20294_/B vssd1 vssd1 vccd1 vccd1 _20298_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__11508__B1_N _11507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22030_ _22030_/A _22030_/B vssd1 vssd1 vccd1 vccd1 _22031_/C sky130_fd_sc_hd__nand2_1
XFILLER_103_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15818__A2 _15727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14161__D _14494_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16369__C _16369_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22932_ _22933_/CLK _22932_/D vssd1 vssd1 vccd1 vccd1 _22932_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18865__B _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13074__B _13519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22863_ _22944_/CLK _22863_/D vssd1 vssd1 vccd1 vccd1 _22863_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14254__A1 _14220_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16666__A _16669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19178__D1 _19687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19042__A _19418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21814_ _21814_/A _21814_/B _21913_/B _21814_/D vssd1 vssd1 vccd1 vccd1 _21837_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_97_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22794_ _22795_/CLK _22794_/D vssd1 vssd1 vccd1 vccd1 _22794_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_189_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19193__A1 _19504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21745_ _21850_/A vssd1 vssd1 vccd1 vccd1 _22176_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13090__A _22843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11603__A _12003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14557__A2 _14843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21676_ _21680_/B _21676_/B _21676_/C vssd1 vssd1 vccd1 vccd1 _21809_/A sky130_fd_sc_hd__nand3b_2
XFILLER_178_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11322__B _22953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22915__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20627_ _20598_/X _20599_/Y _20484_/Y vssd1 vssd1 vccd1 vccd1 _20629_/B sky130_fd_sc_hd__o21ai_2
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11360_ _12008_/A vssd1 vssd1 vccd1 vccd1 _11361_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20558_ _22933_/Q _20566_/A _20566_/B vssd1 vssd1 vccd1 vccd1 _20559_/B sky130_fd_sc_hd__or3_1
XANTENNA__18105__B _18848_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11291_ _11404_/B _11404_/C _11411_/A _11325_/A vssd1 vssd1 vccd1 vccd1 _11295_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_152_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20489_ _20465_/X _20470_/Y _20499_/D vssd1 vssd1 vccd1 vccd1 _20489_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_106_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12725__D1 _12601_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13030_ _12990_/B _13036_/A _12990_/D _12990_/A vssd1 vssd1 vccd1 vccd1 _13031_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_1130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22228_ _22228_/A _22263_/C vssd1 vssd1 vccd1 vccd1 _22271_/A sky130_fd_sc_hd__or2_1
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15809__A2 _12774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11543__A2 _18371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22159_ _22164_/A _22159_/B vssd1 vssd1 vccd1 vccd1 _22160_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_1147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20370__B _20593_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15464__B _16256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A wb_dat_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14981_ _14980_/A _15035_/B _14980_/C vssd1 vssd1 vccd1 vccd1 _14981_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16219__C1 _18193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14493__A1 _14491_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16720_ _20781_/A _20781_/B _16720_/C vssd1 vssd1 vccd1 vccd1 _16720_/Y sky130_fd_sc_hd__nand3_1
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13932_ _22873_/Q vssd1 vssd1 vccd1 vccd1 _14624_/A sky130_fd_sc_hd__clkinv_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16651_ _15646_/X _15645_/X _16431_/B _16444_/A vssd1 vssd1 vccd1 vccd1 _16652_/B
+ sky130_fd_sc_hd__o211ai_2
X_13863_ _13829_/B _13877_/A _13807_/A _13837_/A vssd1 vssd1 vccd1 vccd1 _13866_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15602_ _15449_/X _15505_/X _15502_/C vssd1 vssd1 vccd1 vccd1 _15602_/X sky130_fd_sc_hd__o21a_1
X_12814_ _15633_/B _16450_/C _20341_/C vssd1 vssd1 vccd1 vccd1 _20219_/A sky130_fd_sc_hd__nand3_4
XFILLER_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19370_ _19356_/X _19363_/Y _19369_/Y vssd1 vssd1 vccd1 vccd1 _19379_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__15993__A1 _15904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16582_ _16582_/A vssd1 vssd1 vccd1 vccd1 _16585_/A sky130_fd_sc_hd__clkbuf_2
X_13794_ _13793_/Y _13773_/A _22757_/Q vssd1 vssd1 vccd1 vccd1 _13959_/A sky130_fd_sc_hd__a21o_2
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20098__A _20478_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18321_ _19011_/A vssd1 vssd1 vccd1 vccd1 _19194_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15533_ _15439_/X _15524_/X _15527_/A vssd1 vssd1 vccd1 vccd1 _16215_/A sky130_fd_sc_hd__o21ai_2
XFILLER_16_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13712__B _15114_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12745_ _12745_/A _12745_/B _12745_/C vssd1 vssd1 vccd1 vccd1 _12745_/Y sky130_fd_sc_hd__nand3_1
XFILLER_187_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15630__D _16361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12609__A _20461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17734__A2 _17928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _18251_/A _18257_/B _19443_/A _12258_/A _18251_/Y vssd1 vssd1 vccd1 vccd1
+ _18252_/Y sky130_fd_sc_hd__o221ai_2
X_15464_ _16256_/A _16256_/B _15466_/B _15466_/C vssd1 vssd1 vccd1 vccd1 _15472_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _16256_/C vssd1 vssd1 vccd1 vccd1 _16932_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_31_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17203_ _17036_/A _17036_/C _17036_/B vssd1 vssd1 vccd1 vccd1 _17205_/A sky130_fd_sc_hd__a21bo_1
X_14415_ _22713_/Q _14403_/X _14410_/X _22745_/Q _14414_/X vssd1 vssd1 vccd1 vccd1
+ _14415_/X sky130_fd_sc_hd__a221o_1
X_11627_ _11627_/A vssd1 vssd1 vccd1 vccd1 _18716_/A sky130_fd_sc_hd__buf_2
X_18183_ _18173_/C _18173_/B _18173_/A vssd1 vssd1 vccd1 vccd1 _18183_/Y sky130_fd_sc_hd__a21oi_4
X_15395_ _20323_/A vssd1 vssd1 vccd1 vccd1 _17128_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_168_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17134_ _17134_/A vssd1 vssd1 vccd1 vccd1 _17288_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_128_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14346_ _12320_/A _14344_/X _14337_/X _13095_/X _14345_/X vssd1 vssd1 vccd1 vccd1
+ _14346_/X sky130_fd_sc_hd__a221o_1
X_11558_ _15435_/C vssd1 vssd1 vccd1 vccd1 _11659_/D sky130_fd_sc_hd__inv_2
XFILLER_129_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17065_ _17065_/A vssd1 vssd1 vccd1 vccd1 _17373_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14277_ _14279_/B _14280_/A _14277_/C vssd1 vssd1 vccd1 vccd1 _14280_/B sky130_fd_sc_hd__nand3_1
XFILLER_195_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11489_ _12157_/A _12158_/A vssd1 vssd1 vccd1 vccd1 _18167_/A sky130_fd_sc_hd__nand2_1
X_16016_ _16016_/A vssd1 vssd1 vccd1 vccd1 _16016_/X sky130_fd_sc_hd__buf_4
XFILLER_143_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13228_ _22848_/Q vssd1 vssd1 vccd1 vccd1 _13229_/A sky130_fd_sc_hd__inv_2
XFILLER_143_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14720__A2 _14942_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19772__D _19772_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13161_/A _21336_/C _13161_/C vssd1 vssd1 vccd1 vccd1 _13162_/A sky130_fd_sc_hd__a21oi_4
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15374__B _15382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17967_ _17967_/A _22904_/Q _17967_/C vssd1 vssd1 vccd1 vccd1 _17968_/B sky130_fd_sc_hd__and3_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17292__D _20793_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14484__A1 _13737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19706_ _19708_/A _19708_/B _19789_/A vssd1 vssd1 vccd1 vccd1 _19706_/X sky130_fd_sc_hd__and3_1
XFILLER_84_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16918_ _16911_/X _16913_/X _16915_/Y _17525_/C _19619_/B vssd1 vssd1 vccd1 vccd1
+ _16919_/C sky130_fd_sc_hd__o2111ai_4
X_17898_ _17897_/A _17897_/B _17897_/C vssd1 vssd1 vccd1 vccd1 _17899_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19637_ _19486_/A _19486_/B _19536_/D _19536_/C vssd1 vssd1 vccd1 vccd1 _19637_/Y
+ sky130_fd_sc_hd__o211ai_4
X_16849_ _16742_/Y _16743_/X _16747_/X vssd1 vssd1 vccd1 vccd1 _16849_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16486__A _17139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19568_ _19669_/A _19669_/B _19569_/A _19750_/A vssd1 vssd1 vccd1 vccd1 _19571_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15984__A1 _15427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15984__B2 _15983_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13444__C1 _13475_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16613__A_N _16351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18519_ _18915_/A _18526_/D _18916_/A vssd1 vssd1 vccd1 vccd1 _18519_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__22938__CLK _22948_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19499_ _19350_/X _16799_/X _19497_/A vssd1 vssd1 vccd1 vccd1 _19503_/A sky130_fd_sc_hd__o21ai_1
XFILLER_90_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19012__D _19012_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21530_ _21530_/A vssd1 vssd1 vccd1 vccd1 _21531_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11744__A1_N _11904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21461_ _21651_/B vssd1 vssd1 vccd1 vccd1 _21514_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17748__C _20917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17110__A _17110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20412_ _20408_/Y _20409_/Y _20410_/Y _20411_/Y vssd1 vssd1 vccd1 vccd1 _20413_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_105_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21392_ _21393_/A _21393_/B _21378_/A _21378_/B vssd1 vssd1 vccd1 vccd1 _21404_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_190_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11773__A2 _11771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20343_ _20343_/A _20464_/A vssd1 vssd1 vccd1 vccd1 _20343_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20274_ _20202_/Y _20270_/Y _20272_/Y _20273_/X vssd1 vssd1 vccd1 vccd1 _20274_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20471__A _20471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20245__B1 _16477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12722__A1 _12716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22013_ _22013_/A _22013_/B vssd1 vssd1 vccd1 vccd1 _22014_/B sky130_fd_sc_hd__and2_1
XANTENNA__12722__B2 _12721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22915_ _22915_/CLK _22915_/D vssd1 vssd1 vccd1 vccd1 _22915_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18610__B1 _15530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21733__C _22108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16396__A _20975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12238__B1 _18778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22846_ _22943_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 _22846_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22777_ _22810_/CLK _22777_/D vssd1 vssd1 vccd1 vccd1 _22777_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12771_/A _12773_/A vssd1 vssd1 vccd1 vccd1 _12553_/A sky130_fd_sc_hd__nor2_1
XFILLER_158_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21728_ _21629_/Y _21725_/Y _21724_/Y _21455_/X vssd1 vssd1 vccd1 vccd1 _21728_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_52_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20646__A _20870_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12461_ _12461_/A vssd1 vssd1 vccd1 vccd1 _15569_/A sky130_fd_sc_hd__buf_2
XFILLER_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21659_ _21651_/X _21666_/A _21515_/Y vssd1 vssd1 vccd1 vccd1 _21659_/X sky130_fd_sc_hd__a21o_1
X_14200_ _14200_/A vssd1 vssd1 vccd1 vccd1 _14693_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__18116__A _18116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ _11436_/A _16482_/A _11407_/B vssd1 vssd1 vccd1 vccd1 _11464_/A sky130_fd_sc_hd__a21o_1
XFILLER_32_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1094 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22473__A1 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15180_ _15180_/A _15180_/B vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__nand2_1
XFILLER_149_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14950__A2 _14013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12410__B1 _15325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ _12487_/B _12487_/C _12391_/Y vssd1 vssd1 vccd1 vccd1 _12407_/A sky130_fd_sc_hd__a21o_1
XFILLER_126_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ _14686_/B vssd1 vssd1 vccd1 vccd1 _14131_/X sky130_fd_sc_hd__buf_2
XFILLER_137_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11343_ _22788_/Q _11496_/B vssd1 vssd1 vccd1 vccd1 _11471_/C sky130_fd_sc_hd__nand2_2
XFILLER_152_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16152__A1 _15904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16152__B2 _12774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ _14169_/A _14169_/B _14058_/X _14061_/X vssd1 vssd1 vccd1 vccd1 _14167_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_11274_ _22799_/Q vssd1 vssd1 vccd1 vccd1 _11995_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13013_ _13011_/A _13011_/B _12966_/B _13012_/Y vssd1 vssd1 vccd1 vccd1 _13040_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18870_ _18839_/X _18865_/X _18909_/A vssd1 vssd1 vccd1 vccd1 _18870_/Y sky130_fd_sc_hd__o21ai_1
X_17821_ _19896_/A _17886_/A _17821_/C _17833_/A vssd1 vssd1 vccd1 vccd1 _17886_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__16455__A2 _15531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18786__A _22913_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__B _12938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
X_17752_ _19844_/B _17752_/B _17752_/C _20972_/B vssd1 vssd1 vccd1 vccd1 _17753_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_130_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14964_ _13737_/X _13746_/X _14670_/A vssd1 vssd1 vccd1 vccd1 _14966_/B sky130_fd_sc_hd__a21o_1
X_16703_ _16889_/B _16673_/A _16665_/A vssd1 vssd1 vccd1 vccd1 _16892_/A sky130_fd_sc_hd__a21o_1
XANTENNA__17404__A1 _15903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17404__B2 _16177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13915_ _13924_/A _14618_/A _13937_/A _13903_/Y vssd1 vssd1 vccd1 vccd1 _14021_/B
+ sky130_fd_sc_hd__o211ai_2
X_17683_ _17687_/A _17687_/B _17687_/C vssd1 vssd1 vccd1 vccd1 _17683_/X sky130_fd_sc_hd__and3_1
X_14895_ _14895_/A _14895_/B _14895_/C vssd1 vssd1 vccd1 vccd1 _14965_/A sky130_fd_sc_hd__nand3_1
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19422_ _19422_/A _19556_/A vssd1 vssd1 vccd1 vccd1 _19424_/A sky130_fd_sc_hd__nand2_1
X_16634_ _16634_/A _16634_/B _16634_/C vssd1 vssd1 vccd1 vccd1 _16635_/A sky130_fd_sc_hd__nand3_2
XFILLER_63_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13846_ _13985_/B vssd1 vssd1 vccd1 vccd1 _14013_/B sky130_fd_sc_hd__buf_2
XANTENNA__21362__D _21724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19353_ _19507_/A _19353_/B _19353_/C vssd1 vssd1 vccd1 vccd1 _19368_/B sky130_fd_sc_hd__and3_1
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13442__B _13475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13777_ _14184_/A _14184_/B vssd1 vssd1 vccd1 vccd1 _14042_/A sky130_fd_sc_hd__nand2_1
X_16565_ _15617_/X _16323_/D _16580_/A vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__a21oi_1
XFILLER_188_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18304_ _18305_/A _18305_/D _18459_/A vssd1 vssd1 vccd1 vccd1 _18572_/A sky130_fd_sc_hd__a21o_1
X_15516_ _15755_/A _15439_/X _15448_/X vssd1 vssd1 vccd1 vccd1 _15516_/Y sky130_fd_sc_hd__o21ai_1
X_19284_ _19284_/A _19284_/B vssd1 vssd1 vccd1 vccd1 _19681_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12728_ _20207_/C _15314_/A vssd1 vssd1 vccd1 vccd1 _20096_/A sky130_fd_sc_hd__nand2_1
X_16496_ _16496_/A vssd1 vssd1 vccd1 vccd1 _16496_/X sky130_fd_sc_hd__buf_2
XFILLER_30_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16753__B _16753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18235_ _18249_/A _12249_/A _18231_/Y _18234_/X vssd1 vssd1 vccd1 vccd1 _18251_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_30_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15447_ _19047_/B vssd1 vssd1 vccd1 vccd1 _19694_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_787 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12659_ _16157_/C _20723_/A _12757_/B vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__and3_1
XANTENNA__18026__A _19945_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22464__A1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18668__B1 _15580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18166_ _18172_/A _18383_/B _18132_/Y _18136_/X vssd1 vssd1 vccd1 vccd1 _18173_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_11_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15378_ _15378_/A vssd1 vssd1 vccd1 vccd1 _17111_/A sky130_fd_sc_hd__buf_4
XANTENNA__14273__B _14575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ _20781_/A vssd1 vssd1 vccd1 vccd1 _21019_/A sky130_fd_sc_hd__buf_2
XFILLER_144_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14329_ _14413_/A vssd1 vssd1 vccd1 vccd1 _14361_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18097_ _18092_/Y _18093_/Y _18849_/D _18096_/Y _18810_/A vssd1 vssd1 vccd1 vccd1
+ _18098_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_116_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17048_ _17076_/A _17076_/B _17076_/C _17048_/D vssd1 vssd1 vccd1 vccd1 _17048_/Y
+ sky130_fd_sc_hd__nand4_4
XANTENNA__22921__D _22921_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11507__A2 _11503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12180__A2 _12168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18999_ _18999_/A vssd1 vssd1 vccd1 vccd1 _19614_/C sky130_fd_sc_hd__buf_2
XFILLER_39_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_6_0_bq_clk_i_A clkbuf_3_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21727__B1 _21733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18199__A2 _11503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20961_ _20961_/A _20961_/B _22937_/Q vssd1 vssd1 vccd1 vccd1 _20961_/Y sky130_fd_sc_hd__nand3_1
X_22700_ _22733_/CLK _22700_/D vssd1 vssd1 vccd1 vccd1 _22700_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13633__A _13633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20892_ _20892_/A _20892_/B vssd1 vssd1 vccd1 vccd1 _20892_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22631_ _22631_/A vssd1 vssd1 vccd1 vccd1 _22803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19320__A _19320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22562_ _22562_/A vssd1 vssd1 vccd1 vccd1 _22772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21513_ _21464_/X _21465_/Y _21507_/Y _21512_/Y vssd1 vssd1 vccd1 vccd1 _21537_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_167_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22493_ _22742_/Q input49/X _22497_/S vssd1 vssd1 vccd1 vccd1 _22494_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21444_ _22172_/A vssd1 vssd1 vccd1 vccd1 _22231_/D sky130_fd_sc_hd__buf_2
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21375_ _21177_/Y _21179_/B _21374_/Y vssd1 vssd1 vccd1 vccd1 _21378_/A sky130_fd_sc_hd__a21oi_2
XFILLER_135_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20326_ _12577_/X _12576_/X _20323_/D _17532_/A vssd1 vssd1 vccd1 vccd1 _20326_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_123_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22831__D _22843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20257_ _20262_/C _20262_/B _20262_/A vssd1 vssd1 vccd1 vccd1 _20261_/A sky130_fd_sc_hd__a21oi_4
XFILLER_103_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20188_ _20064_/Y _13045_/Y _20186_/Y vssd1 vssd1 vccd1 vccd1 _20189_/C sky130_fd_sc_hd__a21o_1
XFILLER_130_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11961_ _12219_/A _12220_/A vssd1 vssd1 vccd1 vccd1 _11963_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_982 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17398__B1 _17643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22391__A0 _12378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12474__A3 _12528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_610 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _14808_/D vssd1 vssd1 vccd1 vccd1 _15115_/C sky130_fd_sc_hd__buf_2
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14948_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15948__A1 _15937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ _17313_/D _19455_/C _16130_/B _18305_/B vssd1 vssd1 vccd1 vccd1 _11909_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13631_ _21399_/A _21489_/A _13630_/Y _13595_/Y vssd1 vssd1 vccd1 vccd1 _13666_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22829_ _22850_/CLK _22841_/Q vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14620__A1 _14942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13562_ _13614_/A _13539_/A _13614_/C vssd1 vssd1 vccd1 vccd1 _13608_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__21497__A2 _21220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16350_ _20582_/A vssd1 vssd1 vccd1 vccd1 _17462_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_160_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19587__D _19587_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15301_ _16257_/A _16257_/B _15893_/C vssd1 vssd1 vccd1 vccd1 _15302_/B sky130_fd_sc_hd__nand3_2
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12513_ _12513_/A _22690_/Q vssd1 vssd1 vccd1 vccd1 _12525_/B sky130_fd_sc_hd__nand2_4
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16281_ _16283_/A _16283_/B vssd1 vssd1 vccd1 vccd1 _16288_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13493_ _13493_/A _13493_/B vssd1 vssd1 vccd1 vccd1 _21280_/B sky130_fd_sc_hd__nand2_1
XFILLER_185_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20095__B _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18020_ _18020_/A _18020_/B _18020_/C _18020_/D vssd1 vssd1 vccd1 vccd1 _18042_/A
+ sky130_fd_sc_hd__nor4_2
XFILLER_145_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12444_ _15466_/C vssd1 vssd1 vccd1 vccd1 _15799_/B sky130_fd_sc_hd__buf_2
X_15232_ _15180_/A _15205_/C _15180_/B _14552_/X vssd1 vssd1 vccd1 vccd1 _15233_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19311__A1 _18514_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ _15163_/A _15163_/B _15163_/C vssd1 vssd1 vccd1 vccd1 _15163_/X sky130_fd_sc_hd__or3_1
XANTENNA__13592__D1 _21445_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ _12519_/B vssd1 vssd1 vccd1 vccd1 _15608_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_181_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17322__B1 _17125_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ _14111_/X _14191_/B _14491_/C _14113_/X vssd1 vssd1 vccd1 vccd1 _14115_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11326_ _11324_/X _11315_/B _11325_/Y vssd1 vssd1 vccd1 vccd1 _11372_/A sky130_fd_sc_hd__o21ai_2
X_19971_ _19976_/B _19971_/B vssd1 vssd1 vccd1 vccd1 _19972_/B sky130_fd_sc_hd__and2_1
XFILLER_114_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15094_ _15034_/A _15033_/B _15033_/A vssd1 vssd1 vccd1 vccd1 _15095_/C sky130_fd_sc_hd__o21bai_1
XFILLER_153_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14687__A1 _14998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21638__C _21638_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18922_ _18908_/C _18908_/B _18920_/Y _18921_/X vssd1 vssd1 vccd1 vccd1 _18922_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_14045_ _14044_/B _14273_/C _14044_/C _14044_/A vssd1 vssd1 vccd1 vccd1 _14045_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18853_ _18853_/A vssd1 vssd1 vccd1 vccd1 _18920_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15636__B1 _16720_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17804_ _19844_/D vssd1 vssd1 vccd1 vccd1 _19901_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_94_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15933__A _15933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18784_ _18607_/Y _19281_/A _19138_/D vssd1 vssd1 vccd1 vccd1 _18969_/A sky130_fd_sc_hd__a21oi_1
X_15996_ _15797_/X _15546_/X _16006_/A vssd1 vssd1 vccd1 vccd1 _16000_/A sky130_fd_sc_hd__o21ai_1
XFILLER_95_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17735_ _17638_/X _17734_/X _17633_/Y vssd1 vssd1 vccd1 vccd1 _17736_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__18666__D _19507_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14947_ _14947_/A _14947_/B _14947_/C _14947_/D vssd1 vssd1 vccd1 vccd1 _14959_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_684 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17666_ _17661_/A _17661_/B _17660_/A _17660_/B vssd1 vssd1 vccd1 vccd1 _17666_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11673__B2 _18666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14878_ _14881_/A _14952_/B _14947_/A _14887_/B vssd1 vssd1 vccd1 vccd1 _14883_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20932__A1 _17928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16061__B1 _11845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19405_ _19254_/A _19254_/B _19254_/C _19149_/X vssd1 vssd1 vccd1 vccd1 _19405_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_91_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16617_ _16617_/A _16873_/A _16617_/C _16617_/D vssd1 vssd1 vccd1 vccd1 _16873_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__16600__A2 _16310_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13829_ _13829_/A _13829_/B vssd1 vssd1 vccd1 vccd1 _13829_/Y sky130_fd_sc_hd__nand2_2
X_17597_ _17597_/A _17597_/B _17597_/C vssd1 vssd1 vccd1 vccd1 _17704_/A sky130_fd_sc_hd__nand3_2
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19336_ _19336_/A _19619_/D _19768_/B _19771_/A vssd1 vssd1 vccd1 vccd1 _19336_/X
+ sky130_fd_sc_hd__and4_2
X_16548_ _16548_/A _16548_/B _16548_/C vssd1 vssd1 vccd1 vccd1 _16608_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12622__B1 _12601_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22916__D _22916_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20696__B1 _16996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19267_ _19272_/C vssd1 vssd1 vccd1 vccd1 _19434_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16364__A1 _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16479_ _16479_/A vssd1 vssd1 vccd1 vccd1 _16479_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17561__B1 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18218_ _18417_/B vssd1 vssd1 vccd1 vccd1 _18219_/B sky130_fd_sc_hd__inv_2
XANTENNA__11701__A _11819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22437__A1 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19198_ _19059_/Y _19215_/A _18282_/X _19194_/Y vssd1 vssd1 vccd1 vccd1 _19200_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18149_ _18348_/A _19016_/B _19016_/C vssd1 vssd1 vccd1 vccd1 _18150_/B sky130_fd_sc_hd__and3_1
XFILLER_8_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18656__A3 _18514_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16930__C _16930_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12235__C _22660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21160_ _21165_/A _22948_/Q vssd1 vssd1 vccd1 vccd1 _21164_/B sky130_fd_sc_hd__and2_1
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18203__B _18203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20111_ _16778_/X _16779_/X _20109_/Y _20110_/Y _20593_/D vssd1 vssd1 vccd1 vccd1
+ _20111_/X sky130_fd_sc_hd__o221a_1
XFILLER_131_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12532__A _12532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21091_ _21091_/A _21091_/B vssd1 vssd1 vccd1 vccd1 _21093_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20042_ _20022_/A _20042_/B _20042_/C vssd1 vssd1 vccd1 vccd1 _20042_/Y sky130_fd_sc_hd__nand3b_1
XANTENNA__18813__B1 _18812_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17092__A2 _17435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15642__A3 _16809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21993_ _21993_/A _22029_/B vssd1 vssd1 vccd1 vccd1 _21996_/C sky130_fd_sc_hd__nand2_1
XFILLER_67_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20944_ _20877_/A _20877_/B _20876_/B vssd1 vssd1 vccd1 vccd1 _20946_/A sky130_fd_sc_hd__a21oi_1
XFILLER_54_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21580__A _21580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20875_ _20871_/B _20871_/A _20873_/X _20874_/Y vssd1 vssd1 vccd1 vccd1 _20876_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__13513__D _13519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22614_ _22614_/A vssd1 vssd1 vccd1 vccd1 _22795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22545_ _22765_/Q input39/X _22547_/S vssd1 vssd1 vccd1 vccd1 _22546_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12707__A _12938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18895__A3 _18890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22476_ _22476_/A vssd1 vssd1 vccd1 vccd1 _22734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22615__S _22619_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16107__A1 _16106_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21427_ _21297_/Y _21420_/X _21423_/Y _21820_/A _21426_/Y vssd1 vssd1 vccd1 vccd1
+ _21431_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21739__B _21739_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _19016_/B vssd1 vssd1 vccd1 vccd1 _19490_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21358_ _21342_/X _21344_/X _21321_/A _21386_/B vssd1 vssd1 vccd1 vccd1 _21359_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_146_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20309_ _20309_/A _20553_/A _20553_/B _20764_/A vssd1 vssd1 vccd1 vccd1 _20311_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_151_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12091_ _11431_/A _11431_/B _11605_/A vssd1 vssd1 vccd1 vccd1 _12094_/A sky130_fd_sc_hd__a21oi_2
XFILLER_151_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21289_ _21422_/A _21289_/B vssd1 vssd1 vccd1 vccd1 _21289_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22600__A1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19072__A3 _18830_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15618__B1 _15617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__B1 _11345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15175__D _15175_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18280__A1 _11859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15850_ _15970_/A _15826_/C _15826_/A _15828_/X _15836_/X vssd1 vssd1 vccd1 vccd1
+ _15874_/B sky130_fd_sc_hd__a32o_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input20_A wb_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ _14716_/C _14800_/X _14716_/B vssd1 vssd1 vccd1 vccd1 _14802_/C sky130_fd_sc_hd__o21a_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _20249_/C _15778_/Y _15711_/A _15780_/Y vssd1 vssd1 vccd1 vccd1 _15783_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _12954_/Y _12992_/Y _12937_/Y vssd1 vssd1 vccd1 vccd1 _12993_/X sky130_fd_sc_hd__a21o_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _17520_/A _17523_/A _17520_/C _17520_/D vssd1 vssd1 vccd1 vccd1 _17520_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_18_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14732_ _14731_/B _14731_/C _14731_/A vssd1 vssd1 vccd1 vccd1 _14733_/B sky130_fd_sc_hd__a21oi_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ _12062_/A _11462_/A _11846_/Y _11774_/Y vssd1 vssd1 vccd1 vccd1 _11945_/B
+ sky130_fd_sc_hd__o22ai_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17451_ _17457_/C _17457_/D _17452_/A vssd1 vssd1 vccd1 vccd1 _17454_/A sky130_fd_sc_hd__a21o_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14663_ _14661_/C _14549_/B _14662_/Y vssd1 vssd1 vccd1 vccd1 _14664_/B sky130_fd_sc_hd__o21ai_2
X_11875_ _11922_/C _11873_/Y _11922_/B vssd1 vssd1 vccd1 vccd1 _11896_/C sky130_fd_sc_hd__o21ai_2
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16584__A _16584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output107_A _14333_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16402_ _16402_/A _16402_/B vssd1 vssd1 vccd1 vccd1 _16403_/B sky130_fd_sc_hd__nand2_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20818__B _20818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13614_ _13614_/A _13614_/B _13614_/C vssd1 vssd1 vccd1 vccd1 _13616_/B sky130_fd_sc_hd__nand3_1
X_17382_ _17380_/X _17381_/X _20928_/A _20928_/B _18197_/C vssd1 vssd1 vccd1 vccd1
+ _17382_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_38_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14594_ _14786_/C vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__buf_2
XFILLER_38_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18335__A2 _18330_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19121_ _19121_/A _19121_/B vssd1 vssd1 vccd1 vccd1 _19121_/Y sky130_fd_sc_hd__nand2_1
X_16333_ _15792_/B _16745_/A _16316_/Y _16351_/A vssd1 vssd1 vccd1 vccd1 _16333_/Y
+ sky130_fd_sc_hd__o22ai_2
X_13545_ _13550_/A _13550_/C _13501_/A vssd1 vssd1 vccd1 vccd1 _13559_/C sky130_fd_sc_hd__a21o_1
XFILLER_41_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19052_ _19052_/A _19694_/B _19346_/A vssd1 vssd1 vccd1 vccd1 _19052_/Y sky130_fd_sc_hd__nand3_1
XFILLER_186_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16264_ _16290_/A vssd1 vssd1 vccd1 vccd1 _16595_/A sky130_fd_sc_hd__clkbuf_2
X_13476_ _13215_/A _13215_/B _13443_/A vssd1 vssd1 vccd1 vccd1 _13476_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18003_ _18048_/A _18048_/B _18045_/A _18045_/B vssd1 vssd1 vccd1 vccd1 _18055_/A
+ sky130_fd_sc_hd__nand4_1
X_15215_ _15215_/A vssd1 vssd1 vccd1 vccd1 _15217_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_12427_ _12341_/A _15363_/C _12343_/B vssd1 vssd1 vccd1 vccd1 _20359_/C sky130_fd_sc_hd__a21oi_4
X_16195_ _16195_/A _16195_/B _16195_/C vssd1 vssd1 vccd1 vccd1 _16195_/Y sky130_fd_sc_hd__nand3_1
XFILLER_142_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15146_ _15146_/A vssd1 vssd1 vccd1 vccd1 _15146_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12358_ _12299_/X _12323_/Y _12346_/Y _12357_/Y vssd1 vssd1 vccd1 vccd1 _12358_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_127_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20272__C _20398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11309_ _11709_/B vssd1 vssd1 vccd1 vccd1 _11936_/C sky130_fd_sc_hd__buf_2
X_19954_ _19954_/A _19954_/B vssd1 vssd1 vccd1 vccd1 _19955_/B sky130_fd_sc_hd__or2_1
XFILLER_141_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15077_ _15128_/B _15076_/C _15076_/A vssd1 vssd1 vccd1 vccd1 _15078_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12289_ _16319_/A _12402_/A _12413_/A _12335_/A vssd1 vssd1 vccd1 vccd1 _12294_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18905_ _18905_/A _18905_/B vssd1 vssd1 vccd1 vccd1 _18905_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14028_ _14043_/A _14043_/B _14044_/C _14043_/C vssd1 vssd1 vccd1 vccd1 _14029_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19885_ _22922_/Q _19885_/B _19885_/C vssd1 vssd1 vccd1 vccd1 _19893_/A sky130_fd_sc_hd__nand3b_1
XFILLER_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12071__B _18305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16759__A _16759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18836_ _18836_/A vssd1 vssd1 vccd1 vccd1 _18836_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16821__A2 _15939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15382__B _15382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18767_ _18564_/A _18564_/B _18564_/C _18575_/B _18574_/X vssd1 vssd1 vccd1 vccd1
+ _18768_/C sky130_fd_sc_hd__a32oi_4
XFILLER_49_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15979_ _16010_/A _16010_/B _15977_/Y _15978_/X vssd1 vssd1 vccd1 vccd1 _16003_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14832__A1 _14834_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_632 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17718_ _17720_/C _17718_/B vssd1 vssd1 vccd1 vccd1 _22960_/D sky130_fd_sc_hd__xnor2_1
X_18698_ _18698_/A _18698_/B vssd1 vssd1 vccd1 vccd1 _18699_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11646__B2 _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17649_ _20928_/A _20928_/B _18303_/A _18303_/B vssd1 vssd1 vccd1 vccd1 _17649_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__22679__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_646 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20728__B _20728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16925__C _20675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20660_ _20660_/A vssd1 vssd1 vccd1 vccd1 _20660_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19319_ _12118_/A _18135_/A _19318_/Y vssd1 vssd1 vccd1 vccd1 _19319_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_17_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16337__A1 _12114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13630__B _21878_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20591_ _20704_/A _20704_/B _20591_/C vssd1 vssd1 vccd1 vccd1 _20702_/A sky130_fd_sc_hd__nand3_2
XFILLER_177_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17534__B1 _17401_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19331__A2_N _19334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22330_ _22265_/B _22304_/C _22306_/A vssd1 vssd1 vccd1 vccd1 _22330_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14348__B1 _14337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20744__A _20806_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15838__A _15838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22261_ _22304_/A _22304_/C vssd1 vssd1 vccd1 vccd1 _22308_/B sky130_fd_sc_hd__nand2_1
XFILLER_191_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21212_ _21990_/A _21351_/C _21212_/C _21990_/C vssd1 vssd1 vccd1 vccd1 _21212_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_145_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15557__B _15559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22192_ _22192_/A _22192_/B vssd1 vssd1 vccd1 vccd1 _22193_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21143_ _21143_/A _21143_/B vssd1 vssd1 vccd1 vccd1 _22924_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__15312__A2 _16178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21074_ _21074_/A _21074_/B vssd1 vssd1 vccd1 vccd1 _21124_/B sky130_fd_sc_hd__and2_1
XFILLER_116_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16669__A _16669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20025_ _20025_/A vssd1 vssd1 vccd1 vccd1 _20025_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15573__A _16937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16273__B1 _16040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15615__A3 _20098_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ _21973_/X _21854_/X _21850_/Y _22031_/B _22030_/A vssd1 vssd1 vccd1 vccd1
+ _22036_/C sky130_fd_sc_hd__o2111ai_4
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20927_ _20851_/Y _20863_/B _20863_/C _20850_/Y vssd1 vssd1 vccd1 vccd1 _20937_/A
+ sky130_fd_sc_hd__a31oi_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _11660_/A _15435_/D _16482_/A vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__nand3_1
XFILLER_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20858_ _21009_/A _17444_/A _20857_/Y vssd1 vssd1 vccd1 vccd1 _20860_/C sky130_fd_sc_hd__o21ai_2
XFILLER_30_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19211__C _19211_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11591_ _11591_/A _11591_/B _11591_/C vssd1 vssd1 vccd1 vccd1 _11592_/A sky130_fd_sc_hd__nand3_1
XFILLER_41_189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20124__A2 _15546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20789_ _20788_/B _20871_/A _20871_/B vssd1 vssd1 vccd1 vccd1 _20799_/B sky130_fd_sc_hd__a21bo_1
XFILLER_167_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13330_ _13330_/A vssd1 vssd1 vccd1 vccd1 _21990_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_195_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22528_ _13815_/X input62/X _22536_/S vssd1 vssd1 vccd1 vccd1 _22529_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ _13370_/A _13650_/B _21724_/B _21724_/C vssd1 vssd1 vccd1 vccd1 _13262_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_183_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22459_ _22459_/A vssd1 vssd1 vccd1 vccd1 _22726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ _15486_/C _12212_/B vssd1 vssd1 vccd1 vccd1 _15440_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15000_ _15001_/B _15001_/C _15001_/D _15001_/A vssd1 vssd1 vccd1 vccd1 _15018_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ _13581_/A _13192_/B _21173_/C _21173_/A vssd1 vssd1 vccd1 vccd1 _13210_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_159_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input68_A wb_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17385__D _17525_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12143_ _12143_/A _12143_/B _12143_/C vssd1 vssd1 vccd1 vccd1 _12175_/A sky130_fd_sc_hd__nand3_1
XFILLER_124_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15303__A2 _11704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16951_ _15536_/X _16240_/X _16484_/X _16483_/A _16483_/B vssd1 vssd1 vccd1 vccd1
+ _18814_/A sky130_fd_sc_hd__a32o_4
XFILLER_151_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12074_ _12074_/A _12074_/B _12074_/C _12074_/D vssd1 vssd1 vccd1 vccd1 _12074_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15483__A _22964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15902_ _16006_/B _15900_/Y _15780_/B _15901_/Y vssd1 vssd1 vccd1 vccd1 _15924_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_77_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19670_ _19670_/A _19670_/B vssd1 vssd1 vccd1 vccd1 _19880_/D sky130_fd_sc_hd__nand2_1
X_16882_ _16213_/Y _16214_/X _16378_/X _16391_/A vssd1 vssd1 vccd1 vccd1 _16882_/X
+ sky130_fd_sc_hd__o31a_1
X_18621_ _18610_/X _18611_/Y _18618_/B _17632_/A _19418_/A vssd1 vssd1 vccd1 vccd1
+ _18623_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__17461__C1 _19482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _16613_/C _17652_/B _15921_/A _15834_/A vssd1 vssd1 vccd1 vccd1 _15914_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11516__A _11583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _18553_/A _18553_/B _18553_/C vssd1 vssd1 vccd1 vccd1 _18554_/A sky130_fd_sc_hd__a21o_1
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _15683_/Y _15687_/Y _15763_/Y vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__22821__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _20134_/A vssd1 vssd1 vccd1 vccd1 _15899_/B sky130_fd_sc_hd__buf_2
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17503_ _17060_/B _17229_/Y _17352_/X _17210_/B vssd1 vssd1 vccd1 vccd1 _17503_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_166_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _14716_/A _14696_/A _14716_/C vssd1 vssd1 vccd1 vccd1 _14717_/B sky130_fd_sc_hd__a21o_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _18690_/A _18483_/B _18691_/C vssd1 vssd1 vccd1 vccd1 _18695_/A sky130_fd_sc_hd__nand3_1
X_11927_ _11927_/A _11927_/B _11927_/C vssd1 vssd1 vccd1 vccd1 _11927_/Y sky130_fd_sc_hd__nand3_1
X_15695_ _15298_/Y _15309_/A _15457_/A _19012_/C _16100_/A vssd1 vssd1 vccd1 vccd1
+ _15698_/B sky130_fd_sc_hd__o2111ai_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _17434_/A vssd1 vssd1 vccd1 vccd1 _17442_/A sky130_fd_sc_hd__buf_2
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14646_ _14646_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14646_/Y sky130_fd_sc_hd__nand2_1
X_11858_ _11306_/A _11385_/C _11273_/X _11772_/A _11420_/C vssd1 vssd1 vccd1 vccd1
+ _11859_/A sky130_fd_sc_hd__o311a_1
XANTENNA__19505__A1 _18330_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19505__B2 _11598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13450__B _21476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17365_ _17616_/C _17616_/A _17616_/B vssd1 vssd1 vccd1 vccd1 _17365_/Y sky130_fd_sc_hd__o21ai_1
X_11789_ _11789_/A vssd1 vssd1 vccd1 vccd1 _11789_/X sky130_fd_sc_hd__clkbuf_2
X_14577_ _14684_/C _14684_/A vssd1 vssd1 vccd1 vccd1 _14578_/A sky130_fd_sc_hd__nand2_1
X_19104_ _19104_/A _19254_/C _19104_/C vssd1 vssd1 vccd1 vccd1 _19104_/X sky130_fd_sc_hd__and3_1
XFILLER_192_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16316_ _15988_/A _16563_/A _16563_/B _20593_/B _16563_/C vssd1 vssd1 vccd1 vccd1
+ _16316_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13528_ _13528_/A vssd1 vssd1 vccd1 vccd1 _13528_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17296_ _17275_/Y _17285_/Y _17291_/Y _17591_/A vssd1 vssd1 vccd1 vccd1 _17304_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_9_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19035_ _19037_/A _19037_/B _19013_/X _19012_/X vssd1 vssd1 vccd1 vccd1 _19035_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_16247_ _16247_/A _16247_/B vssd1 vssd1 vccd1 vccd1 _16250_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15542__A2 _15541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13459_ _13434_/A _13436_/Y _21621_/C _13433_/C _13572_/A vssd1 vssd1 vccd1 vccd1
+ _13460_/B sky130_fd_sc_hd__o2111a_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput104 _14328_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput115 _22951_/Q vssd1 vssd1 vccd1 vccd1 y[10] sky130_fd_sc_hd__buf_2
X_16178_ _16178_/A vssd1 vssd1 vccd1 vccd1 _16179_/A sky130_fd_sc_hd__buf_2
XFILLER_126_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1098 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15129_ _15129_/A _15128_/Y vssd1 vssd1 vccd1 vccd1 _15145_/B sky130_fd_sc_hd__or2b_1
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18688__B _18691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19937_ _19937_/A _19937_/B vssd1 vssd1 vccd1 vccd1 _19955_/A sky130_fd_sc_hd__nor2_1
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16489__A _16489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15393__A _15714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19868_ _19866_/A _19866_/B _19862_/X _19863_/Y vssd1 vssd1 vccd1 vccd1 _19894_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_68_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18200__C _18453_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18819_ _18819_/A _18825_/B vssd1 vssd1 vccd1 vccd1 _18823_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19799_ _19864_/B _19799_/B vssd1 vssd1 vccd1 vccd1 _19799_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21830_ _21832_/A _21832_/B _21831_/B vssd1 vssd1 vccd1 vccd1 _21922_/B sky130_fd_sc_hd__nand3_1
XFILLER_37_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21761_ _21761_/A _21761_/B vssd1 vssd1 vccd1 vccd1 _21762_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17113__A _19619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20712_ _20702_/A _20702_/B _20702_/C _20702_/D vssd1 vssd1 vccd1 vccd1 _20712_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_169_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21692_ _21809_/A _21814_/A _21809_/B vssd1 vssd1 vccd1 vccd1 _21693_/C sky130_fd_sc_hd__nand3_1
XFILLER_180_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20643_ _20568_/B _20567_/Y _20568_/A vssd1 vssd1 vccd1 vccd1 _20645_/B sky130_fd_sc_hd__o21ai_1
XFILLER_177_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12257__A _22909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20574_ _20734_/B _20637_/A _20728_/A _20449_/B vssd1 vssd1 vccd1 vccd1 _20574_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_164_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22313_ _22313_/A _22313_/B vssd1 vssd1 vccd1 vccd1 _22314_/C sky130_fd_sc_hd__and2_1
XFILLER_11_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15533__A2 _15524_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22244_ _22244_/A _22244_/B vssd1 vssd1 vccd1 vccd1 _22244_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17286__A2 _11563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22175_ _22229_/B vssd1 vssd1 vccd1 vccd1 _22265_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21126_ _21150_/A _21127_/B _21127_/C vssd1 vssd1 vccd1 vccd1 _21128_/A sky130_fd_sc_hd__a21oi_1
XFILLER_87_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13847__A2 _14013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__B1 _11306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13816__A _22867_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21057_ _21095_/C vssd1 vssd1 vccd1 vccd1 _21057_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22844__CLK _22937_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12720__A _20255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20008_ _20008_/A _20008_/B _22925_/Q vssd1 vssd1 vccd1 vccd1 _20010_/A sky130_fd_sc_hd__nor3b_1
XFILLER_189_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18110__C _18367_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12830_ _15362_/D _15370_/A vssd1 vssd1 vccd1 vccd1 _20213_/A sky130_fd_sc_hd__nand2_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18538__A2 _18371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _20415_/A vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ _22108_/C vssd1 vssd1 vccd1 vccd1 _22182_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14500_/A _14500_/B _14500_/C vssd1 vssd1 vccd1 vccd1 _14607_/B sky130_fd_sc_hd__nand3_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11712_/A _11712_/B _11712_/C _15482_/C vssd1 vssd1 vccd1 vccd1 _11718_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _15502_/A _15502_/B _15501_/A _15502_/D vssd1 vssd1 vccd1 vccd1 _15597_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _20471_/C vssd1 vssd1 vccd1 vccd1 _20584_/C sky130_fd_sc_hd__clkbuf_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14431_/A vssd1 vssd1 vccd1 vccd1 _14432_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11698_/A _11698_/B _11698_/C vssd1 vssd1 vccd1 vccd1 _11643_/Y sky130_fd_sc_hd__nand3_2
XFILLER_187_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15772__A2 _15646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17150_ _16952_/X _17136_/X _17146_/Y _17149_/Y vssd1 vssd1 vccd1 vccd1 _17168_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_11_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13783__A1 _14079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11574_ _19619_/B _18629_/A _11565_/B _11565_/A vssd1 vssd1 vccd1 vccd1 _11899_/B
+ sky130_fd_sc_hd__a22o_2
X_14362_ _22763_/Q vssd1 vssd1 vccd1 vccd1 _14362_/X sky130_fd_sc_hd__buf_2
XFILLER_156_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18171__B1 _19504_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput17 wb_adr_i[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16101_ _12716_/X _11912_/A _11541_/X _15890_/A vssd1 vssd1 vccd1 vccd1 _16103_/C
+ sky130_fd_sc_hd__o22ai_2
Xinput28 wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_1
X_13313_ _13316_/A _21202_/A _13324_/B _13300_/Y vssd1 vssd1 vccd1 vccd1 _13314_/C
+ sky130_fd_sc_hd__o211ai_1
Xinput39 wb_dat_i[13] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17081_ _17081_/A _17591_/B vssd1 vssd1 vccd1 vccd1 _17081_/Y sky130_fd_sc_hd__nor2_2
X_14293_ _14553_/B _14553_/A vssd1 vssd1 vccd1 vccd1 _14843_/A sky130_fd_sc_hd__xnor2_4
XFILLER_196_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16032_ _15966_/X _15921_/X _16024_/Y _16200_/C vssd1 vssd1 vccd1 vccd1 _16038_/B
+ sky130_fd_sc_hd__o31a_2
X_13244_ _22722_/Q vssd1 vssd1 vccd1 vccd1 _13257_/B sky130_fd_sc_hd__buf_2
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17277__A2 _15808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ _13465_/A _13169_/X _13465_/B vssd1 vssd1 vccd1 vccd1 _13221_/A sky130_fd_sc_hd__a21boi_1
XFILLER_123_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12120__A1_N _18208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12126_ _12126_/A vssd1 vssd1 vccd1 vccd1 _12126_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17983_ _21017_/A _21017_/B _19945_/B _17039_/C _19454_/C vssd1 vssd1 vccd1 vccd1
+ _18030_/D sky130_fd_sc_hd__a32o_1
XFILLER_111_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19722_ _19611_/X _19613_/Y _19631_/Y _19724_/A vssd1 vssd1 vccd1 vccd1 _19723_/B
+ sky130_fd_sc_hd__o31a_1
X_16934_ _16934_/A vssd1 vssd1 vccd1 vccd1 _16934_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12057_ _12054_/X _12056_/Y _12039_/Y _12081_/A vssd1 vssd1 vccd1 vccd1 _12245_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__19423__B1 _19211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12630__A _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A3 _11404_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19653_ _19740_/A _19656_/B _19652_/Y vssd1 vssd1 vccd1 vccd1 _19653_/Y sky130_fd_sc_hd__a21boi_1
X_16865_ _16866_/A _16866_/B _16863_/Y _16864_/X vssd1 vssd1 vccd1 vccd1 _16867_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16788__A1 _15530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16788__B2 _12294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18604_ _18268_/A _18268_/B _18434_/A vssd1 vssd1 vccd1 vccd1 _18604_/Y sky130_fd_sc_hd__o21ai_1
X_15816_ _15825_/B _15825_/C vssd1 vssd1 vccd1 vccd1 _15817_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15941__A _15941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19584_ _19350_/X _17400_/X _17647_/A _11639_/X vssd1 vssd1 vccd1 vccd1 _19602_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_19_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16796_ _16796_/A _16796_/B _16796_/C vssd1 vssd1 vccd1 vccd1 _16834_/A sky130_fd_sc_hd__nand3_1
XFILLER_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18535_ _18664_/B _18533_/Y _18534_/X vssd1 vssd1 vccd1 vccd1 _18535_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _15516_/Y _15517_/Y _15746_/Y vssd1 vssd1 vccd1 vccd1 _15747_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12959_ _13004_/B _12959_/B vssd1 vssd1 vccd1 vccd1 _12960_/B sky130_fd_sc_hd__nor2_1
XANTENNA__18029__A _21086_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18466_ _18451_/A _18451_/B _19046_/C _17525_/D _18450_/B vssd1 vssd1 vccd1 vccd1
+ _18466_/Y sky130_fd_sc_hd__o2111ai_4
X_15678_ _15678_/A _15678_/B _15678_/C _15678_/D vssd1 vssd1 vccd1 vccd1 _15680_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_763 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17417_ _17298_/A _17298_/C _17377_/Y vssd1 vssd1 vccd1 vccd1 _17420_/A sky130_fd_sc_hd__a21o_1
XFILLER_53_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14629_ _14917_/C _14629_/B _14911_/A _15010_/C vssd1 vssd1 vccd1 vccd1 _14629_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_159_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18397_ _18408_/C _18397_/B vssd1 vssd1 vccd1 vccd1 _18397_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16772__A _16772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17348_ _17330_/Y _17337_/X _17339_/X vssd1 vssd1 vccd1 vccd1 _17350_/B sky130_fd_sc_hd__a21o_1
XFILLER_158_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17279_ _17293_/A vssd1 vssd1 vccd1 vccd1 _17449_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19018_ _19014_/X _19015_/Y _19017_/Y vssd1 vssd1 vccd1 vccd1 _19026_/A sky130_fd_sc_hd__o21ai_1
XFILLER_161_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20290_ _20290_/A _20290_/B _20290_/C vssd1 vssd1 vccd1 vccd1 _20294_/B sky130_fd_sc_hd__nand3_1
XFILLER_161_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18465__A1 _19043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22867__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15835__B _16613_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18849__D _18849_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18217__A1 _18208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17108__A _19012_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21221__B1 _13350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21853__A _21853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22931_ _22933_/CLK _22931_/D vssd1 vssd1 vccd1 vccd1 _22931_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16947__A _16947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18865__C _19602_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22862_ _22933_/CLK _22874_/Q vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfxtp_2
XFILLER_83_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16666__B _16670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19717__A1 _16015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19178__C1 _19334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14254__A2 _15154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21813_ _21805_/X _21677_/A _21797_/Y _21804_/A vssd1 vssd1 vccd1 vccd1 _21913_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_58_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19042__B _19504_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22793_ _22795_/CLK _22793_/D vssd1 vssd1 vccd1 vccd1 _22793_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19193__A2 _19694_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21744_ _21383_/X _21958_/A _21743_/Y vssd1 vssd1 vccd1 vccd1 _21761_/A sky130_fd_sc_hd__o21ai_1
XFILLER_58_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13214__B1 _13350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21675_ _21664_/X _21674_/Y _21671_/Y vssd1 vssd1 vccd1 vccd1 _21676_/C sky130_fd_sc_hd__a21o_1
XFILLER_178_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13765__A1 _14892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20626_ _20626_/A vssd1 vssd1 vccd1 vccd1 _20630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22834__D _22846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17928__D _17928_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20557_ _20566_/A _20566_/B _22933_/Q vssd1 vssd1 vccd1 vccd1 _20559_/A sky130_fd_sc_hd__o21ai_1
XFILLER_192_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18105__C _19317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ _22955_/Q vssd1 vssd1 vccd1 vccd1 _11325_/A sky130_fd_sc_hd__inv_2
X_20488_ _12721_/X _15939_/A _12832_/Y _20481_/Y _20482_/Y vssd1 vssd1 vccd1 vccd1
+ _20488_/X sky130_fd_sc_hd__o221a_1
XFILLER_106_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22227_ _22186_/X _22225_/Y _22222_/X _22224_/Y vssd1 vssd1 vccd1 vccd1 _22263_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_156_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22158_ _21698_/B _21698_/C _21838_/B vssd1 vssd1 vccd1 vccd1 _22158_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20370__C _20608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21109_ _16585_/A _16585_/B _20843_/X vssd1 vssd1 vccd1 vccd1 _21109_/X sky130_fd_sc_hd__a21o_1
X_22089_ _22089_/A vssd1 vssd1 vccd1 vccd1 _22284_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14980_ _14980_/A _15035_/B _14980_/C vssd1 vssd1 vccd1 vccd1 _15039_/A sky130_fd_sc_hd__and3_1
XFILLER_102_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16219__B1 _18192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13931_ _14765_/A _14506_/B _14765_/C _14117_/A _14107_/A vssd1 vssd1 vccd1 vccd1
+ _13931_/X sky130_fd_sc_hd__a32o_2
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16650_ _16895_/A _16895_/B _16650_/C vssd1 vssd1 vccd1 vccd1 _16653_/B sky130_fd_sc_hd__nand3_1
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13862_ _13862_/A _14061_/A _14061_/D vssd1 vssd1 vccd1 vccd1 _13862_/X sky130_fd_sc_hd__and3_1
XFILLER_47_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15601_ _15474_/C _15474_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15601_/Y sky130_fd_sc_hd__a21oi_2
X_12813_ _12813_/A vssd1 vssd1 vccd1 vccd1 _16450_/C sky130_fd_sc_hd__buf_2
X_16581_ _16435_/B _16579_/X _16580_/X _22702_/Q vssd1 vssd1 vccd1 vccd1 _16582_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_90_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13793_ _13810_/A _13963_/B _13810_/B vssd1 vssd1 vccd1 vccd1 _13793_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__15993__A2 _15905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19184__A2 _19162_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18320_ _18512_/B _18512_/C vssd1 vssd1 vccd1 vccd1 _19011_/A sky130_fd_sc_hd__nor2_1
X_15532_ _15530_/X _15531_/X _12571_/A _12571_/B vssd1 vssd1 vccd1 vccd1 _15532_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14808__C _14808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12744_ _12739_/A _12739_/B _12739_/C _13002_/C vssd1 vssd1 vccd1 vccd1 _12744_/Y
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__13712__C _15115_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18251_ _18251_/A _18251_/B _18251_/C vssd1 vssd1 vccd1 vccd1 _18251_/Y sky130_fd_sc_hd__nand3_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15755_/A _15439_/X _15448_/X _15517_/A _15517_/B vssd1 vssd1 vccd1 vccd1
+ _15756_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_124_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12675_/A vssd1 vssd1 vccd1 vccd1 _12749_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17202_ _17197_/Y _17201_/Y _17198_/X vssd1 vssd1 vccd1 vccd1 _17205_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14414_ _22809_/Q _14411_/X _14412_/X _14413_/X _22777_/Q vssd1 vssd1 vccd1 vccd1
+ _14414_/X sky130_fd_sc_hd__a32o_1
XFILLER_156_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18182_ _18182_/A vssd1 vssd1 vccd1 vccd1 _18277_/A sky130_fd_sc_hd__clkbuf_2
X_11626_ _11394_/A _11378_/X _11306_/X vssd1 vssd1 vccd1 vccd1 _11626_/X sky130_fd_sc_hd__o21a_4
X_15394_ _15394_/A vssd1 vssd1 vccd1 vccd1 _15909_/A sky130_fd_sc_hd__buf_2
XFILLER_11_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17133_ _17133_/A _17631_/A vssd1 vssd1 vccd1 vccd1 _17133_/Y sky130_fd_sc_hd__nand2_2
X_14345_ _18115_/A _14338_/X _14339_/X _14334_/X _13736_/C vssd1 vssd1 vccd1 vccd1
+ _14345_/X sky130_fd_sc_hd__a32o_1
X_11557_ _22959_/Q vssd1 vssd1 vccd1 vccd1 _15435_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__12625__A _16486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17064_ _17215_/D _17064_/B _17064_/C vssd1 vssd1 vccd1 vccd1 _17222_/B sky130_fd_sc_hd__nand3b_1
XFILLER_128_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14276_ _14279_/C _14276_/B _14276_/C _14276_/D vssd1 vssd1 vccd1 vccd1 _14277_/C
+ sky130_fd_sc_hd__and4b_1
X_11488_ _11608_/A _11608_/B _11980_/C vssd1 vssd1 vccd1 vccd1 _12158_/A sky130_fd_sc_hd__nand3_1
XFILLER_6_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16015_ _16015_/A vssd1 vssd1 vccd1 vccd1 _16015_/X sky130_fd_sc_hd__buf_4
XANTENNA__18447__A1 _11634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15936__A _15936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13227_ _13396_/A _13396_/B _13396_/C vssd1 vssd1 vccd1 vccd1 _13484_/A sky130_fd_sc_hd__nand3_1
XFILLER_170_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18312__A _22796_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20254__A1 _20241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16458__B1 _15997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18998__A2 _18678_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13158_ _13158_/A vssd1 vssd1 vccd1 vccd1 _13161_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _15714_/B _18510_/A _12094_/A _12001_/Y _12004_/B vssd1 vssd1 vccd1 vccd1
+ _12110_/C sky130_fd_sc_hd__a32oi_4
XFILLER_2_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17966_ _17967_/C _17967_/A _22904_/Q vssd1 vssd1 vccd1 vccd1 _17968_/A sky130_fd_sc_hd__a21oi_1
X_13089_ _13050_/X _21341_/A _13139_/A vssd1 vssd1 vccd1 vccd1 _13122_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__15374__C _15912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18966__B _22914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14484__A2 _13746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19705_ _19705_/A _19705_/B vssd1 vssd1 vccd1 vccd1 _19708_/B sky130_fd_sc_hd__nor2_1
X_16917_ _15580_/X _17443_/A _16926_/A vssd1 vssd1 vccd1 vccd1 _16919_/B sky130_fd_sc_hd__o21ai_1
XFILLER_78_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17897_ _17897_/A _17897_/B _17897_/C vssd1 vssd1 vccd1 vccd1 _17899_/A sky130_fd_sc_hd__nand3_1
X_19636_ _19636_/A _19636_/B vssd1 vssd1 vccd1 vccd1 _19636_/X sky130_fd_sc_hd__and2_1
X_16848_ _16853_/A vssd1 vssd1 vccd1 vccd1 _16848_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22919__D _22919_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16486__B _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19567_ _19681_/A _19681_/C _19681_/B vssd1 vssd1 vccd1 vccd1 _19569_/A sky130_fd_sc_hd__nand3_4
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16779_ _16779_/A vssd1 vssd1 vccd1 vccd1 _16779_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13444__B1 _13475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15984__A2 _12716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18518_ _18518_/A vssd1 vssd1 vccd1 vccd1 _18916_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19498_ _19365_/X _19489_/X _19492_/Y _19497_/Y vssd1 vssd1 vccd1 vccd1 _19511_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__16918__D1 _19619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12519__B _12519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18449_ _18795_/A _15839_/A _18448_/Y vssd1 vssd1 vccd1 vccd1 _18450_/B sky130_fd_sc_hd__o21ai_2
XFILLER_179_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16933__A1 _16059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21460_ _21460_/A _21460_/B _21460_/C _21460_/D vssd1 vssd1 vccd1 vccd1 _21651_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_159_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18206__B _18571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20411_ _20395_/A _20395_/B _20396_/A vssd1 vssd1 vccd1 vccd1 _20411_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17110__B _17110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21391_ _21247_/A _21247_/B _21380_/Y vssd1 vssd1 vccd1 vccd1 _21404_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12535__A _22824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20493__A1 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20342_ _20342_/A vssd1 vssd1 vccd1 vccd1 _20464_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__20493__B2 _12967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19318__A _19318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20273_ _20397_/A _20397_/B _20398_/A vssd1 vssd1 vccd1 vccd1 _20273_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12183__B1 _12123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20471__B _20471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22012_ _21915_/Y _21932_/Y _22011_/X vssd1 vssd1 vccd1 vccd1 _22014_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12722__A2 _12718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12270__A _22703_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18876__B _18876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_546 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18595__C _22912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22914_ _22915_/CLK _22914_/D vssd1 vssd1 vccd1 vccd1 _22914_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__18610__B2 _15531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22829__D _22841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21733__D _22106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12238__A1 _12234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22845_ _22943_/CLK hold17/X vssd1 vssd1 vccd1 vccd1 _22845_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__18892__A _19587_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22776_ _22808_/CLK _22776_/D vssd1 vssd1 vccd1 vccd1 _22776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21727_ _21724_/Y _21455_/X _21733_/A _21638_/B _21726_/Y vssd1 vssd1 vccd1 vccd1
+ _21730_/C sky130_fd_sc_hd__o2111ai_4
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21658_ _21658_/A _21658_/B _21658_/C vssd1 vssd1 vccd1 vccd1 _21658_/X sky130_fd_sc_hd__and3_1
X_12460_ _16477_/C _17144_/A _20694_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _12460_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11411_ _11411_/A vssd1 vssd1 vccd1 vccd1 _16482_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12410__A1 _15631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12391_ _17141_/A _12683_/A vssd1 vssd1 vccd1 vccd1 _12391_/Y sky130_fd_sc_hd__nand2_1
X_20609_ _16267_/X _16266_/X _20241_/A _16268_/X vssd1 vssd1 vccd1 vccd1 _20609_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21589_ _21596_/A _21596_/B vssd1 vssd1 vccd1 vccd1 _21589_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12445__A _15394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14950__A3 _14013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14130_ _13829_/A _14123_/X _13873_/X _14085_/Y _14727_/A vssd1 vssd1 vccd1 vccd1
+ _14237_/B sky130_fd_sc_hd__o2111ai_2
X_11342_ _11764_/B vssd1 vssd1 vccd1 vccd1 _12148_/B sky130_fd_sc_hd__buf_2
XFILLER_4_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16152__A2 _15905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14061_ _14061_/A _14491_/C _14512_/A _14061_/D vssd1 vssd1 vccd1 vccd1 _14061_/X
+ sky130_fd_sc_hd__and4_1
X_11273_ _11374_/A vssd1 vssd1 vccd1 vccd1 _11273_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19626__B1 _19476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_75 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input50_A wb_dat_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13910__A1 _13904_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13012_ _13012_/A _13012_/B vssd1 vssd1 vccd1 vccd1 _13012_/Y sky130_fd_sc_hd__nand2_1
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17101__B2 _16727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17820_ _17731_/A _19839_/C _17927_/A _15941_/X vssd1 vssd1 vccd1 vccd1 _17821_/C
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19929__A1 _19293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17751_ _19772_/D vssd1 vssd1 vccd1 vccd1 _19844_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_130_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_14963_ _14963_/A _14963_/B _14963_/C vssd1 vssd1 vccd1 vccd1 _14969_/A sky130_fd_sc_hd__and3_1
XANTENNA__12477__A1 _12500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16702_ _16702_/A _16702_/B vssd1 vssd1 vccd1 vccd1 _16702_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17404__A2 _20255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13914_ _13923_/A vssd1 vssd1 vccd1 vccd1 _14618_/A sky130_fd_sc_hd__clkbuf_2
X_17682_ _17687_/C _17687_/A _17687_/B vssd1 vssd1 vccd1 vccd1 _17682_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14894_ _14895_/A _14895_/B _14895_/C vssd1 vssd1 vccd1 vccd1 _14966_/A sky130_fd_sc_hd__a21o_1
X_19421_ _19304_/Y _19305_/Y _19417_/Y _19420_/Y vssd1 vssd1 vccd1 vccd1 _19428_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16612__B1 _15645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16633_ _16630_/A _16630_/B _16637_/B _16637_/A vssd1 vssd1 vccd1 vccd1 _16634_/C
+ sky130_fd_sc_hd__o211ai_1
X_13845_ _13849_/B _13845_/B _13896_/A vssd1 vssd1 vccd1 vccd1 _13985_/B sky130_fd_sc_hd__nand3_1
XFILLER_74_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19352_ _19352_/A vssd1 vssd1 vccd1 vccd1 _19352_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13977__A1 _22858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16564_ _16563_/Y _16564_/B _16996_/A vssd1 vssd1 vccd1 vccd1 _16586_/A sky130_fd_sc_hd__nand3b_2
X_13776_ _13776_/A _13776_/B _14699_/B vssd1 vssd1 vccd1 vccd1 _14184_/B sky130_fd_sc_hd__nand3_2
XFILLER_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18303_ _18303_/A _18303_/B _18303_/C vssd1 vssd1 vccd1 vccd1 _18459_/A sky130_fd_sc_hd__and3_2
XFILLER_188_543 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15515_ _15385_/A _15512_/Y _15514_/X vssd1 vssd1 vccd1 vccd1 _15859_/B sky130_fd_sc_hd__a21o_1
X_19283_ _19134_/A _19134_/B _19138_/Y vssd1 vssd1 vccd1 vccd1 _19681_/C sky130_fd_sc_hd__a21oi_2
X_12727_ _12727_/A vssd1 vssd1 vccd1 vccd1 _15890_/A sky130_fd_sc_hd__buf_2
X_16495_ _16506_/A _16762_/A _16496_/A _16100_/D _19507_/B vssd1 vssd1 vccd1 vccd1
+ _16512_/A sky130_fd_sc_hd__o2111ai_4
XANTENNA__16915__A1 _16275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18234_ _18232_/X _18233_/Y _18224_/Y _18230_/Y vssd1 vssd1 vccd1 vccd1 _18234_/X
+ sky130_fd_sc_hd__o211a_1
X_15446_ _15528_/A vssd1 vssd1 vccd1 vccd1 _19047_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_176_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12658_ _12742_/A _12640_/B _12640_/A vssd1 vssd1 vccd1 vccd1 _12757_/B sky130_fd_sc_hd__a21boi_2
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14554__B _14554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18668__A1 _11979_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18165_ _18165_/A _18165_/B vssd1 vssd1 vccd1 vccd1 _18173_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11609_ _22791_/Q vssd1 vssd1 vccd1 vccd1 _11616_/C sky130_fd_sc_hd__inv_2
XFILLER_156_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18668__B2 _11639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15377_ _15377_/A vssd1 vssd1 vccd1 vccd1 _15918_/A sky130_fd_sc_hd__buf_2
XFILLER_11_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14941__A3 _15004_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12589_ _20346_/C vssd1 vssd1 vccd1 vccd1 _20471_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_144_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17116_ _17116_/A _17116_/B vssd1 vssd1 vccd1 vccd1 _17120_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14273__C _14273_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14328_ _12470_/X _14308_/X _14313_/X _13257_/B _14327_/X vssd1 vssd1 vccd1 vccd1
+ _14328_/X sky130_fd_sc_hd__a221o_1
X_18096_ _12018_/A _16276_/A _18091_/Y vssd1 vssd1 vccd1 vccd1 _18096_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_128_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20572__A _20575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17047_ _17229_/A vssd1 vssd1 vccd1 vccd1 _17603_/B sky130_fd_sc_hd__buf_2
XANTENNA__15351__B1 _15350_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14259_ _14259_/A _14259_/B vssd1 vssd1 vccd1 vccd1 _14259_/X sky130_fd_sc_hd__or2_1
XFILLER_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20227__A1 _12697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17881__A _19585_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18840__A1 _19504_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ _18698_/B _18678_/D _15427_/X vssd1 vssd1 vccd1 vccd1 _19000_/C sky130_fd_sc_hd__a21oi_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17949_ _17949_/A _17949_/B vssd1 vssd1 vccd1 vccd1 _17950_/B sky130_fd_sc_hd__or2_1
XFILLER_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20960_ _20832_/Y _20902_/Y _20773_/B _20903_/Y vssd1 vssd1 vccd1 vccd1 _20960_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19619_ _19792_/A _19619_/B _19900_/A _19619_/D vssd1 vssd1 vccd1 vccd1 _19621_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_398 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20891_ _20891_/A _20891_/B vssd1 vssd1 vccd1 vccd1 _20892_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21850__B _22108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22630_ _22803_/Q input45/X _22630_/S vssd1 vssd1 vccd1 vccd1 _22631_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11979__B1 _11980_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22561_ _22772_/Q input47/X _22569_/S vssd1 vssd1 vccd1 vccd1 _22562_/A sky130_fd_sc_hd__mux2_1
XANTENNA__19320__B _19490_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21512_ _21508_/Y _21485_/X _21650_/C _21650_/B vssd1 vssd1 vccd1 vccd1 _21512_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_179_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22492_ _22492_/A vssd1 vssd1 vccd1 vccd1 _22741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21443_ _21522_/D vssd1 vssd1 vccd1 vccd1 _22172_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21374_ _21374_/A _21374_/B vssd1 vssd1 vccd1 vccd1 _21374_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15576__A _16912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20325_ _20508_/A _15909_/A _20323_/Y _20324_/Y vssd1 vssd1 vccd1 vccd1 _20328_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14911__C _14911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20256_ _20255_/X _20109_/Y _20098_/Y vssd1 vssd1 vccd1 vccd1 _20262_/A sky130_fd_sc_hd__o21ai_4
XFILLER_131_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20187_ _12754_/X _12894_/Y _13045_/Y _20186_/Y vssd1 vssd1 vccd1 vccd1 _20189_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_62_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _11751_/X _11703_/X _11935_/X _12219_/A _12220_/A vssd1 vssd1 vccd1 vccd1
+ _12054_/A sky130_fd_sc_hd__o2111ai_4
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22391__A1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_622 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15948__A2 _15942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _18629_/A vssd1 vssd1 vccd1 vccd1 _18305_/B sky130_fd_sc_hd__buf_2
XANTENNA__11682__A2 _15297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ _13630_/A _21878_/C _13664_/A _13635_/A vssd1 vssd1 vccd1 vccd1 _13630_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11419__C1 _11430_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22828_ _22933_/CLK hold7/X vssd1 vssd1 vccd1 vccd1 _22828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13561_ _13677_/A _13677_/B _13677_/C vssd1 vssd1 vccd1 vccd1 _13611_/B sky130_fd_sc_hd__a21bo_1
XFILLER_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22759_ _22762_/CLK _22759_/D vssd1 vssd1 vccd1 vccd1 _22759_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15300_ _18107_/B _18107_/C _15901_/C vssd1 vssd1 vccd1 vccd1 _15302_/A sky130_fd_sc_hd__nand3_2
X_12512_ _12520_/A _12518_/A _12324_/X vssd1 vssd1 vccd1 vccd1 _12513_/A sky130_fd_sc_hd__o21ai_1
XFILLER_157_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16280_ _16595_/B _16596_/A _16595_/A vssd1 vssd1 vccd1 vccd1 _16283_/B sky130_fd_sc_hd__nand3b_2
XFILLER_160_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13492_ _13492_/A _13492_/B vssd1 vssd1 vccd1 vccd1 _13493_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17570__A1 _17442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15231_ _15231_/A _15231_/B vssd1 vssd1 vccd1 vccd1 _15233_/A sky130_fd_sc_hd__xor2_4
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12443_ _15466_/B vssd1 vssd1 vccd1 vccd1 _15799_/A sky130_fd_sc_hd__buf_2
XFILLER_173_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15581__B1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19311__A2 _19308_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15162_ _15163_/A _15163_/B _15163_/C vssd1 vssd1 vccd1 vccd1 _15162_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_165_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12374_ _12374_/A _12374_/B vssd1 vssd1 vccd1 vccd1 _12487_/B sky130_fd_sc_hd__nand2_1
XFILLER_193_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14113_ _14963_/A _14113_/B _14963_/B _14191_/C vssd1 vssd1 vccd1 vccd1 _14113_/X
+ sky130_fd_sc_hd__and4_1
X_11325_ _11325_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11325_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15333__B1 _17532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19970_ _19970_/A _22923_/Q _19970_/C vssd1 vssd1 vccd1 vccd1 _19976_/B sky130_fd_sc_hd__nand3_1
XFILLER_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15093_ _15093_/A vssd1 vssd1 vccd1 vccd1 _15095_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12903__A _20133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20209__A1 _20210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18921_ _18839_/X _18865_/X _18912_/A _18870_/Y _18853_/A vssd1 vssd1 vccd1 vccd1
+ _18921_/X sky130_fd_sc_hd__o311a_1
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14044_ _14044_/A _14044_/B _14044_/C vssd1 vssd1 vccd1 vccd1 _14044_/Y sky130_fd_sc_hd__nand3_2
XFILLER_141_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12698__A1 _12696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18797__A _19351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17086__B1 _17085_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11519__A _11968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18852_ _18862_/A _18854_/A _18861_/A _18861_/B vssd1 vssd1 vccd1 vccd1 _18853_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_79_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15636__A1 _15319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17803_ _17760_/A _17760_/B _17760_/C _17765_/A vssd1 vssd1 vccd1 vccd1 _17900_/B
+ sky130_fd_sc_hd__a31o_1
X_18783_ _18783_/A _18958_/A vssd1 vssd1 vccd1 vccd1 _19138_/D sky130_fd_sc_hd__nand2_1
X_15995_ _16047_/C _16047_/D vssd1 vssd1 vccd1 vccd1 _15995_/Y sky130_fd_sc_hd__nand2_1
X_17734_ _17873_/A _17928_/A _17928_/D _17876_/A vssd1 vssd1 vccd1 vccd1 _17734_/X
+ sky130_fd_sc_hd__o22a_1
X_14946_ _14947_/A _14947_/B _14947_/C _14947_/D vssd1 vssd1 vccd1 vccd1 _14959_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17389__A1 _15941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17665_ _17665_/A _17665_/B _17665_/C vssd1 vssd1 vccd1 vccd1 _17687_/C sky130_fd_sc_hd__nand3_1
XANTENNA__11673__A2 _11666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14877_ _14880_/A _14880_/B _14877_/C vssd1 vssd1 vccd1 vccd1 _14887_/B sky130_fd_sc_hd__nand3_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19404_ _19248_/A _19248_/B _19403_/Y _19106_/B vssd1 vssd1 vccd1 vccd1 _19404_/Y
+ sky130_fd_sc_hd__a22oi_1
X_16616_ _16873_/A _16617_/C _16615_/Y _16310_/Y vssd1 vssd1 vccd1 vccd1 _16624_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__16061__B2 _16177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13828_ _13959_/A _13828_/B vssd1 vssd1 vccd1 vccd1 _13829_/B sky130_fd_sc_hd__nand2_1
XFILLER_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17596_ _17597_/B _17597_/C _17597_/A vssd1 vssd1 vccd1 vccd1 _17600_/B sky130_fd_sc_hd__a21oi_1
XFILLER_91_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19335_ _19587_/B vssd1 vssd1 vccd1 vccd1 _19768_/B sky130_fd_sc_hd__buf_2
X_16547_ _16541_/X _16546_/Y _16534_/B _16536_/B vssd1 vssd1 vccd1 vccd1 _16548_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__21244__A1_N _13339_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ _22753_/Q _13707_/B _13733_/B vssd1 vssd1 vccd1 vccd1 _13766_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11404__D _11404_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19266_ _19043_/X _19899_/B _19265_/X _19065_/X vssd1 vssd1 vccd1 vccd1 _19272_/C
+ sky130_fd_sc_hd__o31ai_2
XANTENNA__20696__B2 _20792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16478_ _15455_/A _16786_/A _16782_/A vssd1 vssd1 vccd1 vccd1 _16479_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__16364__A2 _16627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17561__A1 _16579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18217_ _18208_/A _18208_/B _18216_/B vssd1 vssd1 vccd1 vccd1 _18417_/B sky130_fd_sc_hd__a21oi_1
X_15429_ _15427_/X _15933_/A _15331_/Y _15329_/X _15344_/X vssd1 vssd1 vccd1 vccd1
+ _15430_/C sky130_fd_sc_hd__o221ai_2
XANTENNA__14375__A1 _22798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19197_ _19197_/A _19496_/B _19197_/C _19197_/D vssd1 vssd1 vccd1 vccd1 _19215_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_129_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14375__B2 _22766_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_1_bq_clk_i clkbuf_1_0_1_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__16780__A _18445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12386__B1 _12387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18148_ _12126_/X _12128_/X _12131_/Y _12134_/B vssd1 vssd1 vccd1 vccd1 _18389_/A
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_144_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15396__A _19329_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18079_ _18079_/A _18079_/B vssd1 vssd1 vccd1 vccd1 _22967_/D sky130_fd_sc_hd__xor2_1
XFILLER_171_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20110_ _20110_/A _20110_/B vssd1 vssd1 vccd1 vccd1 _20110_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18203__C _18203_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19066__A1 _11308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21090_ _21090_/A _21090_/B _21090_/C vssd1 vssd1 vccd1 vccd1 _21091_/B sky130_fd_sc_hd__and3_1
XFILLER_125_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20041_ _20041_/A _20041_/B vssd1 vssd1 vccd1 vccd1 _20042_/C sky130_fd_sc_hd__xnor2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21992_ _21987_/Y _21989_/Y _22075_/B vssd1 vssd1 vccd1 vccd1 _22029_/B sky130_fd_sc_hd__o21ai_2
XFILLER_66_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20384__B1 _20337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20943_ _20877_/A _20877_/B _20945_/A _20945_/B _20876_/B vssd1 vssd1 vccd1 vccd1
+ _20949_/B sky130_fd_sc_hd__a221oi_2
XFILLER_27_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20874_ _20787_/B _20787_/C _20706_/X vssd1 vssd1 vccd1 vccd1 _20874_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22613_ _18128_/C input37/X _22619_/S vssd1 vssd1 vccd1 vccd1 _22614_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22544_ _22544_/A vssd1 vssd1 vccd1 vccd1 _22764_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__19985__B _20012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12707__B _16489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22475_ _22734_/Q input40/X _22475_/S vssd1 vssd1 vccd1 vccd1 _22476_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21426_ _21426_/A _21426_/B _21426_/C vssd1 vssd1 vccd1 vccd1 _21426_/Y sky130_fd_sc_hd__nand3_1
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21357_ _21321_/A _21333_/A _21509_/A _21509_/B vssd1 vssd1 vccd1 vccd1 _21359_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_146_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12129__B1 _11771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20308_ _20314_/B vssd1 vssd1 vccd1 vccd1 _20764_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12090_ _12090_/A _12090_/B _12090_/C vssd1 vssd1 vccd1 vccd1 _12090_/X sky130_fd_sc_hd__or3_1
X_21288_ _21422_/A _21559_/A _21424_/C vssd1 vssd1 vccd1 vccd1 _21288_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_146_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17068__B1 _22895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20239_ _20237_/X _20238_/Y _20118_/B _20119_/B vssd1 vssd1 vccd1 vccd1 _20240_/C
+ sky130_fd_sc_hd__a22oi_4
XFILLER_118_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15618__A1 _15904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16815__B1 _17131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15618__B2 _12827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18280__A2 _11861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _14681_/X _14682_/X _14687_/X _14689_/Y vssd1 vssd1 vccd1 vccd1 _14800_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _15780_/A _15780_/B vssd1 vssd1 vccd1 vccd1 _15780_/Y sky130_fd_sc_hd__nor2_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12992_ _12705_/X _12737_/D _12942_/Y _12943_/X vssd1 vssd1 vccd1 vccd1 _12992_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_A wb_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ _14731_/A _14731_/B _14731_/C vssd1 vssd1 vccd1 vccd1 _14733_/A sky130_fd_sc_hd__and3_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _11943_/A _11943_/B vssd1 vssd1 vccd1 vccd1 _11947_/A sky130_fd_sc_hd__nand2_1
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_806 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17450_ _17457_/A _17523_/C vssd1 vssd1 vccd1 vccd1 _17452_/A sky130_fd_sc_hd__nand2_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14553_/A _14553_/B _14661_/Y vssd1 vssd1 vccd1 vccd1 _14662_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11874_ _11874_/A _12074_/A _12074_/B vssd1 vssd1 vccd1 vccd1 _11922_/B sky130_fd_sc_hd__nand3_1
XFILLER_189_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _16397_/X _16400_/X _16429_/A _16431_/C vssd1 vssd1 vccd1 vccd1 _16433_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13613_ _13552_/A _13512_/B _13614_/B _13614_/A vssd1 vssd1 vccd1 vccd1 _13616_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_17381_ _17381_/A vssd1 vssd1 vccd1 vccd1 _17381_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14593_ _14863_/B _14593_/B _22764_/Q vssd1 vssd1 vccd1 vccd1 _14786_/C sky130_fd_sc_hd__nand3_1
XFILLER_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19120_ _19303_/B _19117_/X _19118_/X _18927_/Y _19119_/X vssd1 vssd1 vccd1 vccd1
+ _19121_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_111_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16332_ _16332_/A _16332_/B vssd1 vssd1 vccd1 vccd1 _16351_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_1074 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13544_ _13614_/C _13614_/B _13548_/A vssd1 vssd1 vccd1 vccd1 _13559_/B sky130_fd_sc_hd__a21bo_1
XFILLER_186_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_855 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19051_ _12157_/X _12158_/X _15530_/X _15531_/X vssd1 vssd1 vccd1 vccd1 _19051_/X
+ sky130_fd_sc_hd__a22o_2
XANTENNA__14357__A1 _16322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16263_ _16265_/A _16265_/B _16263_/C _16263_/D vssd1 vssd1 vccd1 vccd1 _16290_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11521__B _18875_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13475_ _13475_/A _13475_/B _13475_/C vssd1 vssd1 vccd1 vccd1 _13475_/Y sky130_fd_sc_hd__nand3_1
X_18002_ _18002_/A _18044_/A _18002_/C vssd1 vssd1 vccd1 vccd1 _18045_/B sky130_fd_sc_hd__nand3_1
XFILLER_127_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15214_ _15238_/A _15240_/C _15216_/A vssd1 vssd1 vccd1 vccd1 _15214_/X sky130_fd_sc_hd__o21a_1
XANTENNA__21627__B1 _21853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12426_ _12403_/A _15631_/B _15631_/C _12377_/A vssd1 vssd1 vccd1 vccd1 _20359_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16194_ _16145_/A _16145_/C _16146_/Y vssd1 vssd1 vccd1 vccd1 _16195_/C sky130_fd_sc_hd__a21oi_1
XFILLER_138_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21011__A _21011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15145_ _15145_/A _15145_/B vssd1 vssd1 vccd1 vccd1 _15145_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12357_ _12334_/X _12350_/Y _12734_/A _15409_/A vssd1 vssd1 vccd1 vccd1 _12357_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_154_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11308_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11709_/B sky130_fd_sc_hd__nand2_1
X_19953_ _19991_/A _19952_/B _19991_/B vssd1 vssd1 vccd1 vccd1 _19954_/B sky130_fd_sc_hd__a21oi_1
X_15076_ _15076_/A _15128_/B _15076_/C vssd1 vssd1 vccd1 vccd1 _15078_/A sky130_fd_sc_hd__nand3_1
XFILLER_142_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12288_ _12288_/A vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__buf_2
X_18904_ _18705_/A _18705_/B _18707_/A _18707_/B vssd1 vssd1 vccd1 vccd1 _18904_/Y
+ sky130_fd_sc_hd__a22oi_1
X_14027_ _14043_/A _14043_/B _14044_/C _14043_/C vssd1 vssd1 vccd1 vccd1 _14029_/A
+ sky130_fd_sc_hd__nand4_1
X_19884_ _19885_/B _19885_/C _22922_/Q vssd1 vssd1 vccd1 vccd1 _19976_/A sky130_fd_sc_hd__a21bo_1
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18320__A _18512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16759__B _17139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12071__C _16192_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18835_ _18835_/A _18933_/B _18835_/C _19112_/A vssd1 vssd1 vccd1 vccd1 _18929_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18766_ _18757_/X _18758_/Y _18754_/X _18765_/X vssd1 vssd1 vccd1 vccd1 _18768_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15382__C _16062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15978_ _15978_/A _15978_/B _15978_/C _17645_/D vssd1 vssd1 vccd1 vccd1 _15978_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_49_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14832__A2 _14834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17717_ _17608_/X _17610_/Y _17619_/B _17722_/A vssd1 vssd1 vccd1 vccd1 _17718_/B
+ sky130_fd_sc_hd__a22o_1
X_14929_ _14929_/A _14929_/B _14929_/C _14845_/A vssd1 vssd1 vccd1 vccd1 _15046_/A
+ sky130_fd_sc_hd__or4b_2
X_18697_ _11770_/X _18500_/Y _18841_/B _18678_/D vssd1 vssd1 vccd1 vccd1 _18699_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18574__A3 _18572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22927__D _22927_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17648_ _17645_/D _19689_/C _17817_/A _15919_/X vssd1 vssd1 vccd1 vccd1 _17648_/Y
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_1_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14596__A1 _13748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17579_ _17524_/Y _17579_/B _17579_/C vssd1 vssd1 vccd1 vccd1 _17579_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_51_658 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14295__A input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19318_ _19318_/A _19322_/B _19322_/C vssd1 vssd1 vccd1 vccd1 _19318_/Y sky130_fd_sc_hd__nand3_2
X_20590_ _20464_/B _20697_/B _20695_/A _20579_/X vssd1 vssd1 vccd1 vccd1 _20591_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16337__A2 _16179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14348__A1 _12343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19249_ _19082_/Y _19089_/A _19033_/X _19039_/Y vssd1 vssd1 vccd1 vccd1 _19249_/Y
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22260_ _22306_/B _21970_/X _22233_/B _22232_/B vssd1 vssd1 vccd1 vccd1 _22301_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21211_ _21211_/A vssd1 vssd1 vccd1 vccd1 _21238_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__20463__C _20463_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22191_ _22190_/D _22190_/A _22190_/B _22219_/B vssd1 vssd1 vccd1 vccd1 _22192_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__19692__D1 _18197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15557__C _15558_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21142_ _21142_/A _21150_/C vssd1 vssd1 vccd1 vccd1 _21143_/B sky130_fd_sc_hd__or2b_1
XFILLER_105_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22043__B1 _21963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19326__A _19326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21073_ _21065_/X _21071_/Y _21072_/Y vssd1 vssd1 vccd1 vccd1 _21074_/B sky130_fd_sc_hd__o21ai_1
XFILLER_132_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21397__A2 _21445_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20024_ _20024_/A _20024_/B _20024_/C vssd1 vssd1 vccd1 vccd1 _20029_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13874__A3 _13736_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input5_A wb_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16273__A1 _16016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16273__B2 _15580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21975_ _22031_/B _22030_/A _22030_/B vssd1 vssd1 vccd1 vccd1 _22036_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16685__A _16685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18801__A1_N _12170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19061__A _19061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20926_ _20925_/Y _20936_/B _20936_/C _20936_/D vssd1 vssd1 vccd1 vccd1 _20926_/X
+ sky130_fd_sc_hd__and4b_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12047__C1 _11721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ _20782_/B _20854_/Y _20855_/Y vssd1 vssd1 vccd1 vccd1 _20857_/Y sky130_fd_sc_hd__o21ai_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11590_ _11528_/Y _11793_/A _18797_/C _15988_/A _11589_/X vssd1 vssd1 vccd1 vccd1
+ _11591_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20124__A3 _20123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20788_ _20871_/B _20788_/B _20871_/A vssd1 vssd1 vccd1 vccd1 _20799_/A sky130_fd_sc_hd__nand3b_1
XFILLER_70_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11341__B _22786_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22527_ _22584_/S vssd1 vssd1 vccd1 vccd1 _22536_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_195_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ _21367_/C vssd1 vssd1 vccd1 vccd1 _21724_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22458_ _13055_/A input63/X _22464_/S vssd1 vssd1 vccd1 vccd1 _22459_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12211_ _12211_/A vssd1 vssd1 vccd1 vccd1 _17381_/A sky130_fd_sc_hd__clkbuf_4
X_21409_ _21547_/B _21401_/B _21403_/Y _21404_/Y _21390_/Y vssd1 vssd1 vccd1 vccd1
+ _21410_/C sky130_fd_sc_hd__o221ai_2
XFILLER_68_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13191_ _13450_/A vssd1 vssd1 vccd1 vccd1 _21173_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22389_ _12343_/B input65/X _22391_/S vssd1 vssd1 vccd1 vccd1 _22390_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12142_ _12126_/X _12128_/X _12131_/Y _18510_/A _15357_/A vssd1 vssd1 vccd1 vccd1
+ _12143_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_135_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15186__D _15186_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18778__C _19983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14511__A1 _15008_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16950_ _16225_/X _16227_/X _17144_/C vssd1 vssd1 vccd1 vccd1 _17403_/A sky130_fd_sc_hd__o21ai_2
X_12073_ _17039_/D _19046_/C vssd1 vssd1 vccd1 vccd1 _12074_/D sky130_fd_sc_hd__xnor2_1
XFILLER_173_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_75 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15901_ _15901_/A _15901_/B _15901_/C vssd1 vssd1 vccd1 vccd1 _15901_/Y sky130_fd_sc_hd__nand3_4
X_16881_ _17042_/A _16885_/B _16879_/X _16880_/X vssd1 vssd1 vccd1 vccd1 _17049_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15832_ _17385_/B vssd1 vssd1 vccd1 vccd1 _17652_/B sky130_fd_sc_hd__clkbuf_4
X_18620_ _12064_/A _17526_/X _18616_/A vssd1 vssd1 vccd1 vccd1 _18623_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__17461__B1 _20972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _15514_/X _15512_/Y _15682_/Y vssd1 vssd1 vccd1 vccd1 _15763_/Y sky130_fd_sc_hd__a21oi_1
X_18551_ _18360_/X _18367_/A _18544_/X vssd1 vssd1 vccd1 vccd1 _18553_/C sky130_fd_sc_hd__a21oi_2
XFILLER_66_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12989_/A _13024_/B _16106_/A _12975_/D vssd1 vssd1 vccd1 vccd1 _12989_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _17502_/A vssd1 vssd1 vccd1 vccd1 _17502_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14714_ _14714_/A _14714_/B _14714_/C vssd1 vssd1 vccd1 vccd1 _14737_/A sky130_fd_sc_hd__nand3_2
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _18482_/A _18482_/B _19165_/A _19168_/C vssd1 vssd1 vccd1 vccd1 _18482_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11926_ _11693_/X _11565_/Y _12059_/B _12247_/B vssd1 vssd1 vccd1 vccd1 _11927_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_166_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15694_ _15694_/A vssd1 vssd1 vccd1 vccd1 _19012_/C sky130_fd_sc_hd__clkbuf_4
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16567__A2 _16324_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17430_/Y _17433_/B _17433_/C vssd1 vssd1 vccd1 vccd1 _17523_/B sky130_fd_sc_hd__nand3b_4
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _22863_/D vssd1 vssd1 vccd1 vccd1 _14963_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _19418_/A _16564_/B _11399_/Y _11393_/Y vssd1 vssd1 vccd1 vccd1 _12074_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19505__A2 _17400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11532__A _18706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17364_ _22897_/Q vssd1 vssd1 vccd1 vccd1 _17616_/B sky130_fd_sc_hd__inv_2
XFILLER_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14576_ _14576_/A vssd1 vssd1 vccd1 vccd1 _14576_/X sky130_fd_sc_hd__buf_2
X_11788_ _11595_/X _11589_/X _11583_/Y vssd1 vssd1 vccd1 vccd1 _11799_/A sky130_fd_sc_hd__a21boi_2
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19103_ _19104_/A _19254_/C _19104_/C vssd1 vssd1 vccd1 vccd1 _19103_/Y sky130_fd_sc_hd__a21oi_1
X_16315_ _16311_/X _16314_/Y _16309_/Y _16301_/Y vssd1 vssd1 vccd1 vccd1 _16315_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15939__A _15939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13527_ _13563_/A _13563_/B _13563_/C vssd1 vssd1 vccd1 vccd1 _13527_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_186_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17295_ _17464_/B _17464_/A _17292_/X _17294_/X vssd1 vssd1 vccd1 vccd1 _17591_/A
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_174_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14843__A _14843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19034_ _18899_/B _18899_/C _18899_/A vssd1 vssd1 vccd1 vccd1 _19034_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_174_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16246_ _19197_/C _19197_/D _16515_/A vssd1 vssd1 vccd1 vccd1 _16247_/B sky130_fd_sc_hd__and3_1
XFILLER_12_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _13572_/A _21621_/C _13457_/Y _13433_/C vssd1 vssd1 vccd1 vccd1 _13460_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_103_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12409_ _12409_/A vssd1 vssd1 vccd1 vccd1 _15325_/A sky130_fd_sc_hd__clkbuf_4
X_16177_ _16177_/A vssd1 vssd1 vccd1 vccd1 _20449_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput105 _14426_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[30] sky130_fd_sc_hd__buf_2
X_13389_ _13339_/Y _13353_/Y _13359_/A vssd1 vssd1 vccd1 vccd1 _13391_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12363__A _12378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput116 _22952_/Q vssd1 vssd1 vccd1 vccd1 y[11] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_891 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15128_ _15128_/A _15128_/B _15128_/C _15128_/D vssd1 vssd1 vccd1 vccd1 _15128_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_5_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19936_ _19894_/A _19921_/A _19922_/B vssd1 vssd1 vccd1 vccd1 _19962_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__18688__C _18690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15059_ _14503_/X _15057_/A _15005_/Y vssd1 vssd1 vccd1 vccd1 _15059_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_68_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16489__B _16770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21233__D1 _21805_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19441__A1 _19293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19867_ _19862_/X _19863_/Y _19866_/X vssd1 vssd1 vccd1 vccd1 _19867_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18985__A _19480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__A _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18818_ _18818_/A _18818_/B vssd1 vssd1 vccd1 vccd1 _18825_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19798_ _19725_/C _19860_/A _19798_/C vssd1 vssd1 vccd1 vccd1 _19866_/A sky130_fd_sc_hd__nand3b_2
XFILLER_110_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18749_ _18608_/Y _18609_/Y _18738_/Y _18748_/Y vssd1 vssd1 vccd1 vccd1 _18763_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_110_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21760_ _21760_/A _21760_/B vssd1 vssd1 vccd1 vccd1 _21762_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20711_ _20709_/B _20709_/C _20709_/A vssd1 vssd1 vccd1 vccd1 _20711_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_196_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21691_ _21809_/A _21814_/A _21809_/B vssd1 vssd1 vccd1 vccd1 _21693_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12538__A _22824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20642_ _20631_/Y _20737_/A _20574_/X _20575_/X vssd1 vssd1 vccd1 vccd1 _20645_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_149_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18704__B1 _11800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15781__A3 _15711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20573_ _20449_/A _20728_/B _20519_/C _20512_/Y _20519_/B vssd1 vssd1 vccd1 vccd1
+ _20637_/A sky130_fd_sc_hd__o221ai_4
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_622 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22312_ _22304_/B _22263_/B _22263_/C _22302_/Y _22310_/X vssd1 vssd1 vccd1 vccd1
+ _22313_/B sky130_fd_sc_hd__a311o_1
XFILLER_30_1111 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_666 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22243_ _22243_/A _22243_/B vssd1 vssd1 vccd1 vccd1 _22244_/B sky130_fd_sc_hd__and2_1
XFILLER_180_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22174_ _22231_/D _22173_/B _22173_/D _22173_/A vssd1 vssd1 vccd1 vccd1 _22176_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_87_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11960__D1 _12220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21125_ _22942_/Q _21122_/X _21130_/B _21130_/A vssd1 vssd1 vccd1 vccd1 _21127_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_120_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21056_ _21061_/B _21061_/A vssd1 vssd1 vccd1 vccd1 _21095_/C sky130_fd_sc_hd__xor2_1
XFILLER_115_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20007_ _20008_/A _20008_/B _22925_/Q vssd1 vssd1 vccd1 vccd1 _20057_/B sky130_fd_sc_hd__o21bai_1
XFILLER_115_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18110__D _18848_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12760_ _22826_/Q vssd1 vssd1 vccd1 vccd1 _20415_/A sky130_fd_sc_hd__inv_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21958_ _21958_/A vssd1 vssd1 vccd1 vccd1 _21958_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _22959_/Q _22960_/Q vssd1 vssd1 vccd1 vccd1 _15482_/C sky130_fd_sc_hd__nor2_2
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _20892_/A _20908_/Y _20894_/B vssd1 vssd1 vccd1 vccd1 _20950_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__20750__B1 _20751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12691_ _12749_/A _13007_/A vssd1 vssd1 vccd1 vccd1 _12920_/C sky130_fd_sc_hd__xor2_1
XFILLER_14_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21889_ _21889_/A _21889_/B _21889_/C vssd1 vssd1 vccd1 vccd1 _21896_/A sky130_fd_sc_hd__nand3_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12448__A _15394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14430_/A vssd1 vssd1 vccd1 vccd1 _14431_/A sky130_fd_sc_hd__buf_4
XANTENNA__13768__C1 _13761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11635_/X _11641_/X _11647_/A _11647_/B vssd1 vssd1 vccd1 vccd1 _11698_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_74_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _14361_/A vssd1 vssd1 vccd1 vccd1 _14361_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13783__A2 _14489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11573_ _11664_/D vssd1 vssd1 vccd1 vccd1 _18629_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__18135__A _18135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16100_ _16100_/A _19000_/A _16106_/C _16100_/D vssd1 vssd1 vccd1 vccd1 _16150_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_7_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 wb_adr_i[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input80_A x[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13312_ _21213_/A _21480_/B _21214_/A vssd1 vssd1 vccd1 vccd1 _13324_/B sky130_fd_sc_hd__and3_1
X_17080_ _16580_/X _16579_/X _16711_/C _17462_/A vssd1 vssd1 vccd1 vccd1 _17591_/B
+ sky130_fd_sc_hd__o211ai_4
Xinput29 wb_adr_i[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_1
X_14292_ _14180_/Y _14289_/Y _14290_/X _14291_/Y vssd1 vssd1 vccd1 vccd1 _14553_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_10_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_0_0_bq_clk_i_A clkbuf_2_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16031_ _16043_/A _16043_/B _16028_/Y _16030_/Y vssd1 vssd1 vccd1 vccd1 _16200_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__15909__D _15988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13243_ _13243_/A vssd1 vssd1 vccd1 vccd1 _21584_/C sky130_fd_sc_hd__buf_4
XFILLER_136_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13174_ _13170_/Y _13172_/Y _13173_/Y vssd1 vssd1 vccd1 vccd1 _13465_/B sky130_fd_sc_hd__o21ai_2
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16485__A1 _14429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ _12006_/Y _11986_/X _11972_/Y _11976_/Y vssd1 vssd1 vccd1 vccd1 _12177_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__22669__CLK _22964_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17982_ _19842_/D vssd1 vssd1 vccd1 vccd1 _19945_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_151_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19721_ _19725_/B _19725_/C vssd1 vssd1 vccd1 vccd1 _19723_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19423__A1 _12064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16933_ _16059_/A _17634_/A _16932_/Y vssd1 vssd1 vccd1 vccd1 _16934_/A sky130_fd_sc_hd__o21ai_4
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ _12088_/B _12055_/Y _11930_/X _11933_/Y vssd1 vssd1 vccd1 vccd1 _12056_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19652_ _19652_/A _19652_/B vssd1 vssd1 vccd1 vccd1 _19652_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16864_ _16753_/A _16753_/B _16733_/Y _16740_/Y _16848_/X vssd1 vssd1 vccd1 vccd1
+ _16864_/X sky130_fd_sc_hd__o221a_1
XANTENNA__16788__A2 _15531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18603_ _19443_/A _18599_/X _18602_/Y vssd1 vssd1 vccd1 vccd1 _18603_/Y sky130_fd_sc_hd__o21bai_1
X_15815_ _15714_/X _15814_/Y _15752_/B _15752_/C vssd1 vssd1 vccd1 vccd1 _15825_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_19_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19583_ _19689_/A _19687_/B _19687_/C _19836_/C vssd1 vssd1 vccd1 vccd1 _19602_/A
+ sky130_fd_sc_hd__nand4_1
X_16795_ _16508_/X _16510_/Y _16493_/Y _16517_/Y vssd1 vssd1 vccd1 vccd1 _16796_/C
+ sky130_fd_sc_hd__o22ai_1
XFILLER_93_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15746_ _15748_/A _15746_/B _19772_/D _15748_/B vssd1 vssd1 vccd1 vccd1 _15746_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_34_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18534_ _11431_/A _11431_/B _17421_/X _17422_/X vssd1 vssd1 vccd1 vccd1 _18534_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12958_ _12958_/A _12958_/B _12958_/C vssd1 vssd1 vccd1 vccd1 _12959_/B sky130_fd_sc_hd__and3_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11909_ _11909_/A _11909_/B _11909_/C vssd1 vssd1 vccd1 vccd1 _12077_/C sky130_fd_sc_hd__nand3_1
X_18465_ _19043_/A _17730_/A _18451_/Y _18452_/X vssd1 vssd1 vccd1 vccd1 _18465_/X
+ sky130_fd_sc_hd__o22a_1
X_15677_ _15677_/A _15677_/B _15677_/C vssd1 vssd1 vccd1 vccd1 _15680_/A sky130_fd_sc_hd__nand3_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _12889_/A _12889_/B _12889_/C vssd1 vssd1 vccd1 vccd1 _13043_/B sky130_fd_sc_hd__nand3_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17416_ _17416_/A _17416_/B _17416_/C vssd1 vssd1 vccd1 vccd1 _17457_/C sky130_fd_sc_hd__nand3_1
X_14628_ _15008_/C vssd1 vssd1 vccd1 vccd1 _15061_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18396_ _18396_/A _18396_/B _18396_/C _18559_/A vssd1 vssd1 vccd1 vccd1 _18396_/Y
+ sky130_fd_sc_hd__nand4_2
XANTENNA__20575__A _20734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21297__A1 _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17347_ _17346_/Y _17350_/A _17206_/B vssd1 vssd1 vccd1 vccd1 _17347_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_14_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14559_ _22875_/Q vssd1 vssd1 vccd1 vccd1 _14560_/A sky130_fd_sc_hd__inv_2
XFILLER_174_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17278_ _16275_/A _16708_/X _17277_/Y vssd1 vssd1 vccd1 vccd1 _17293_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__21049__A1 _21017_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16229_ _14429_/A _16241_/C _16228_/Y _11714_/A vssd1 vssd1 vccd1 vccd1 _17251_/A
+ sky130_fd_sc_hd__o211ai_4
X_19017_ _11702_/X _19176_/A _19016_/Y vssd1 vssd1 vccd1 vccd1 _19017_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_174_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15920__B1 _15918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1070 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18465__A2 _17730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15835__C _17652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19919_ _19919_/A _19919_/B vssd1 vssd1 vccd1 vccd1 _19919_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16228__A1 _16482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11437__A _22957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17425__B1 _17423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22930_ _22933_/CLK _22930_/D vssd1 vssd1 vccd1 vccd1 _22930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16947__B _17139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22861_ _22915_/CLK _22873_/Q vssd1 vssd1 vccd1 vccd1 _22861_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19178__B1 _18849_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19717__A2 _19838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21812_ _21797_/Y _21913_/A _21806_/X vssd1 vssd1 vccd1 vccd1 _21814_/B sky130_fd_sc_hd__a21o_1
XFILLER_97_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19042__C _19504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22792_ _22795_/CLK _22792_/D vssd1 vssd1 vccd1 vccd1 _22792_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21743_ _21610_/B _21740_/X _21742_/Y vssd1 vssd1 vccd1 vccd1 _21743_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_58_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19977__C _22924_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21674_ _21650_/X _21653_/Y _21673_/Y _21656_/Y vssd1 vssd1 vccd1 vccd1 _21674_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_178_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13765__A2 _14079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20625_ _20501_/X _20623_/Y _20624_/X vssd1 vssd1 vccd1 vccd1 _20631_/B sky130_fd_sc_hd__a21o_1
XFILLER_193_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20556_ _20548_/X _20551_/Y _20554_/Y _20764_/A vssd1 vssd1 vccd1 vccd1 _20566_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_153_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18105__D _18367_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20487_ _20479_/Y _20476_/Y _20486_/X vssd1 vssd1 vccd1 vccd1 _20487_/X sky130_fd_sc_hd__o21a_1
XFILLER_152_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22226_ _22186_/A _22186_/B _22222_/X _22224_/Y _22225_/Y vssd1 vssd1 vccd1 vccd1
+ _22228_/A sky130_fd_sc_hd__o221a_1
XANTENNA__22850__D hold22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16467__A1 _16269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22157_ _22212_/A _22212_/B vssd1 vssd1 vccd1 vccd1 _22157_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21108_ _21097_/A _21095_/Y _21094_/Y vssd1 vssd1 vccd1 vccd1 _21108_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_191_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22961__CLK _22964_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22088_ _22145_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _22088_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16219__A1 _12500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14493__A3 _14963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13930_ _13930_/A _13930_/B vssd1 vssd1 vccd1 vccd1 _14117_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21039_ _21039_/A _21039_/B _22940_/Q vssd1 vssd1 vccd1 vccd1 _21076_/D sky130_fd_sc_hd__nand3_1
XFILLER_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13861_ _14061_/A _14061_/D _13862_/A vssd1 vssd1 vccd1 vccd1 _13861_/Y sky130_fd_sc_hd__a21oi_1
X_15600_ _15678_/A _15678_/B vssd1 vssd1 vccd1 vccd1 _15677_/A sky130_fd_sc_hd__nand2_1
X_12812_ _12428_/Y _12334_/X _12350_/Y vssd1 vssd1 vccd1 vccd1 _12818_/A sky130_fd_sc_hd__a21boi_1
XFILLER_90_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16580_ _16580_/A vssd1 vssd1 vccd1 vccd1 _16580_/X sky130_fd_sc_hd__clkbuf_4
X_13792_ _14273_/A _15082_/A vssd1 vssd1 vccd1 vccd1 _14049_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15531_ _15531_/A vssd1 vssd1 vccd1 vccd1 _15531_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_12_0_bq_clk_i clkbuf_3_6_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _22948_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _13007_/D _13007_/A vssd1 vssd1 vccd1 vccd1 _13002_/C sky130_fd_sc_hd__xor2_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13712__D _14273_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _18772_/B _18250_/B vssd1 vssd1 vccd1 vccd1 _18251_/C sky130_fd_sc_hd__nand2_1
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _15449_/X _15502_/B _15457_/Y _15461_/Y vssd1 vssd1 vccd1 vccd1 _15517_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_31_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12674_ _12742_/A _12742_/B vssd1 vssd1 vccd1 vccd1 _12675_/A sky130_fd_sc_hd__or2_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17187_/X _17191_/Y _17200_/Y _17192_/X vssd1 vssd1 vccd1 vccd1 _17201_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14413_/A vssd1 vssd1 vccd1 vccd1 _14413_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15489__A _15489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18181_ _18181_/A _18181_/B _18181_/C vssd1 vssd1 vccd1 vccd1 _18182_/A sky130_fd_sc_hd__nand3_1
X_11625_ _11450_/A _11395_/A _18674_/A _11299_/X vssd1 vssd1 vccd1 vccd1 _11625_/X
+ sky130_fd_sc_hd__o211a_4
X_15393_ _15714_/A vssd1 vssd1 vccd1 vccd1 _19329_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_8_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12906__A _15901_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19341__B1 _19512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17132_ _17128_/Y _17134_/A _17131_/Y vssd1 vssd1 vccd1 vccd1 _17270_/A sky130_fd_sc_hd__a21o_1
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14344_ _14370_/A vssd1 vssd1 vccd1 vccd1 _14344_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11556_ _11712_/A _11659_/B _11712_/C vssd1 vssd1 vccd1 vccd1 _11668_/A sky130_fd_sc_hd__nand3_4
XFILLER_10_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17063_ _17226_/A _17227_/A _17371_/A vssd1 vssd1 vccd1 vccd1 _17064_/B sky130_fd_sc_hd__o21ai_1
XFILLER_183_474 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14275_ _14998_/A _14272_/C _14203_/X _14185_/X _14206_/Y vssd1 vssd1 vccd1 vccd1
+ _14276_/C sky130_fd_sc_hd__o221a_1
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21938__B _21938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11487_ _18115_/D vssd1 vssd1 vccd1 vccd1 _11980_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_170_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16014_ _16014_/A vssd1 vssd1 vccd1 vccd1 _16015_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13226_ _13223_/Y _13225_/X _13340_/A _13286_/B vssd1 vssd1 vccd1 vccd1 _13396_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__18447__A2 _17635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16458__A1 _18445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16458__B2 _16471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21451__A1 _21853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20254__A2 _15450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ _13157_/A vssd1 vssd1 vccd1 vccd1 _21336_/C sky130_fd_sc_hd__buf_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12108_ _12108_/A _12108_/B vssd1 vssd1 vccd1 vccd1 _18510_/A sky130_fd_sc_hd__nand2_2
XFILLER_111_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _17961_/Y _17962_/Y _17963_/X _17964_/Y vssd1 vssd1 vccd1 vccd1 _17967_/A
+ sky130_fd_sc_hd__o22ai_2
X_13088_ _13120_/B _13316_/A _13300_/A _13105_/A vssd1 vssd1 vccd1 vccd1 _13139_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15374__D _17281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12360__B _12687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19704_ _19705_/A _19705_/B _19789_/A _19708_/A vssd1 vssd1 vccd1 vccd1 _19704_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__21203__A1 _13305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22400__A0 _14369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16916_ _16911_/X _16913_/X _16915_/Y vssd1 vssd1 vccd1 vccd1 _16926_/A sky130_fd_sc_hd__o21ai_1
X_12039_ _12039_/A _12039_/B _12039_/C vssd1 vssd1 vccd1 vccd1 _12039_/Y sky130_fd_sc_hd__nand3_2
X_17896_ _17896_/A _17896_/B vssd1 vssd1 vccd1 vccd1 _17897_/C sky130_fd_sc_hd__nand2_1
XFILLER_19_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19635_ _19635_/A _19724_/B vssd1 vssd1 vccd1 vccd1 _19635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16847_ _16847_/A _16866_/B _16866_/A vssd1 vssd1 vccd1 vccd1 _16860_/B sky130_fd_sc_hd__nand3_1
XFILLER_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16486__C _16486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19566_ _19561_/A _19561_/B _19565_/Y vssd1 vssd1 vccd1 vccd1 _19669_/B sky130_fd_sc_hd__a21o_1
XFILLER_18_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16778_ _16778_/A vssd1 vssd1 vccd1 vccd1 _16778_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12101__D1 _18453_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14641__B1 _14512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18517_ _18526_/A _18526_/B vssd1 vssd1 vccd1 vccd1 _18518_/A sky130_fd_sc_hd__nand2_1
X_15729_ _15713_/A _15728_/X _15714_/X vssd1 vssd1 vccd1 vccd1 _15733_/A sky130_fd_sc_hd__a21oi_2
XFILLER_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13995__A2 _14686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19497_ _19497_/A _19497_/B vssd1 vssd1 vccd1 vccd1 _19497_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16918__C1 _17525_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12519__C _12669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18448_ _17381_/X _17380_/X _18107_/A _18200_/A vssd1 vssd1 vccd1 vccd1 _18448_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16933__A2 _17634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15399__A _16257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18379_ _18389_/A _18389_/B _18389_/C _18310_/Y _18383_/A vssd1 vssd1 vccd1 vccd1
+ _18381_/B sky130_fd_sc_hd__a32oi_1
XFILLER_193_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22834__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18206__C _18571_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20410_ _20378_/Y _20381_/Y _20396_/B _20388_/Y vssd1 vssd1 vccd1 vccd1 _20410_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_175_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21390_ _21535_/A _21535_/B _21535_/C vssd1 vssd1 vccd1 vccd1 _21390_/Y sky130_fd_sc_hd__nand3_2
XFILLER_179_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21690__A1 _22167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20341_ _20341_/A _20341_/B _20341_/C vssd1 vssd1 vccd1 vccd1 _20342_/A sky130_fd_sc_hd__nand3_1
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21848__B _21848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20272_ _20397_/A _20397_/B _20398_/A vssd1 vssd1 vccd1 vccd1 _20272_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__19318__B _19322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12183__A1 _18208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20245__A2 _16932_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22011_ _22008_/A _22007_/A _21908_/C _21911_/A vssd1 vssd1 vccd1 vccd1 _22011_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__20471__C _20471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17119__A _19012_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16958__A _20129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19334__A _19334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18876__C _18876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_992 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13085__C _21476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22913_ _22916_/CLK _22913_/D vssd1 vssd1 vccd1 vccd1 _22913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22844_ _22937_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 _22844_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12238__A2 _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11614__B _18665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22775_ _22807_/CLK _22775_/D vssd1 vssd1 vccd1 vccd1 _22775_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21726_ _13423_/A _21183_/X _21725_/Y vssd1 vssd1 vccd1 vccd1 _21726_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22458__A0 _13055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21657_ _21650_/X _21653_/Y _21656_/Y vssd1 vssd1 vccd1 vccd1 _21657_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11410_ _11712_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _11436_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11630__A _11647_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20608_ _20608_/A _20608_/B _20608_/C _20917_/A vssd1 vssd1 vccd1 vccd1 _20608_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_137_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12390_ _22822_/Q vssd1 vssd1 vccd1 vccd1 _12683_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21588_ _21936_/A _21588_/B _21588_/C vssd1 vssd1 vccd1 vccd1 _21596_/B sky130_fd_sc_hd__nand3_2
XANTENNA__12445__B _15799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11341_ _22787_/Q _22786_/Q vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20539_ _20658_/A vssd1 vssd1 vccd1 vccd1 _20539_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ _14117_/A vssd1 vssd1 vccd1 vccd1 _14512_/A sky130_fd_sc_hd__buf_2
XANTENNA__19626__A1 _16015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11272_ _22785_/Q vssd1 vssd1 vccd1 vccd1 _11374_/A sky130_fd_sc_hd__buf_2
XFILLER_180_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13371__B1 _21584_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ _13011_/A _13011_/B _13011_/C _13011_/D vssd1 vssd1 vccd1 vccd1 _13045_/A
+ sky130_fd_sc_hd__nand4_4
XANTENNA__17637__B1 _17732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22209_ _22290_/D vssd1 vssd1 vccd1 vccd1 _22209_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15648__C1 _16400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A wb_dat_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19929__A2 _19294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__D _20576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17750_ _17752_/B _17752_/C _15840_/X _17981_/D vssd1 vssd1 vccd1 vccd1 _17753_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__21493__B _21725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14962_ _14930_/A _14930_/B _14961_/B vssd1 vssd1 vccd1 vccd1 _14971_/A sky130_fd_sc_hd__a21o_1
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12477__A2 _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16701_ _16889_/B _16673_/A _16665_/X _17065_/A vssd1 vssd1 vccd1 vccd1 _16702_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13913_ _14069_/C _14069_/A vssd1 vssd1 vccd1 vccd1 _13924_/A sky130_fd_sc_hd__nand2_4
XFILLER_75_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17681_ _17681_/A _17681_/B vssd1 vssd1 vccd1 vccd1 _17687_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17404__A3 _17647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14893_ _14893_/A _14955_/B vssd1 vssd1 vccd1 vccd1 _14895_/C sky130_fd_sc_hd__nand2_1
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16612__A1 _11541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19420_ _19411_/X _19555_/A _19418_/X _19419_/X vssd1 vssd1 vccd1 vccd1 _19420_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16632_ _16391_/B _16636_/B _16636_/A vssd1 vssd1 vccd1 vccd1 _16634_/B sky130_fd_sc_hd__a21o_1
X_13844_ _22760_/Q vssd1 vssd1 vccd1 vccd1 _13896_/A sky130_fd_sc_hd__buf_2
XFILLER_74_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19351_ _19351_/A _19351_/B _19351_/C vssd1 vssd1 vccd1 vccd1 _19352_/A sky130_fd_sc_hd__nand3_2
XFILLER_74_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16563_ _16563_/A _16563_/B _16563_/C vssd1 vssd1 vccd1 vccd1 _16563_/Y sky130_fd_sc_hd__nand3_1
X_13775_ _13845_/B vssd1 vssd1 vccd1 vccd1 _14699_/B sky130_fd_sc_hd__buf_2
XANTENNA__13977__A2 _14911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18302_ _18309_/B vssd1 vssd1 vccd1 vccd1 _18571_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__22857__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15514_ _15397_/Y _15513_/Y _15700_/C _15707_/B vssd1 vssd1 vccd1 vccd1 _15514_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12726_ _12583_/A _12630_/A _12721_/X _12716_/X vssd1 vssd1 vccd1 vccd1 _12916_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_19282_ _19284_/A _19284_/B _19282_/C _19750_/A vssd1 vssd1 vccd1 vccd1 _19286_/A
+ sky130_fd_sc_hd__nand4_1
X_16494_ _16494_/A vssd1 vssd1 vccd1 vccd1 _16494_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16915__A2 _15919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15445_ _15445_/A _15445_/B vssd1 vssd1 vccd1 vccd1 _15528_/A sky130_fd_sc_hd__nand2_2
X_18233_ _18275_/A _18275_/B vssd1 vssd1 vccd1 vccd1 _18233_/Y sky130_fd_sc_hd__nand2_2
X_12657_ _20390_/B vssd1 vssd1 vccd1 vccd1 _20723_/A sky130_fd_sc_hd__clkbuf_4
X_11608_ _11608_/A _11608_/B _11616_/B _18115_/A vssd1 vssd1 vccd1 vccd1 _11611_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ _15382_/B vssd1 vssd1 vccd1 vccd1 _15389_/C sky130_fd_sc_hd__clkbuf_2
X_18164_ _12173_/Y _12174_/X _18162_/A vssd1 vssd1 vccd1 vccd1 _18165_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18668__A2 _11980_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12588_ _12701_/A _12704_/A _12587_/Y vssd1 vssd1 vccd1 vccd1 _12588_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__20853__A _20853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17115_ _16976_/B _16934_/X _16937_/Y vssd1 vssd1 vccd1 vccd1 _17122_/A sky130_fd_sc_hd__a21boi_1
X_14327_ _11306_/X _14317_/X _14320_/X _14322_/X _13761_/B vssd1 vssd1 vccd1 vccd1
+ _14327_/X sky130_fd_sc_hd__a32o_2
XFILLER_8_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19419__A _19651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18095_ _12116_/X _12114_/X _18108_/A vssd1 vssd1 vccd1 vccd1 _18098_/B sky130_fd_sc_hd__o21ai_1
X_11539_ _15357_/A vssd1 vssd1 vccd1 vccd1 _16058_/C sky130_fd_sc_hd__buf_4
XFILLER_8_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17046_ _17042_/Y _17045_/X _17208_/B _17041_/X vssd1 vssd1 vccd1 vccd1 _17229_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15351__A1 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14258_ _14576_/A _14258_/B _14259_/B _14258_/D vssd1 vssd1 vccd1 vccd1 _14272_/A
+ sky130_fd_sc_hd__or4_1
X_13209_ _21398_/B _13456_/A _21398_/A vssd1 vssd1 vccd1 vccd1 _13210_/C sky130_fd_sc_hd__and3_1
XFILLER_48_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20227__A2 _15378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1081 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _14198_/A _14198_/B vssd1 vssd1 vccd1 vccd1 _14197_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17881__B _21019_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18840__A2 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18997_ _11511_/A _18889_/X _18890_/X _18333_/X _15887_/A vssd1 vssd1 vccd1 vccd1
+ _19007_/B sky130_fd_sc_hd__o32a_2
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16778__A _16778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19154__A _19614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17948_ _18020_/C _17948_/B vssd1 vssd1 vccd1 vccd1 _17950_/A sky130_fd_sc_hd__xnor2_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11676__B1 _15435_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17879_ _17731_/A _17927_/A _19839_/C _17733_/A vssd1 vssd1 vccd1 vccd1 _17883_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_686 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11715__A _22961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19618_ _19618_/A vssd1 vssd1 vccd1 vccd1 _19900_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20890_ _20890_/A _20890_/B _20890_/C vssd1 vssd1 vccd1 vccd1 _20891_/B sky130_fd_sc_hd__and3_1
XFILLER_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19549_ _19552_/A _19552_/C _19552_/B vssd1 vssd1 vccd1 vccd1 _19549_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13930__A _13930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22665__D _22665_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22560_ _22571_/A vssd1 vssd1 vccd1 vccd1 _22569_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__19320__C _19490_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21511_ _21485_/X _21492_/Y _21508_/B vssd1 vssd1 vccd1 vccd1 _21650_/B sky130_fd_sc_hd__o21bai_2
XFILLER_181_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22491_ _22741_/Q input48/X _22497_/S vssd1 vssd1 vccd1 vccd1 _22492_/A sky130_fd_sc_hd__mux2_1
X_21442_ _21442_/A vssd1 vssd1 vccd1 vccd1 _21522_/D sky130_fd_sc_hd__buf_2
XANTENNA__14393__A2 _14370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15590__B2 _15524_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15327__D1 _16257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19329__A _19329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21373_ _21369_/A _21369_/B _21371_/Y _21372_/X vssd1 vssd1 vccd1 vccd1 _21374_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_107_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15342__A1 _15891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20324_ _20514_/A _12420_/X _20244_/A vssd1 vssd1 vccd1 vccd1 _20324_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_162_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19048__B _19490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20255_ _20255_/A _20255_/B _20255_/C vssd1 vssd1 vccd1 vccd1 _20255_/X sky130_fd_sc_hd__or3_1
XFILLER_27_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17095__A1 _19615_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20186_ _20314_/C _20442_/A vssd1 vssd1 vccd1 vccd1 _20186_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _16157_/D vssd1 vssd1 vccd1 vccd1 _16130_/B sky130_fd_sc_hd__buf_4
XFILLER_72_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22827_ _22929_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _22827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17312__A _17312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13560_ _13677_/C _13677_/A _13677_/B vssd1 vssd1 vccd1 vccd1 _13611_/A sky130_fd_sc_hd__nand3b_1
XFILLER_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22758_ _22762_/CLK _22758_/D vssd1 vssd1 vccd1 vccd1 _22758_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_185_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12511_ _12520_/A _12518_/A _12303_/A _12550_/A vssd1 vssd1 vccd1 vccd1 _12525_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_73_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18127__B _18127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21709_ _21562_/Y _21707_/X _21708_/X _22675_/Q vssd1 vssd1 vccd1 vccd1 _21709_/X
+ sky130_fd_sc_hd__o211a_1
X_13491_ _13491_/A _13491_/B _13556_/C _13496_/B vssd1 vssd1 vccd1 vccd1 _13493_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22689_ _22690_/CLK _22689_/D vssd1 vssd1 vccd1 vccd1 _22689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11360__A _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15230_ _15230_/A _15230_/B vssd1 vssd1 vccd1 vccd1 _15231_/B sky130_fd_sc_hd__nor2_2
XFILLER_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12442_ _12457_/A vssd1 vssd1 vccd1 vccd1 _15394_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19847__A1 _19353_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15581__A1 _16016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15581__B2 _15580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15318__D1 _17532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15161_ _15161_/A _15161_/B vssd1 vssd1 vccd1 vccd1 _15163_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__13592__B1 _21874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12373_ _20089_/A _20605_/B _12579_/C vssd1 vssd1 vccd1 vccd1 _12374_/B sky130_fd_sc_hd__nand3_1
XFILLER_193_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17322__A2 _17122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14112_ _14112_/A vssd1 vssd1 vccd1 vccd1 _14963_/A sky130_fd_sc_hd__clkbuf_2
X_11324_ _11675_/A vssd1 vssd1 vccd1 vccd1 _11324_/X sky130_fd_sc_hd__buf_2
XANTENNA__15333__A1 _12576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15092_ _15092_/A _15092_/B _15092_/C vssd1 vssd1 vccd1 vccd1 _15093_/A sky130_fd_sc_hd__nand3_1
XFILLER_181_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18920_ _19091_/B _18920_/B vssd1 vssd1 vccd1 vccd1 _18920_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__20209__A2 _20210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14043_ _14043_/A _14043_/B _14043_/C vssd1 vssd1 vccd1 vccd1 _14044_/A sky130_fd_sc_hd__nand3_1
XANTENNA__18807__C1 _17525_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12698__A2 _13022_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18797__B _18797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18851_ _19013_/B _18849_/C _18330_/X _17434_/A vssd1 vssd1 vccd1 vccd1 _18861_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_133_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17802_ _17768_/A _17768_/B _17768_/C vssd1 vssd1 vccd1 vccd1 _17843_/A sky130_fd_sc_hd__o21bai_4
XFILLER_121_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18782_ _19132_/A _19132_/C vssd1 vssd1 vccd1 vccd1 _18958_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15994_ _15907_/Y _15993_/Y _15649_/X _16049_/A _17539_/D vssd1 vssd1 vccd1 vccd1
+ _16047_/D sky130_fd_sc_hd__o2111ai_4
XFILLER_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17733_ _17733_/A vssd1 vssd1 vccd1 vccd1 _17928_/D sky130_fd_sc_hd__buf_2
X_14945_ _14945_/A _15001_/A _14945_/C _15080_/C vssd1 vssd1 vccd1 vccd1 _14947_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_36_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17389__A2 _17388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17664_ _17663_/Y _17544_/Y _17541_/Y vssd1 vssd1 vccd1 vccd1 _17665_/C sky130_fd_sc_hd__a21boi_1
XFILLER_47_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14876_ _14880_/B _14877_/C _14880_/A vssd1 vssd1 vccd1 vccd1 _14947_/A sky130_fd_sc_hd__a21o_1
XFILLER_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11673__A3 _11672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19403_ _19103_/Y _19104_/X _19106_/A vssd1 vssd1 vccd1 vccd1 _19403_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16615_ _16617_/D vssd1 vssd1 vccd1 vccd1 _16615_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13827_ _14069_/A _13989_/A _14069_/C vssd1 vssd1 vccd1 vccd1 _13829_/A sky130_fd_sc_hd__nand3_2
X_17595_ _17474_/C _17474_/A _17474_/B _17484_/X vssd1 vssd1 vccd1 vccd1 _17597_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18318__A _18691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12069__C _16130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19334_ _19334_/A _19334_/B _19842_/A vssd1 vssd1 vccd1 vccd1 _19334_/X sky130_fd_sc_hd__and3_1
X_16546_ _16524_/Y _16545_/Y _16530_/D vssd1 vssd1 vccd1 vccd1 _16546_/Y sky130_fd_sc_hd__o21ai_2
X_13758_ _13707_/A _13707_/B _13773_/A _13766_/A vssd1 vssd1 vccd1 vccd1 _13948_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__21342__B1 _21767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12709_ _12700_/Y _12705_/X _12950_/C vssd1 vssd1 vccd1 vccd1 _12709_/Y sky130_fd_sc_hd__o21ai_1
X_19265_ _11345_/X _11351_/X _19941_/A _19941_/B _12064_/X vssd1 vssd1 vccd1 vccd1
+ _19265_/X sky130_fd_sc_hd__o32a_1
XFILLER_148_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16477_ _16477_/A _16477_/B _16477_/C vssd1 vssd1 vccd1 vccd1 _16513_/A sky130_fd_sc_hd__and3_1
X_13689_ _13689_/A _13689_/B vssd1 vssd1 vccd1 vccd1 _22929_/D sky130_fd_sc_hd__nand2_1
XFILLER_188_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17561__A2 _16580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11270__A _22786_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18216_ _18216_/A _18216_/B vssd1 vssd1 vccd1 vccd1 _18219_/A sky130_fd_sc_hd__nand2_1
X_15428_ _15718_/A vssd1 vssd1 vccd1 vccd1 _15933_/A sky130_fd_sc_hd__clkbuf_4
X_19196_ _18156_/X _17635_/A _18282_/X _19194_/Y _19195_/Y vssd1 vssd1 vccd1 vccd1
+ _19201_/B sky130_fd_sc_hd__o221ai_4
XFILLER_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16780__B _18797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18147_ _18172_/A vssd1 vssd1 vccd1 vccd1 _18383_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15046__C_N _15175_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15359_ _22699_/Q vssd1 vssd1 vccd1 vccd1 _15369_/C sky130_fd_sc_hd__inv_2
XFILLER_191_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18078_ _18015_/C _18051_/Y _18053_/Y _18077_/Y vssd1 vssd1 vccd1 vccd1 _18079_/B
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__15396__B _18130_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17029_ _16733_/Y _16740_/Y _16853_/C _16848_/X vssd1 vssd1 vccd1 vccd1 _17031_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_171_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19066__A2 _11308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20040_ _20037_/B _20012_/X _20013_/X _20039_/Y vssd1 vssd1 vccd1 vccd1 _20041_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__21948__A2 _21594_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21991_ _21987_/A _21988_/X _21990_/X vssd1 vssd1 vccd1 vccd1 _22075_/B sky130_fd_sc_hd__a21bo_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21861__B _21963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20942_ _20941_/A _20941_/B _20941_/C vssd1 vssd1 vccd1 vccd1 _20945_/B sky130_fd_sc_hd__a21o_1
XFILLER_94_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14162__A1_N _14147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ _12379_/A _12379_/B _12761_/X vssd1 vssd1 vccd1 vccd1 _20873_/X sky130_fd_sc_hd__a21o_1
XANTENNA__20435__A2_N _20554_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22612_ _22612_/A vssd1 vssd1 vccd1 vccd1 _22794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22543_ _14366_/X input38/X _22547_/S vssd1 vssd1 vccd1 vccd1 _22544_/A sky130_fd_sc_hd__mux2_1
XANTENNA__20687__A2 _15935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15563__A1 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22474_ _22474_/A vssd1 vssd1 vccd1 vccd1 _22733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16690__B _22891_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21425_ _21559_/A _21424_/C _21424_/A vssd1 vssd1 vccd1 vccd1 _21426_/C sky130_fd_sc_hd__a21o_1
XFILLER_182_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15315__A1 _15714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15315__B2 _18680_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21356_ _21346_/X _21198_/Y _21204_/Y _21211_/A _21237_/Y vssd1 vssd1 vccd1 vccd1
+ _21359_/A sky130_fd_sc_hd__a32o_1
XFILLER_136_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20307_ _20432_/B vssd1 vssd1 vccd1 vccd1 _20553_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21287_ _21423_/A vssd1 vssd1 vccd1 vccd1 _21559_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20238_ _20093_/A _20093_/B _20107_/C vssd1 vssd1 vccd1 vccd1 _20238_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15079__B1 _15182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16815__A1 _19461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15618__A2 _15905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17307__A _17307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16815__B2 _18839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20169_ _20169_/A _20169_/B vssd1 vssd1 vccd1 vccd1 _20170_/C sky130_fd_sc_hd__nand2_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12991_ _12954_/C _12954_/A _12954_/B _12937_/A _12958_/C vssd1 vssd1 vccd1 vccd1
+ _12991_/X sky130_fd_sc_hd__a32o_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11355__A _22968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11942_ _11942_/A _18107_/B _18107_/C vssd1 vssd1 vccd1 vccd1 _11943_/B sky130_fd_sc_hd__and3_1
X_14730_ _14727_/X _14728_/X _14729_/Y vssd1 vssd1 vccd1 vccd1 _14731_/C sky130_fd_sc_hd__o21ai_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14548_/A _14661_/B _14661_/C vssd1 vssd1 vccd1 vccd1 _14661_/Y sky130_fd_sc_hd__nand3b_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11873_ _12074_/A _12074_/B _11874_/A vssd1 vssd1 vccd1 vccd1 _11873_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17791__A2 _18044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16400_ _16400_/A _21050_/D _16400_/C vssd1 vssd1 vccd1 vccd1 _16400_/X sky130_fd_sc_hd__and3_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13570__A _21739_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13612_ _13612_/A _13612_/B vssd1 vssd1 vccd1 vccd1 _13612_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17380_ _17380_/A vssd1 vssd1 vccd1 vccd1 _17380_/X sky130_fd_sc_hd__buf_4
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _14729_/A _14605_/D _14591_/X vssd1 vssd1 vccd1 vccd1 _14712_/A sky130_fd_sc_hd__a21oi_1
XFILLER_164_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_823 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13543_ _13543_/A _13543_/B _13543_/C vssd1 vssd1 vccd1 vccd1 _13548_/A sky130_fd_sc_hd__nand3_1
X_16331_ _16331_/A vssd1 vssd1 vccd1 vccd1 _16745_/A sky130_fd_sc_hd__buf_2
XFILLER_38_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18740__A1 _18666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19050_ _18371_/X _16799_/X _19062_/A vssd1 vssd1 vccd1 vccd1 _19231_/A sky130_fd_sc_hd__o21ai_1
X_16262_ _16258_/Y _16261_/Y _11820_/A _15723_/A vssd1 vssd1 vccd1 vccd1 _16263_/D
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__15554__A1 _12913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13474_ _13471_/Y _13473_/X _13537_/B vssd1 vssd1 vccd1 vccd1 _13474_/X sky130_fd_sc_hd__o21a_1
XFILLER_185_355 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18001_ _18048_/C _17910_/Y _17960_/D vssd1 vssd1 vccd1 vccd1 _18045_/A sky130_fd_sc_hd__a21boi_1
XFILLER_139_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15213_ _15213_/A vssd1 vssd1 vccd1 vccd1 _15238_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12425_ _12734_/A _12420_/X _12461_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _12425_/X
+ sky130_fd_sc_hd__o22a_1
X_16193_ _16192_/X _15978_/X _16043_/C _16090_/Y _16188_/Y vssd1 vssd1 vccd1 vccd1
+ _16195_/B sky130_fd_sc_hd__o221ai_2
XFILLER_166_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15144_ _15134_/A _15132_/Y _15133_/A vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__a21oi_1
X_12356_ _15633_/B _12813_/A vssd1 vssd1 vccd1 vccd1 _15409_/A sky130_fd_sc_hd__nand2_2
XFILLER_5_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11307_ _11377_/A _11420_/A _11306_/X vssd1 vssd1 vccd1 vccd1 _11308_/B sky130_fd_sc_hd__o21ai_4
X_19952_ _19991_/A _19952_/B _19991_/B vssd1 vssd1 vccd1 vccd1 _19954_/A sky130_fd_sc_hd__and3_1
X_15075_ _15074_/B _15074_/C _15074_/A vssd1 vssd1 vccd1 vccd1 _15076_/C sky130_fd_sc_hd__o21ai_1
XFILLER_126_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12287_ _22703_/Q vssd1 vssd1 vccd1 vccd1 _12288_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__11328__C1 _11860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18903_ _18891_/X _18893_/X _19085_/A _19009_/A vssd1 vssd1 vccd1 vccd1 _18907_/B
+ sky130_fd_sc_hd__o211ai_1
X_14026_ _14061_/A _14026_/B _14026_/C _14026_/D vssd1 vssd1 vccd1 vccd1 _14043_/C
+ sky130_fd_sc_hd__nand4_1
X_19883_ _19750_/X _19880_/Y _19881_/X _19882_/Y vssd1 vssd1 vccd1 vccd1 _19885_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__18320__B _18512_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__D _16157_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16759__C _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18834_ _18835_/C _19112_/A _18833_/Y vssd1 vssd1 vccd1 vccd1 _18929_/A sky130_fd_sc_hd__a21o_1
XFILLER_121_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18008__B1 _22904_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18765_ _18765_/A _18765_/B vssd1 vssd1 vccd1 vccd1 _18765_/X sky130_fd_sc_hd__and2_1
X_15977_ _16011_/A vssd1 vssd1 vccd1 vccd1 _15977_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15382__D _17530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20528__A1_N _20378_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17716_ _17716_/A _17716_/B vssd1 vssd1 vccd1 vccd1 _17720_/C sky130_fd_sc_hd__nor2_1
XANTENNA__15960__A _15960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14928_ _14928_/A _14929_/C vssd1 vssd1 vccd1 vccd1 _22677_/D sky130_fd_sc_hd__xor2_1
X_18696_ _18877_/A vssd1 vssd1 vccd1 vccd1 _18696_/X sky130_fd_sc_hd__buf_2
XFILLER_48_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_656 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17647_ _17647_/A vssd1 vssd1 vccd1 vccd1 _17817_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14859_ _14859_/A vssd1 vssd1 vccd1 vccd1 _15050_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19508__B1 _19651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20728__D _20818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17578_ _17578_/A _17628_/A _17580_/A vssd1 vssd1 vccd1 vccd1 _17579_/C sky130_fd_sc_hd__nand3_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19317_ _19317_/A _19329_/B _19461_/C _19317_/D vssd1 vssd1 vccd1 vccd1 _19317_/Y
+ sky130_fd_sc_hd__nand4_2
X_16529_ _16530_/D _16529_/B _16529_/C vssd1 vssd1 vccd1 vccd1 _16529_/X sky130_fd_sc_hd__and3_1
XANTENNA__11712__B _11712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19248_ _19248_/A _19248_/B vssd1 vssd1 vccd1 vccd1 _19248_/Y sky130_fd_sc_hd__nand2_2
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19179_ _19179_/A _19179_/B _19179_/C vssd1 vssd1 vccd1 vccd1 _19190_/B sky130_fd_sc_hd__nand3_2
XFILLER_145_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11567__C1 _11566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21210_ _21210_/A _21210_/B _21210_/C vssd1 vssd1 vccd1 vccd1 _21211_/A sky130_fd_sc_hd__nand3_1
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22190_ _22190_/A _22190_/B _22219_/B _22190_/D vssd1 vssd1 vccd1 vccd1 _22192_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19692__C1 _19461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15557__D _20133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21141_ _21141_/A _21141_/B _22944_/Q vssd1 vssd1 vccd1 vccd1 _21150_/C sky130_fd_sc_hd__or3b_1
XFILLER_120_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21072_ _22941_/Q vssd1 vssd1 vccd1 vccd1 _21072_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18798__A1 _18156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20023_ _20024_/A _20024_/B _20024_/C vssd1 vssd1 vccd1 vccd1 _20042_/B sky130_fd_sc_hd__a21o_1
XFILLER_141_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16273__A2 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15870__A _17039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21591__B _21591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21974_ _21964_/X _21958_/X _21725_/Y _21854_/X _21973_/X vssd1 vssd1 vccd1 vccd1
+ _22030_/B sky130_fd_sc_hd__o32a_1
XFILLER_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19061__B _19199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20925_ _20923_/B _20923_/C _20923_/A vssd1 vssd1 vccd1 vccd1 _20925_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11903__A _11909_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12047__B1 _22660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20109__A1 _12680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20856_ _20782_/B _20854_/Y _20913_/A _20855_/Y _17525_/C vssd1 vssd1 vccd1 vccd1
+ _20860_/B sky130_fd_sc_hd__o2111ai_4
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22918__CLK _22922_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20787_ _20706_/X _20787_/B _20787_/C vssd1 vssd1 vccd1 vccd1 _20871_/A sky130_fd_sc_hd__nand3b_2
XFILLER_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22526_ _22526_/A vssd1 vssd1 vccd1 vccd1 _22756_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__22853__D _22865_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16733__B1 _16732_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22457_ _22457_/A vssd1 vssd1 vccd1 vccd1 _22725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12210_ _12210_/A _22662_/B vssd1 vssd1 vccd1 vccd1 _12211_/A sky130_fd_sc_hd__nand2_2
XFILLER_109_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21408_ _21266_/A _21266_/B _21265_/Y vssd1 vssd1 vccd1 vccd1 _21410_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__21085__A2 _17839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13190_ _13110_/Y _21580_/A _13131_/X vssd1 vssd1 vccd1 vccd1 _13450_/A sky130_fd_sc_hd__a21o_1
XFILLER_163_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22388_ _22388_/A vssd1 vssd1 vccd1 vccd1 _22695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12141_ _11361_/A _18655_/A _12134_/A vssd1 vssd1 vccd1 vccd1 _12143_/B sky130_fd_sc_hd__o21ai_1
XFILLER_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19517__A _19517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21339_ _21725_/A _21725_/B _21498_/B _21454_/A _21739_/B vssd1 vssd1 vccd1 vccd1
+ _21348_/A sky130_fd_sc_hd__a32o_1
XFILLER_163_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12072_ _17006_/D vssd1 vssd1 vccd1 vccd1 _17039_/D sky130_fd_sc_hd__buf_2
XANTENNA__14511__A2 _14834_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18778__D _18778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18140__B _18691_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19986__B1 _18023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15900_ _15900_/A _15900_/B vssd1 vssd1 vccd1 vccd1 _15900_/Y sky130_fd_sc_hd__nand2_2
XFILLER_173_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16880_ _17039_/D _21050_/D _17039_/C _17039_/A vssd1 vssd1 vccd1 vccd1 _16880_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_131_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17461__A1 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _16809_/B vssd1 vssd1 vccd1 vccd1 _17385_/B sky130_fd_sc_hd__buf_2
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14275__A1 _14998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _18519_/Y _18523_/Y _18527_/Y vssd1 vssd1 vccd1 vccd1 _18557_/B sky130_fd_sc_hd__o21ai_1
XFILLER_18_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _16402_/A vssd1 vssd1 vccd1 vccd1 _16209_/A sky130_fd_sc_hd__clkbuf_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _20792_/C _16067_/B _16067_/D _13016_/C vssd1 vssd1 vccd1 vccd1 _12975_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20398__A _20398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17501_ _17507_/A _17853_/A _17959_/C _22898_/Q vssd1 vssd1 vccd1 vccd1 _17501_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _14712_/Y _14600_/Y _14580_/X vssd1 vssd1 vccd1 vccd1 _14714_/C sky130_fd_sc_hd__a21oi_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18481_ _18337_/X _18343_/X _18340_/Y _18349_/B vssd1 vssd1 vccd1 vccd1 _18490_/A
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_73_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11925_ _11897_/Y _11900_/Y _12079_/C _11924_/X vssd1 vssd1 vccd1 vccd1 _11927_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _15693_/A _15693_/B vssd1 vssd1 vccd1 vccd1 _15698_/A sky130_fd_sc_hd__nor2_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12909__A _20207_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17432_ _17129_/Y _17237_/Y _17238_/X _17236_/X vssd1 vssd1 vccd1 vccd1 _17433_/C
+ sky130_fd_sc_hd__o22ai_4
XFILLER_127_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ _15991_/D vssd1 vssd1 vccd1 vccd1 _16564_/B sky130_fd_sc_hd__clkbuf_4
X_14644_ _13948_/X _13949_/X _14646_/A _14646_/B _14560_/A vssd1 vssd1 vccd1 vccd1
+ _14750_/B sky130_fd_sc_hd__a221o_1
XFILLER_127_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17363_ _17361_/Y _17959_/C _17372_/C vssd1 vssd1 vccd1 vccd1 _17616_/A sky130_fd_sc_hd__a21oi_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14575_ _14575_/A _14575_/B _15010_/A vssd1 vssd1 vccd1 vccd1 _14602_/B sky130_fd_sc_hd__nand3_1
XFILLER_82_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11787_ _11782_/Y _12165_/A _11786_/X _11779_/X _11945_/A vssd1 vssd1 vccd1 vccd1
+ _11809_/B sky130_fd_sc_hd__o311a_2
X_19102_ _18829_/X _18830_/X _18819_/A _19079_/A vssd1 vssd1 vccd1 vccd1 _19104_/C
+ sky130_fd_sc_hd__o31a_1
X_16314_ _15638_/X _16312_/X _16313_/X vssd1 vssd1 vccd1 vccd1 _16314_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_119_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13526_ _13526_/A _13526_/B vssd1 vssd1 vccd1 vccd1 _13526_/X sky130_fd_sc_hd__or2_1
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17294_ _17293_/Y _17286_/X _17290_/B vssd1 vssd1 vccd1 vccd1 _17294_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14843__B _14843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19033_ _19004_/Y _19010_/X _19028_/X _19032_/Y vssd1 vssd1 vccd1 vccd1 _19033_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_146_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16245_ _15804_/C _16530_/C _19507_/C _16234_/X vssd1 vssd1 vccd1 vccd1 _16250_/A
+ sky130_fd_sc_hd__a31o_1
X_13457_ _21177_/A _21498_/D _21498_/B _13579_/A vssd1 vssd1 vccd1 vccd1 _13457_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_174_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12408_ _16319_/A vssd1 vssd1 vccd1 vccd1 _15631_/A sky130_fd_sc_hd__buf_4
XANTENNA__20808__C1 _15935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16176_ _16186_/A _16186_/B _16175_/Y vssd1 vssd1 vccd1 vccd1 _16176_/Y sky130_fd_sc_hd__o21ai_1
X_13388_ _13339_/Y _13353_/Y _13359_/X _13387_/X vssd1 vssd1 vccd1 vccd1 _13392_/B
+ sky130_fd_sc_hd__o211ai_1
Xoutput106 _14428_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_86_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput117 _22665_/Q vssd1 vssd1 vccd1 vccd1 y[1] sky130_fd_sc_hd__buf_2
XFILLER_115_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11564__A2 _18371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15127_ _15128_/A _15128_/B _15128_/C _15128_/D vssd1 vssd1 vccd1 vccd1 _15129_/A
+ sky130_fd_sc_hd__a22oi_2
X_12339_ _16319_/A _12402_/A _15631_/C _12361_/A vssd1 vssd1 vccd1 vccd1 _12339_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_142_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19935_ _19935_/A vssd1 vssd1 vccd1 vccd1 _22903_/D sky130_fd_sc_hd__clkbuf_1
X_15058_ _15058_/A _15058_/B _15058_/C vssd1 vssd1 vccd1 vccd1 _15058_/X sky130_fd_sc_hd__and3_1
XFILLER_141_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21233__C1 _21944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14009_ _14497_/A _14009_/B _14009_/C _14009_/D vssd1 vssd1 vccd1 vccd1 _14033_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_68_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16489__C _16771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19866_ _19866_/A _19866_/B vssd1 vssd1 vccd1 vccd1 _19866_/X sky130_fd_sc_hd__and2_1
XFILLER_96_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19441__A2 _19294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18985__B _19481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18817_ _18825_/A _19079_/A vssd1 vssd1 vccd1 vccd1 _18819_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19797_ _19615_/A _19795_/X _19790_/Y _19796_/X vssd1 vssd1 vccd1 vccd1 _19798_/C
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__15999__D1 _15577_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15690__A _16257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18748_ _18748_/A _18748_/B vssd1 vssd1 vccd1 vccd1 _18748_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18679_ _18841_/A _22798_/Q _18679_/C vssd1 vssd1 vccd1 vccd1 _18858_/A sky130_fd_sc_hd__nand3_2
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11723__A _16447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20710_ _20718_/A _20713_/B _20720_/B _20720_/C vssd1 vssd1 vccd1 vccd1 _20710_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21690_ _22167_/A _13434_/X _21539_/B _21524_/A vssd1 vssd1 vccd1 vccd1 _21809_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20641_ _20567_/Y _20568_/X _20636_/Y _20640_/Y vssd1 vssd1 vccd1 vccd1 _20650_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_149_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18506__A _18876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20572_ _20575_/B vssd1 vssd1 vccd1 vccd1 _20734_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22311_ _22302_/A _22302_/Y _22310_/X vssd1 vssd1 vccd1 vccd1 _22313_/A sky130_fd_sc_hd__o21ai_1
XFILLER_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22264__A1 _22231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22242_ _22243_/B _22243_/A vssd1 vssd1 vccd1 vccd1 _22244_/A sky130_fd_sc_hd__nor2_1
XFILLER_192_678 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12273__B _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20275__B1 _20125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15865__A _16192_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22173_ _22173_/A _22173_/B _22304_/B _22173_/D vssd1 vssd1 vccd1 vccd1 _22238_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_106_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11960__C1 _12219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21124_ _21124_/A _21124_/B vssd1 vssd1 vccd1 vccd1 _21130_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17428__D1 _20854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21055_ _21055_/A _21055_/B vssd1 vssd1 vccd1 vccd1 _21061_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__20578__A1 _12967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20006_ _20024_/B _20026_/B _20005_/A vssd1 vssd1 vccd1 vccd1 _20008_/B sky130_fd_sc_hd__a21oi_1
XFILLER_189_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19196__A1 _18156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14928__B _14929_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17304__B _17304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21957_ _21957_/A _22037_/C vssd1 vssd1 vccd1 vccd1 _21957_/Y sky130_fd_sc_hd__nor2_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11633__A _11633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ _11938_/A vssd1 vssd1 vccd1 vccd1 _11935_/C sky130_fd_sc_hd__clkbuf_2
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20908_ _20891_/A _20891_/B _20842_/X vssd1 vssd1 vccd1 vccd1 _20908_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_743 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12690_ _12682_/X _20793_/B _16067_/D _12689_/X vssd1 vssd1 vccd1 vccd1 _13007_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_153_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21888_ _21891_/A _21891_/B _21892_/B _21892_/C vssd1 vssd1 vccd1 vccd1 _21889_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12448__B _16257_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11636_/X _11606_/X _11639_/X _11745_/B _11623_/X vssd1 vssd1 vccd1 vccd1
+ _11641_/X sky130_fd_sc_hd__o311a_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _20839_/A _20839_/B vssd1 vssd1 vccd1 vccd1 _22916_/D sky130_fd_sc_hd__xnor2_2
XANTENNA__19499__A2 _16799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22890__CLK _22952_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14360_ _22795_/Q vssd1 vssd1 vccd1 vccd1 _18128_/C sky130_fd_sc_hd__buf_2
X_11572_ _18303_/C vssd1 vssd1 vccd1 vccd1 _11664_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_156_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13311_ _21495_/A _21476_/C _13311_/C vssd1 vssd1 vccd1 vccd1 _21202_/A sky130_fd_sc_hd__nand3_2
XFILLER_128_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 wb_adr_i[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_1
X_22509_ _22509_/A vssd1 vssd1 vccd1 vccd1 _22749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ _14180_/B _14180_/C _14180_/A vssd1 vssd1 vccd1 vccd1 _14291_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16030_ _16093_/A _16134_/B _16133_/B vssd1 vssd1 vccd1 vccd1 _16030_/Y sky130_fd_sc_hd__a21boi_1
X_13242_ _22720_/Q vssd1 vssd1 vccd1 vccd1 _13623_/A sky130_fd_sc_hd__buf_2
XFILLER_196_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input73_A x[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15775__A _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ _13449_/A _13449_/B _13519_/B vssd1 vssd1 vccd1 vccd1 _13173_/Y sky130_fd_sc_hd__nand3_1
XFILLER_184_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12124_ _12184_/A vssd1 vssd1 vccd1 vccd1 _18208_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_184_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17981_ _21044_/B _18023_/A _19983_/B _17981_/D vssd1 vssd1 vccd1 vccd1 _18030_/C
+ sky130_fd_sc_hd__or4_2
X_19720_ _19719_/X _19799_/B _19720_/C vssd1 vssd1 vccd1 vccd1 _19725_/C sky130_fd_sc_hd__nand3b_1
XFILLER_133_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1032 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16932_ _18445_/A _17129_/B _16932_/C _20502_/B vssd1 vssd1 vccd1 vccd1 _16932_/Y
+ sky130_fd_sc_hd__nand4_4
X_12055_ _12055_/A _12055_/B vssd1 vssd1 vccd1 vccd1 _12055_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__19423__A2 _18023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_707 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12630__C _12630_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19651_ _19651_/A _19651_/B _19651_/C _19945_/B vssd1 vssd1 vccd1 vccd1 _19652_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__18631__B1 _19504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18092__D1 _15810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16863_ _16848_/X _16853_/B _16853_/C vssd1 vssd1 vccd1 vccd1 _16863_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_78_887 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18602_ _19281_/A _18430_/A _18601_/Y vssd1 vssd1 vccd1 vccd1 _18602_/Y sky130_fd_sc_hd__a21oi_1
X_15814_ _15406_/X _15813_/Y _15795_/X vssd1 vssd1 vccd1 vccd1 _15814_/Y sky130_fd_sc_hd__a21oi_1
X_19582_ _19687_/D vssd1 vssd1 vccd1 vccd1 _19836_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__15996__A1 _15797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16794_ _16972_/A _16971_/A _16803_/A _16803_/B vssd1 vssd1 vccd1 vccd1 _16796_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18533_ _19194_/D _19465_/A _19317_/D _19199_/A vssd1 vssd1 vccd1 vccd1 _18533_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__21017__A _21017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _15693_/A _15693_/B _15743_/X _15744_/Y vssd1 vssd1 vccd1 vccd1 _15748_/B
+ sky130_fd_sc_hd__o22ai_2
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _12957_/A _12957_/B _12957_/C vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__nand3_1
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18029__C _20012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18464_ _18464_/A vssd1 vssd1 vccd1 vccd1 _18770_/C sky130_fd_sc_hd__buf_2
X_11908_ _11909_/C _11909_/A _11782_/Y _11907_/Y vssd1 vssd1 vccd1 vccd1 _12077_/D
+ sky130_fd_sc_hd__o2bb2ai_1
X_15676_ _15859_/C _15679_/B _15676_/C _15676_/D vssd1 vssd1 vccd1 vccd1 _15681_/C
+ sky130_fd_sc_hd__nand4_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20741__A1 _20818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12776_/X _12886_/X _12887_/X _12868_/X _20169_/A vssd1 vssd1 vccd1 vccd1
+ _12889_/C sky130_fd_sc_hd__o2111ai_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _17399_/Y _17410_/X _17413_/Y _17414_/X vssd1 vssd1 vccd1 vccd1 _17416_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_14627_ _14623_/X _14625_/X _14626_/Y vssd1 vssd1 vccd1 vccd1 _14635_/B sky130_fd_sc_hd__o21ai_2
X_18395_ _18404_/A _18395_/B _18395_/C vssd1 vssd1 vccd1 vccd1 _18395_/X sky130_fd_sc_hd__and3_1
X_11839_ _11839_/A vssd1 vssd1 vccd1 vccd1 _11902_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20575__B _20575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17346_ _17345_/X _17330_/Y _17340_/Y vssd1 vssd1 vccd1 vccd1 _17346_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_147_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14558_ _14544_/A _14544_/B _14544_/C _14547_/B _14547_/A vssd1 vssd1 vccd1 vccd1
+ _14758_/C sky130_fd_sc_hd__a32oi_4
XFILLER_14_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _13664_/B _22106_/A _13664_/D _22108_/C vssd1 vssd1 vccd1 vccd1 _13509_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17277_ _14431_/A _15808_/A _11672_/A _20781_/A _20781_/B vssd1 vssd1 vccd1 vccd1
+ _17277_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_146_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14489_ _15006_/A _14489_/B _14489_/C _15006_/C vssd1 vssd1 vccd1 vccd1 _14494_/B
+ sky130_fd_sc_hd__nand4_4
X_19016_ _19016_/A _19016_/B _19016_/C vssd1 vssd1 vccd1 vccd1 _19016_/Y sky130_fd_sc_hd__nand3_4
X_16228_ _16482_/A _22965_/Q _16242_/B vssd1 vssd1 vccd1 vccd1 _16228_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__21049__A2 _17839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15920__B2 _15919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ _16157_/C _16997_/C _16166_/B _16160_/A vssd1 vssd1 vccd1 vccd1 _16159_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_1082 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19918_ _19922_/A _19922_/B vssd1 vssd1 vccd1 vccd1 _19919_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__17108__C _20593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12540__C _12540_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16228__A2 _22965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17425__A1 _17421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19849_ _19850_/B _19850_/C _19850_/A vssd1 vssd1 vccd1 vccd1 _19851_/A sky130_fd_sc_hd__a21o_1
XANTENNA__17425__B2 _17424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16947__C _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22860_ _22943_/CLK _22872_/Q vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21811_ _21807_/Y _21808_/X _21810_/Y vssd1 vssd1 vccd1 vccd1 _21837_/C sky130_fd_sc_hd__o21ai_2
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19717__A3 _19793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_762 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22791_ _22791_/CLK _22791_/D vssd1 vssd1 vccd1 vccd1 _22791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1020 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19042__D _19202_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21742_ _21742_/A _21742_/B vssd1 vssd1 vccd1 vccd1 _21742_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20732__A1 _20818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17456__A1_N _17304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21673_ _21618_/Y _21624_/Y _21662_/B _21647_/Y vssd1 vssd1 vccd1 vccd1 _21673_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__17140__A _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20624_ _20455_/X _20459_/Y _20485_/Y _20490_/Y vssd1 vssd1 vccd1 vccd1 _20624_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20555_ _20834_/A _20835_/A _20548_/X _20551_/Y _20554_/Y vssd1 vssd1 vccd1 vccd1
+ _20566_/A sky130_fd_sc_hd__o2111a_1
XFILLER_138_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20486_ _20605_/A _20608_/C _20486_/C vssd1 vssd1 vccd1 vccd1 _20486_/X sky130_fd_sc_hd__and3_1
XFILLER_152_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12725__A1 _12602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22225_ _22108_/Y _22181_/Y _22304_/A _22183_/Y _22265_/C vssd1 vssd1 vccd1 vccd1
+ _22225_/Y sky130_fd_sc_hd__o2111ai_2
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22156_ _22156_/A _22156_/B vssd1 vssd1 vccd1 vccd1 _22212_/B sky130_fd_sc_hd__nand2_1
XFILLER_160_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11628__A _18716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21107_ _21138_/A vssd1 vssd1 vccd1 vccd1 _21107_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22087_ _22142_/B _22090_/B _22145_/A _22145_/B _22155_/A vssd1 vssd1 vccd1 vccd1
+ _22092_/A sky130_fd_sc_hd__a221o_1
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16219__A2 _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21038_ _21039_/A _21039_/B _22940_/Q vssd1 vssd1 vccd1 vccd1 _21076_/C sky130_fd_sc_hd__a21o_1
XFILLER_75_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17315__A _17523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13860_ _13930_/A _13930_/B _13923_/A vssd1 vssd1 vccd1 vccd1 _13862_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20971__A1 _15355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19169__A1 _12118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12811_ _12852_/A vssd1 vssd1 vccd1 vccd1 _20120_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12459__A _16465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13791_ _14044_/B vssd1 vssd1 vccd1 vccd1 _15082_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15530_ _15530_/A vssd1 vssd1 vccd1 vccd1 _15530_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20098__D _20098_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12742_ _12742_/A _12742_/B vssd1 vssd1 vccd1 vccd1 _13007_/D sky130_fd_sc_hd__nor2_1
XANTENNA__17969__B _22903_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15461_ _15461_/A _15461_/B vssd1 vssd1 vccd1 vccd1 _15461_/Y sky130_fd_sc_hd__nand2_1
X_12673_ _12968_/B _12671_/X _20514_/A _12719_/A vssd1 vssd1 vccd1 vccd1 _12742_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17200_/A _17200_/B _17200_/C vssd1 vssd1 vccd1 vccd1 _17200_/Y sky130_fd_sc_hd__nand3_1
XFILLER_24_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11624_ _18810_/D _18328_/A _11614_/Y _11623_/X vssd1 vssd1 vccd1 vccd1 _11647_/C
+ sky130_fd_sc_hd__a22o_1
X_14412_ _22442_/B vssd1 vssd1 vccd1 vccd1 _14412_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18180_ _12189_/A _18208_/B _12182_/D _12185_/Y vssd1 vssd1 vccd1 vccd1 _18181_/C
+ sky130_fd_sc_hd__a31oi_1
X_15392_ _15664_/A _15665_/A _15392_/C vssd1 vssd1 vccd1 vccd1 _15512_/C sky130_fd_sc_hd__nand3_2
XFILLER_196_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19341__A1 _19336_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17131_ _19587_/A _17131_/B vssd1 vssd1 vccd1 vccd1 _17131_/Y sky130_fd_sc_hd__nand2_1
X_11555_ _22957_/Q _22958_/Q vssd1 vssd1 vccd1 vccd1 _11712_/C sky130_fd_sc_hd__nor2_2
XANTENNA__17985__A _19419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14343_ _13799_/X _14330_/X _14337_/X _13055_/A _14342_/X vssd1 vssd1 vccd1 vccd1
+ _14343_/X sky130_fd_sc_hd__a221o_1
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17062_ _17061_/X _16672_/X _16660_/Y _17215_/B vssd1 vssd1 vccd1 vccd1 _17371_/A
+ sky130_fd_sc_hd__o211ai_4
X_14274_ _14274_/A vssd1 vssd1 vccd1 vccd1 _14998_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ _11418_/A _11349_/X _11772_/A vssd1 vssd1 vccd1 vccd1 _11608_/B sky130_fd_sc_hd__o21ai_1
XFILLER_137_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16560__D1 _15711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16013_ _16007_/X _16008_/Y _16009_/Y _16012_/Y vssd1 vssd1 vccd1 vccd1 _16133_/A
+ sky130_fd_sc_hd__o211ai_2
X_13225_ _21383_/A _13162_/C _13162_/A _13384_/B _13385_/A vssd1 vssd1 vccd1 vccd1
+ _13225_/X sky130_fd_sc_hd__o311a_1
XANTENNA__12922__A _16059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17655__A1 _17739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16458__A2 _18797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ _21212_/C _21367_/A _21367_/B _21362_/B _21351_/C vssd1 vssd1 vccd1 vccd1
+ _13385_/A sky130_fd_sc_hd__a32o_2
XFILLER_3_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12107_/A _12107_/B _12107_/C vssd1 vssd1 vccd1 vccd1 _12108_/B sky130_fd_sc_hd__nand3_1
XFILLER_112_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11538__A _11583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _17910_/A _17910_/B _17910_/C _17910_/D _17502_/X vssd1 vssd1 vccd1 vccd1
+ _17964_/Y sky130_fd_sc_hd__a41oi_2
XFILLER_112_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13087_ _13087_/A vssd1 vssd1 vccd1 vccd1 _13105_/A sky130_fd_sc_hd__buf_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19703_ _19703_/A _19703_/B _19703_/C vssd1 vssd1 vccd1 vccd1 _19708_/A sky130_fd_sc_hd__nand3_1
X_16915_ _16275_/A _15919_/A _16914_/Y vssd1 vssd1 vccd1 vccd1 _16915_/Y sky130_fd_sc_hd__o21ai_2
X_12038_ _12055_/A _12055_/B _12088_/B vssd1 vssd1 vccd1 vccd1 _12039_/C sky130_fd_sc_hd__nand3_1
XANTENNA__21203__A2 _13305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22400__A1 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17895_ _17895_/A _17895_/B _17895_/C vssd1 vssd1 vccd1 vccd1 _17896_/B sky130_fd_sc_hd__nand3_1
XFILLER_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19634_ _19611_/X _19634_/B _19634_/C _19724_/A vssd1 vssd1 vccd1 vccd1 _19724_/B
+ sky130_fd_sc_hd__nand4b_4
XANTENNA__13753__A _22865_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16846_ _16846_/A _16846_/B _16846_/C vssd1 vssd1 vccd1 vccd1 _16866_/A sky130_fd_sc_hd__nand3_2
XFILLER_168_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16091__B1 _16011_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19565_ _19555_/C _19563_/Y _19564_/Y vssd1 vssd1 vccd1 vccd1 _19565_/Y sky130_fd_sc_hd__a21oi_2
X_16777_ _16777_/A vssd1 vssd1 vccd1 vccd1 _16971_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12101__C1 _17280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13989_ _13989_/A vssd1 vssd1 vccd1 vccd1 _14786_/B sky130_fd_sc_hd__buf_2
XFILLER_81_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18516_ _11511_/A _11786_/X _12001_/B _18514_/Y _18653_/A vssd1 vssd1 vccd1 vccd1
+ _18526_/B sky130_fd_sc_hd__o221ai_4
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ _15988_/B _16781_/B _16308_/C vssd1 vssd1 vccd1 vccd1 _15728_/X sky130_fd_sc_hd__and3_1
XFILLER_34_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19496_ _19496_/A _19496_/B _19496_/C vssd1 vssd1 vccd1 vccd1 _19497_/B sky130_fd_sc_hd__and3_1
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18447_ _11634_/A _17635_/A _18451_/A _18451_/B vssd1 vssd1 vccd1 vccd1 _18450_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_179_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15659_ _15616_/X _15657_/Y _15658_/Y vssd1 vssd1 vccd1 vccd1 _15660_/B sky130_fd_sc_hd__o21ai_1
XFILLER_178_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14584__A _22764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22467__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18378_ _18726_/A _18520_/B _18520_/A vssd1 vssd1 vccd1 vccd1 _18381_/A sky130_fd_sc_hd__a21o_1
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17329_ _17486_/A _17486_/B _17486_/C vssd1 vssd1 vccd1 vccd1 _17485_/B sky130_fd_sc_hd__a21o_1
XFILLER_146_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20340_ _12450_/X _15611_/A _20339_/Y vssd1 vssd1 vccd1 vccd1 _20340_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_135_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21690__A2 _13434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18503__B _18678_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20271_ _20261_/A _20390_/D _20260_/A vssd1 vssd1 vccd1 vccd1 _20398_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__19318__C _19322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16304__A _16304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12183__A2 _12123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22010_ _21908_/X _21911_/X _21915_/Y _21932_/Y _22024_/B vssd1 vssd1 vccd1 vccd1
+ _22086_/A sky130_fd_sc_hd__o221ai_4
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17119__B _21019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15657__B1 _16431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19615__A _19615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19334__B _19334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22912_ _22915_/CLK _22912_/D vssd1 vssd1 vccd1 vccd1 _22912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16621__A2 _16377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22843_ _22937_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _22843_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19350__A _19350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11614__C _15774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22774_ _22808_/CLK _22774_/D vssd1 vssd1 vccd1 vccd1 _22774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21725_ _21725_/A _21725_/B _22041_/B vssd1 vssd1 vccd1 vccd1 _21725_/Y sky130_fd_sc_hd__nand3_2
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11911__A _11911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22458__A1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21656_ _21654_/X _21642_/Y _21662_/A vssd1 vssd1 vccd1 vccd1 _21656_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12946__A1 _20249_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20607_ _20611_/B vssd1 vssd1 vccd1 vccd1 _20917_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11630__B _11647_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21587_ _21936_/A _13521_/B _21937_/A _21757_/D _21749_/A vssd1 vssd1 vccd1 vccd1
+ _21587_/Y sky130_fd_sc_hd__a32oi_2
XFILLER_138_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12445__C _15799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11340_ _11720_/A _11423_/A _11334_/X vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__a21bo_1
X_20538_ _20653_/A _20538_/B _20538_/C vssd1 vssd1 vccd1 vccd1 _20658_/A sky130_fd_sc_hd__nand3_2
XANTENNA__22861__D _22873_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11271_ _22784_/Q vssd1 vssd1 vccd1 vccd1 _11385_/C sky130_fd_sc_hd__buf_2
XFILLER_153_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20469_ _12734_/X _16611_/A _20343_/A _20464_/A vssd1 vssd1 vccd1 vccd1 _20469_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12742__A _12742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13010_ _13000_/X _13039_/A _13009_/Y vssd1 vssd1 vccd1 vccd1 _13011_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__17637__A1 _17730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22208_ _22208_/A _22208_/B vssd1 vssd1 vccd1 vccd1 _22211_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15648__B1 _15645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22139_ _22075_/X _22074_/Y _22079_/B vssd1 vssd1 vccd1 vccd1 _22140_/B sky130_fd_sc_hd__o21ai_1
XFILLER_121_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A wb_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ _14961_/A _14961_/B vssd1 vssd1 vccd1 vccd1 _14971_/C sky130_fd_sc_hd__nand2_1
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21493__C _21741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22394__A0 _16322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16700_ _16700_/A _16700_/B vssd1 vssd1 vccd1 vccd1 _22953_/D sky130_fd_sc_hd__xor2_4
XFILLER_48_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13912_ _13903_/Y _13937_/A _13911_/X vssd1 vssd1 vccd1 vccd1 _14021_/A sky130_fd_sc_hd__a21o_1
X_17680_ _17679_/B _17679_/C _17669_/X vssd1 vssd1 vccd1 vccd1 _17681_/B sky130_fd_sc_hd__a21bo_1
XFILLER_101_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14892_ _14892_/A _14955_/A _14892_/C _14892_/D vssd1 vssd1 vccd1 vccd1 _14955_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_63_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16631_ _16631_/A _16706_/A vssd1 vssd1 vccd1 vccd1 _16634_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16612__A2 _17435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13843_ _13963_/A _13963_/B _13892_/A _13963_/D vssd1 vssd1 vccd1 vccd1 _13849_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_75_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19350_ _19350_/A vssd1 vssd1 vccd1 vccd1 _19350_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16562_ _16751_/A vssd1 vssd1 vccd1 vccd1 _16599_/B sky130_fd_sc_hd__buf_2
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13774_ _13776_/B _14383_/A _13776_/A vssd1 vssd1 vccd1 vccd1 _14184_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13977__A3 _14911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18301_ _18572_/C _18301_/B _18301_/C vssd1 vssd1 vccd1 vccd1 _18309_/B sky130_fd_sc_hd__nand3b_1
XFILLER_188_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15513_ _15513_/A _15513_/B vssd1 vssd1 vccd1 vccd1 _15513_/Y sky130_fd_sc_hd__nand2_1
X_19281_ _19281_/A vssd1 vssd1 vccd1 vccd1 _19750_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12725_ _12602_/Y _12613_/Y _12584_/A _12630_/B _12601_/Y vssd1 vssd1 vccd1 vccd1
+ _12739_/C sky130_fd_sc_hd__o2111ai_4
X_16493_ _16493_/A _16493_/B vssd1 vssd1 vccd1 vccd1 _16493_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11821__A _16014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18232_ _18232_/A _18232_/B _18232_/C vssd1 vssd1 vccd1 vccd1 _18232_/X sky130_fd_sc_hd__and3_2
XFILLER_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15444_ _15804_/C vssd1 vssd1 vccd1 vccd1 _16106_/D sky130_fd_sc_hd__buf_2
XANTENNA__22449__A1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12656_ _22826_/Q vssd1 vssd1 vccd1 vccd1 _20390_/B sky130_fd_sc_hd__buf_2
XFILLER_31_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19314__A1 _16098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18163_ _18163_/A _18163_/B _18163_/C vssd1 vssd1 vccd1 vccd1 _18163_/Y sky130_fd_sc_hd__nand3_2
X_11607_ _22791_/Q vssd1 vssd1 vccd1 vccd1 _18115_/A sky130_fd_sc_hd__clkbuf_4
X_15375_ _15664_/A _15665_/A _15367_/X _15374_/X vssd1 vssd1 vccd1 vccd1 _15384_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_12587_ _15559_/C _15559_/D _12610_/A vssd1 vssd1 vccd1 vccd1 _12587_/Y sky130_fd_sc_hd__nand3_1
XFILLER_168_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18668__A3 _16276_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17114_ _17311_/A _17311_/B _17311_/C vssd1 vssd1 vccd1 vccd1 _17323_/A sky130_fd_sc_hd__nand3_2
XFILLER_172_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14326_ _12528_/A _14308_/X _14313_/X _13230_/X _14325_/X vssd1 vssd1 vccd1 vccd1
+ _14326_/X sky130_fd_sc_hd__a221o_1
XFILLER_183_250 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18094_ _18090_/Y _18091_/Y _18092_/Y _18093_/Y vssd1 vssd1 vccd1 vccd1 _18108_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_11538_ _11583_/B vssd1 vssd1 vccd1 vccd1 _18367_/C sky130_fd_sc_hd__buf_2
XANTENNA__19419__B _19419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17045_ _16880_/X _16879_/X _16885_/B vssd1 vssd1 vccd1 vccd1 _17045_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12074__D _12074_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15351__A2 _16300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14257_ _14256_/C _14256_/A _14256_/B vssd1 vssd1 vccd1 vccd1 _14281_/B sky130_fd_sc_hd__a21o_1
X_11469_ _18115_/C _11429_/A _11783_/C _11418_/A vssd1 vssd1 vccd1 vccd1 _11587_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16124__A _19336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13362__A1 _21964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ _13517_/C vssd1 vssd1 vccd1 vccd1 _21398_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14188_ _14188_/A _14188_/B _14188_/C vssd1 vssd1 vccd1 vccd1 _14198_/B sky130_fd_sc_hd__nand3_1
XFILLER_87_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1063 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ _13139_/A _13139_/B vssd1 vssd1 vccd1 vccd1 _13139_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17881__C _21019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18996_ _18996_/A vssd1 vssd1 vccd1 vccd1 _19179_/C sky130_fd_sc_hd__clkbuf_4
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12090__C _12090_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _18020_/B _18020_/A _17899_/B vssd1 vssd1 vccd1 vccd1 _17948_/B sky130_fd_sc_hd__o21a_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21456__A2_N _21866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19154__B _19614_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22385__A0 _12413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17878_ _19901_/D _17806_/D _17872_/X _17877_/X vssd1 vssd1 vccd1 vccd1 _17889_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_39_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16829_ _16845_/A _17189_/B _16986_/A _16986_/B vssd1 vssd1 vccd1 vccd1 _16906_/B
+ sky130_fd_sc_hd__nand4_1
X_19617_ _19772_/B vssd1 vssd1 vccd1 vccd1 _19985_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14614__B2 _14503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19548_ _19408_/X _19401_/X _19407_/X vssd1 vssd1 vccd1 vccd1 _19552_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19553__A1 _19455_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21850__D _22106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13930__B _13930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19479_ _19477_/X _19479_/B _19479_/C vssd1 vssd1 vccd1 vccd1 _19630_/C sky130_fd_sc_hd__nand3b_4
XFILLER_94_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21510_ _21386_/B _21509_/Y _21386_/A vssd1 vssd1 vccd1 vccd1 _21650_/C sky130_fd_sc_hd__a21boi_2
X_22490_ _22490_/A vssd1 vssd1 vccd1 vccd1 _22740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22951__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21441_ _21440_/Y _21415_/A _21423_/A _21559_/B vssd1 vssd1 vccd1 vccd1 _21576_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_194_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15590__A2 _12727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17316__B1 _17085_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15327__C1 _15776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21372_ _21372_/A _21372_/B _21372_/C vssd1 vssd1 vccd1 vccd1 _21372_/X sky130_fd_sc_hd__and3_1
XFILLER_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20323_ _20323_/A _20323_/B _20675_/C _20323_/D vssd1 vssd1 vccd1 vccd1 _20323_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_135_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15342__A2 _15341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19048__C _19199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20254_ _20241_/A _15450_/X _20249_/A vssd1 vssd1 vccd1 vccd1 _20262_/B sky130_fd_sc_hd__o21ai_4
XFILLER_192_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17095__A2 _17739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20185_ _20304_/B vssd1 vssd1 vccd1 vccd1 _20442_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22376__A0 _12470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14489__A _15006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11906__A _18305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17252__C1 _17401_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14066__C1 _14834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22856__D _22868_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22826_ _22850_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 _22826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22757_ _22757_/CLK _22757_/D vssd1 vssd1 vccd1 vccd1 _22757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ _12510_/A _12510_/B vssd1 vssd1 vccd1 vccd1 _12564_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13490_ _13556_/A _13554_/A vssd1 vssd1 vccd1 vccd1 _13496_/B sky130_fd_sc_hd__nand2_1
X_21708_ _21566_/A _21566_/B _21574_/A _21820_/A vssd1 vssd1 vccd1 vccd1 _21708_/X
+ sky130_fd_sc_hd__a22o_1
X_22688_ _22690_/CLK _22688_/D vssd1 vssd1 vccd1 vccd1 _22688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12441_ _15558_/C _20130_/B _12610_/A _12458_/A _20456_/C vssd1 vssd1 vccd1 vccd1
+ _12441_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21639_ _21449_/B _21629_/Y _21633_/Y _21631_/A vssd1 vssd1 vccd1 vccd1 _21640_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19847__A2 _19353_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15581__A2 _15546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15318__C1 _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15160_ _15160_/A _15160_/B vssd1 vssd1 vccd1 vccd1 _15161_/B sky130_fd_sc_hd__or2_1
X_12372_ _22817_/Q vssd1 vssd1 vccd1 vccd1 _12579_/C sky130_fd_sc_hd__buf_2
XFILLER_153_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17322__A3 _17122_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11323_ _11712_/A vssd1 vssd1 vccd1 vccd1 _11675_/A sky130_fd_sc_hd__clkbuf_2
X_14111_ _14112_/A _14963_/B _14210_/A _14113_/B vssd1 vssd1 vccd1 vccd1 _14111_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_153_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15091_ _15092_/A _15092_/B _15092_/C vssd1 vssd1 vccd1 vccd1 _15095_/A sky130_fd_sc_hd__a21o_1
XANTENNA__15333__A2 _12577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15486__C _15486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18807__B1 _19455_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14042_ _14042_/A vssd1 vssd1 vccd1 vccd1 _14561_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_140_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16879__A _16879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18797__C _18797_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18850_ _18850_/A vssd1 vssd1 vccd1 vccd1 _19013_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17801_ _18044_/A vssd1 vssd1 vccd1 vccd1 _18048_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__16598__B _16598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18781_ _18776_/Y _18779_/Y _18780_/X vssd1 vssd1 vccd1 vccd1 _19132_/C sky130_fd_sc_hd__o21ai_4
X_15993_ _15904_/X _15905_/X _20452_/A _20452_/B vssd1 vssd1 vccd1 vccd1 _15993_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12304__C1 _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17732_ _17732_/A vssd1 vssd1 vccd1 vccd1 _17733_/A sky130_fd_sc_hd__buf_2
XFILLER_85_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14944_ _14945_/A _15001_/A _14943_/X vssd1 vssd1 vccd1 vccd1 _14947_/C sky130_fd_sc_hd__a21o_1
XANTENNA__22824__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17663_ _17663_/A _17663_/B vssd1 vssd1 vccd1 vccd1 _17663_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14875_ _14685_/B _14862_/A _14884_/C vssd1 vssd1 vccd1 vccd1 _14880_/A sky130_fd_sc_hd__o21ai_2
XFILLER_75_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16597__B2 _16598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19402_ _19407_/A _19408_/A _19401_/X vssd1 vssd1 vccd1 vccd1 _19410_/A sky130_fd_sc_hd__a21o_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16614_ _16609_/X _16613_/X _16354_/C vssd1 vssd1 vccd1 vccd1 _16617_/D sky130_fd_sc_hd__o21ai_4
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13826_ _13826_/A _13826_/B _13826_/C vssd1 vssd1 vccd1 vccd1 _14069_/C sky130_fd_sc_hd__nand3_4
XFILLER_91_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17594_ _17624_/B _17624_/A _17625_/A vssd1 vssd1 vccd1 vccd1 _17597_/C sky130_fd_sc_hd__nand3b_1
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19333_ _19687_/A vssd1 vssd1 vccd1 vccd1 _19842_/A sky130_fd_sc_hd__buf_2
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16545_ _16512_/A _16512_/B _16542_/Y _16544_/Y vssd1 vssd1 vccd1 vccd1 _16545_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__12069__D _19046_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13757_ _22754_/Q vssd1 vssd1 vccd1 vccd1 _13766_/A sky130_fd_sc_hd__inv_2
XFILLER_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17546__B1 _17423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21342__B2 _21341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15023__A _15213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17010__A2 _16836_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19264_ _19272_/B vssd1 vssd1 vccd1 vccd1 _19434_/A sky130_fd_sc_hd__clkbuf_2
X_12708_ _12708_/A vssd1 vssd1 vccd1 vccd1 _12950_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16476_ _16476_/A vssd1 vssd1 vccd1 vccd1 _16476_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20696__A3 _13016_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13688_ _21294_/B _22672_/Q vssd1 vssd1 vccd1 vccd1 _13689_/B sky130_fd_sc_hd__nand2_1
X_18215_ _12188_/A _12188_/B _12188_/C _18227_/C vssd1 vssd1 vccd1 vccd1 _18215_/Y
+ sky130_fd_sc_hd__a31oi_2
X_15427_ _15797_/A vssd1 vssd1 vccd1 vccd1 _15427_/X sky130_fd_sc_hd__buf_4
XFILLER_31_587 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19195_ _11786_/X _15839_/A _19059_/Y vssd1 vssd1 vccd1 vccd1 _19195_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_54_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12639_ _12640_/A _12640_/B _12742_/A vssd1 vssd1 vccd1 vccd1 _12668_/A sky130_fd_sc_hd__a21o_1
XFILLER_141_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16780__C _17246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18146_ _18146_/A _18146_/B _18146_/C vssd1 vssd1 vccd1 vccd1 _18172_/A sky130_fd_sc_hd__nand3_2
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ _15377_/A vssd1 vssd1 vccd1 vccd1 _15358_/X sky130_fd_sc_hd__buf_4
XANTENNA__20302__C1 _20314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14309_ input26/X vssd1 vssd1 vccd1 vccd1 _22514_/A sky130_fd_sc_hd__clkbuf_1
X_18077_ _18077_/A vssd1 vssd1 vccd1 vccd1 _18077_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12382__A _22821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15289_ _15288_/A _15271_/B _22884_/Q vssd1 vssd1 vccd1 vccd1 _15290_/B sky130_fd_sc_hd__a21oi_1
XFILLER_172_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17028_ _17028_/A _17028_/B _17028_/C vssd1 vssd1 vccd1 vccd1 _17036_/B sky130_fd_sc_hd__nand3_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13197__B _21494_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20081__A1 _20728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18979_ _18895_/X _19022_/C _19009_/A vssd1 vssd1 vccd1 vccd1 _19085_/B sky130_fd_sc_hd__o21ai_2
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21990_ _21990_/A _21990_/B _21990_/C vssd1 vssd1 vccd1 vccd1 _21990_/X sky130_fd_sc_hd__and3_1
XFILLER_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20941_ _20941_/A _20941_/B _20941_/C vssd1 vssd1 vccd1 vccd1 _20945_/A sky130_fd_sc_hd__nand3_1
XFILLER_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18982__C1 _17313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20872_ _17816_/A _20806_/B _20871_/Y _20788_/B vssd1 vssd1 vccd1 vccd1 _20876_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22611_ _18127_/B input36/X _22619_/S vssd1 vssd1 vccd1 vccd1 _22612_/A sky130_fd_sc_hd__mux2_1
XANTENNA__22530__A0 _13799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20136__A2 _20126_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11461__A _12090_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22542_ _22542_/A vssd1 vssd1 vccd1 vccd1 _22763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15868__A _17385_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22473_ _21580_/B input39/X _22475_/S vssd1 vssd1 vccd1 vccd1 _22474_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12707__D _20576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15563__A2 _16274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14772__A _22766_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18244__A _18259_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21424_ _21424_/A _21559_/A _21424_/C vssd1 vssd1 vccd1 vccd1 _21426_/B sky130_fd_sc_hd__nand3_1
XFILLER_135_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21355_ _21387_/A _21387_/B _21355_/C vssd1 vssd1 vccd1 vccd1 _21393_/A sky130_fd_sc_hd__nand3_2
XANTENNA__15315__A2 _16932_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20306_ _20304_/Y _20195_/Y _20305_/X vssd1 vssd1 vccd1 vccd1 _20432_/B sky130_fd_sc_hd__o21ai_4
XFILLER_190_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21286_ _21700_/A _21701_/A vssd1 vssd1 vccd1 vccd1 _21558_/A sky130_fd_sc_hd__nor2_1
XFILLER_146_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22597__A0 _11349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18265__A1 _18088_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20237_ _20678_/B _20579_/C _20219_/Y _20085_/X vssd1 vssd1 vccd1 vccd1 _20237_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22847__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15079__A1 _13851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20072__A1 _12522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16815__A2 _15960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20168_ _12875_/X _12879_/Y _12868_/X vssd1 vssd1 vccd1 vccd1 _20169_/B sky130_fd_sc_hd__o21ai_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_67 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20099_ _20486_/C _16261_/B _20096_/Y _20098_/Y vssd1 vssd1 vccd1 vccd1 _20119_/C
+ sky130_fd_sc_hd__a22o_2
X_12990_ _12990_/A _12990_/B _13036_/A _12990_/D vssd1 vssd1 vccd1 vccd1 _13031_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _11941_/A vssd1 vssd1 vccd1 vccd1 _18107_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21572__A1 _22674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13851__A _13851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14660_ _14758_/C _14660_/B vssd1 vssd1 vccd1 vccd1 _14664_/A sky130_fd_sc_hd__xnor2_2
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11868_/Y _11869_/X _11871_/X vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__a21boi_1
XFILLER_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15251__A1 _15180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13611_ _13611_/A _13611_/B _13611_/C vssd1 vssd1 vccd1 vccd1 _13612_/B sky130_fd_sc_hd__nand3_1
XFILLER_38_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22809_ _22810_/CLK _22809_/D vssd1 vssd1 vccd1 vccd1 _22809_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22521__A0 _13761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14591_ _13737_/X _13746_/X _13923_/X vssd1 vssd1 vccd1 vccd1 _14591_/X sky130_fd_sc_hd__a21o_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12467__A _12467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16330_ _16579_/A _16580_/A _20357_/A vssd1 vssd1 vccd1 vccd1 _16331_/A sky130_fd_sc_hd__o21ai_2
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13542_ _13533_/Y _13534_/Y _13471_/Y _13473_/X _13537_/B vssd1 vssd1 vccd1 vccd1
+ _13543_/C sky130_fd_sc_hd__o221ai_1
XFILLER_186_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16261_ _19322_/A _16261_/B _17280_/A _17246_/A vssd1 vssd1 vccd1 vccd1 _16261_/Y
+ sky130_fd_sc_hd__nand4_4
XANTENNA__15554__A2 _19687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13473_ _13447_/X _13169_/X _13446_/X _13563_/B _13454_/B vssd1 vssd1 vccd1 vccd1
+ _13473_/X sky130_fd_sc_hd__a32o_1
XFILLER_13_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11521__D _18875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18000_ _17950_/A _17950_/B _17999_/Y _18002_/A vssd1 vssd1 vccd1 vccd1 _18048_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_185_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15212_ _15212_/A vssd1 vssd1 vccd1 vccd1 _15224_/A sky130_fd_sc_hd__clkbuf_2
X_12424_ _12437_/A _12904_/A _12424_/C vssd1 vssd1 vccd1 vccd1 _12424_/Y sky130_fd_sc_hd__nand3_4
X_16192_ _20734_/A _16192_/B _17401_/A _16192_/D vssd1 vssd1 vccd1 vccd1 _16192_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_154_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15143_ _15175_/B _15143_/B vssd1 vssd1 vccd1 vccd1 _22681_/D sky130_fd_sc_hd__xor2_1
X_12355_ _12401_/A _12284_/A _15631_/C _12377_/A vssd1 vssd1 vccd1 vccd1 _12813_/A
+ sky130_fd_sc_hd__a31o_2
XANTENNA__14109__A3 _15115_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21011__C _21011_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11306_ _11306_/A vssd1 vssd1 vccd1 vccd1 _11306_/X sky130_fd_sc_hd__buf_4
X_19951_ _20037_/C _19951_/B vssd1 vssd1 vccd1 vccd1 _19991_/B sky130_fd_sc_hd__or2_1
XFILLER_153_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15074_ _15074_/A _15074_/B _15074_/C vssd1 vssd1 vccd1 vccd1 _15128_/B sky130_fd_sc_hd__or3_1
X_12286_ _12368_/D vssd1 vssd1 vccd1 vccd1 _12413_/A sky130_fd_sc_hd__buf_2
XFILLER_141_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22404__A _22426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__A1_N _11897_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18902_ _19085_/A _19009_/A _18895_/X _19022_/C vssd1 vssd1 vccd1 vccd1 _18907_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_113_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14025_ _13862_/A _14014_/X _14061_/D _14024_/Y vssd1 vssd1 vccd1 vccd1 _14044_/C
+ sky130_fd_sc_hd__o211ai_4
X_19882_ _19881_/A _19881_/B _19881_/C vssd1 vssd1 vccd1 vccd1 _19882_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12930__A _12930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18833_ _18633_/Y _18619_/Y _18835_/A vssd1 vssd1 vccd1 vccd1 _18833_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_1_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11546__A _11644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19205__B1 _18629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18764_ _18764_/A _18764_/B vssd1 vssd1 vccd1 vccd1 _18768_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15976_ _15976_/A _15976_/B _15976_/C vssd1 vssd1 vccd1 vccd1 _16010_/A sky130_fd_sc_hd__nand3_2
XFILLER_64_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21012__B1 _12671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17715_ _17721_/C _17721_/A _22900_/Q vssd1 vssd1 vccd1 vccd1 _17716_/B sky130_fd_sc_hd__and3_1
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14927_ _14927_/A _14927_/B vssd1 vssd1 vccd1 vccd1 _14929_/C sky130_fd_sc_hd__xor2_4
XFILLER_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18695_ _18695_/A vssd1 vssd1 vccd1 vccd1 _18695_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14832__A4 _15186_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14857__A _14857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17646_ _17646_/A vssd1 vssd1 vccd1 vccd1 _19689_/C sky130_fd_sc_hd__buf_2
X_14858_ _14858_/A vssd1 vssd1 vccd1 vccd1 _15050_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14045__A2 _14273_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19508__A1 _19346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13809_ _22756_/Q vssd1 vssd1 vccd1 vccd1 _13826_/C sky130_fd_sc_hd__buf_2
X_17577_ _17628_/A _17580_/A _17578_/A vssd1 vssd1 vccd1 vccd1 _17579_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13253__B1 _21629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16990__A1 _16822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15793__A2 _15834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14789_ _14576_/X _15240_/C _14788_/Y vssd1 vssd1 vccd1 vccd1 _14884_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__14596__A3 _14942_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19316_ _19316_/A _19316_/B vssd1 vssd1 vccd1 vccd1 _19317_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11281__A _22799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16528_ _16526_/X _16527_/X _16493_/Y _16502_/Y vssd1 vssd1 vccd1 vccd1 _16529_/C
+ sky130_fd_sc_hd__o22ai_1
XFILLER_91_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11712__C _11712_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19247_ _19244_/Y _19245_/Y _19246_/Y vssd1 vssd1 vccd1 vccd1 _19248_/B sky130_fd_sc_hd__o21ai_1
XFILLER_104_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16459_ _15589_/X _16474_/A _16455_/X _16458_/Y vssd1 vssd1 vccd1 vccd1 _16463_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_177_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19178_ _19016_/Y _19167_/Y _18849_/D _19334_/A _19687_/A vssd1 vssd1 vccd1 vccd1
+ _19179_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_157_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11567__B1 _11565_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18129_ _18129_/A _18129_/B vssd1 vssd1 vccd1 vccd1 _19587_/D sky130_fd_sc_hd__nand2_4
XANTENNA__19692__B1 _19461_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22028__C1 _21220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21140_ _21141_/A _21141_/B _22944_/Q vssd1 vssd1 vccd1 vccd1 _21142_/A sky130_fd_sc_hd__o21ba_1
XFILLER_172_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21071_ _21037_/D _21079_/A _21079_/B vssd1 vssd1 vccd1 vccd1 _21071_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_160_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20022_ _20022_/A _20022_/B vssd1 vssd1 vccd1 vccd1 _20024_/C sky130_fd_sc_hd__or2_1
XANTENNA__18798__A2 _16940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16695__A_N _22890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_602 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15870__B _20806_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21973_ _22182_/B _22176_/A _21964_/X _21606_/X vssd1 vssd1 vccd1 vccd1 _21973_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20924_ _20922_/X _20936_/D _12928_/X _17922_/A vssd1 vssd1 vccd1 vccd1 _20924_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__19061__C _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16430__B1 _16400_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12047__A1 _22658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _20514_/X _17435_/A _20780_/Y vssd1 vssd1 vccd1 vccd1 _20855_/Y sky130_fd_sc_hd__o21ai_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12287__A _22703_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20109__A2 _16715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20786_ _20210_/B _20680_/X _20787_/B _20787_/C vssd1 vssd1 vccd1 vccd1 _20788_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_195_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22525_ _13826_/C input61/X _22525_/S vssd1 vssd1 vccd1 vccd1 _22526_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16733__A1 _16723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17930__B1 _17928_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22456_ _13131_/X input62/X _22464_/S vssd1 vssd1 vccd1 vccd1 _22457_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21407_ _21390_/Y _21394_/Y _21401_/Y vssd1 vssd1 vccd1 vccd1 _21410_/A sky130_fd_sc_hd__a21bo_1
X_22387_ _12320_/A input64/X _22391_/S vssd1 vssd1 vccd1 vccd1 _22388_/A sky130_fd_sc_hd__mux2_1
XANTENNA__21085__A3 _17839_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12140_ _11977_/Y _11970_/Y _12137_/A vssd1 vssd1 vccd1 vccd1 _12143_/A sky130_fd_sc_hd__a21boi_1
XFILLER_191_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21338_ _21338_/A _21338_/B vssd1 vssd1 vccd1 vccd1 _21454_/A sky130_fd_sc_hd__nand2_1
XFILLER_151_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12071_ _18830_/A _18305_/B _16192_/D _16157_/D vssd1 vssd1 vccd1 vccd1 _12074_/C
+ sky130_fd_sc_hd__and4_1
X_21269_ _21269_/A vssd1 vssd1 vccd1 vccd1 _21841_/A sky130_fd_sc_hd__buf_2
XANTENNA__14511__A3 _14834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _15978_/C vssd1 vssd1 vccd1 vccd1 _16613_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_106_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17461__A2 _17981_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _15761_/A _15761_/B _15761_/C vssd1 vssd1 vccd1 vccd1 _16402_/A sky130_fd_sc_hd__nand3_1
XFILLER_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12973_ _12973_/A vssd1 vssd1 vccd1 vccd1 _20792_/C sky130_fd_sc_hd__buf_2
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17749__B1 _17880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17500_ _17507_/A _18044_/A _17853_/A vssd1 vssd1 vccd1 vccd1 _17500_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _14712_/A _14712_/B vssd1 vssd1 vccd1 vccd1 _14712_/Y sky130_fd_sc_hd__nor2_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _18376_/Y _18396_/C _18559_/A vssd1 vssd1 vccd1 vccd1 _18556_/A sky130_fd_sc_hd__a21boi_4
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11924_ _12077_/D _12077_/C _11924_/C _11924_/D vssd1 vssd1 vccd1 vccd1 _11924_/X
+ sky130_fd_sc_hd__and4_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _11935_/B _12930_/A _15302_/A _15691_/Y vssd1 vssd1 vccd1 vccd1 _15693_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _19615_/C _17431_/B _17431_/C _17431_/D vssd1 vssd1 vccd1 vccd1 _17433_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _14669_/A _14057_/X _14642_/Y vssd1 vssd1 vccd1 vccd1 _14646_/B sky130_fd_sc_hd__o21ai_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _18706_/A vssd1 vssd1 vccd1 vccd1 _15991_/D sky130_fd_sc_hd__buf_4
XFILLER_61_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output105_A _14426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17362_ _17373_/A vssd1 vssd1 vccd1 vccd1 _17959_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11532__C _18093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14574_ _14688_/A vssd1 vssd1 vccd1 vccd1 _15010_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11786_ _12010_/A vssd1 vssd1 vccd1 vccd1 _11786_/X sky130_fd_sc_hd__buf_4
X_19101_ _18914_/A _18914_/B _18914_/C _18931_/B _18977_/B vssd1 vssd1 vccd1 vccd1
+ _19257_/A sky130_fd_sc_hd__a32oi_4
XFILLER_13_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16313_ _20092_/A _20092_/B _16313_/C vssd1 vssd1 vccd1 vccd1 _16313_/X sky130_fd_sc_hd__and3_1
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ _13350_/A _13633_/B _13633_/C _13506_/C _13506_/B vssd1 vssd1 vccd1 vccd1
+ _13526_/B sky130_fd_sc_hd__o32a_1
XFILLER_41_682 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17293_ _17293_/A _17293_/B vssd1 vssd1 vccd1 vccd1 _17293_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17382__D1 _18197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19032_ _19037_/A _19037_/B _19031_/X vssd1 vssd1 vccd1 vccd1 _19032_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_51_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14843__C _14843_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16244_ _16498_/C vssd1 vssd1 vccd1 vccd1 _19507_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__15301__A _16257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ _13456_/A vssd1 vssd1 vccd1 vccd1 _21621_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11549__B1 _11895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20808__B1 _20178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18477__A1 _18765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12407_ _12407_/A _12407_/B vssd1 vssd1 vccd1 vccd1 _12432_/A sky130_fd_sc_hd__nand2_1
X_16175_ _16143_/Y _16173_/Y _16118_/C _16174_/X vssd1 vssd1 vccd1 vccd1 _16175_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_13387_ _21249_/B _13390_/B vssd1 vssd1 vccd1 vccd1 _13387_/X sky130_fd_sc_hd__xor2_1
XFILLER_126_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput107 _14333_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[3] sky130_fd_sc_hd__buf_2
Xoutput118 _22666_/Q vssd1 vssd1 vccd1 vccd1 y[2] sky130_fd_sc_hd__buf_2
XFILLER_127_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15126_ _15122_/X _15124_/Y _15118_/C vssd1 vssd1 vccd1 vccd1 _15128_/D sky130_fd_sc_hd__o21ai_1
XFILLER_154_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338_ _22696_/Q vssd1 vssd1 vccd1 vccd1 _12361_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13756__A _22858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19934_ _19971_/B _19934_/B vssd1 vssd1 vccd1 vccd1 _19935_/A sky130_fd_sc_hd__and2_1
X_15057_ _15057_/A vssd1 vssd1 vccd1 vccd1 _15185_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12660__A _15586_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ _22692_/Q vssd1 vssd1 vccd1 vccd1 _12396_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14008_ _13916_/Y _14021_/C _13886_/Y _13879_/X vssd1 vssd1 vccd1 vccd1 _14033_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__13475__B _13475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19865_ _19865_/A _19865_/B vssd1 vssd1 vccd1 vccd1 _19866_/B sky130_fd_sc_hd__nand2_1
XFILLER_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19443__A _19443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18816_ _18825_/A _19079_/A _18818_/A _18818_/B vssd1 vssd1 vccd1 vccd1 _18823_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18985__C _18985_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19796_ _19796_/A _19796_/B _19796_/C vssd1 vssd1 vccd1 vccd1 _19796_/X sky130_fd_sc_hd__and3_1
XANTENNA__15463__A1 _15755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18747_ _18646_/B _18746_/Y _18645_/Y vssd1 vssd1 vccd1 vccd1 _18748_/B sky130_fd_sc_hd__a21oi_2
X_15959_ _15959_/A _16400_/C _17816_/A vssd1 vssd1 vccd1 vccd1 _15959_/X sky130_fd_sc_hd__and3_2
XFILLER_49_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14671__C1 _15213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18678_ _18319_/A _18678_/B _18678_/C _18678_/D vssd1 vssd1 vccd1 vccd1 _18841_/A
+ sky130_fd_sc_hd__nand4b_2
XANTENNA__20101__B _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17629_ _17627_/X _17581_/B _17580_/Y vssd1 vssd1 vccd1 vccd1 _17629_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13226__B1 _13340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17113__D _17530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20640_ _20631_/Y _20737_/A _20638_/Y _20639_/X vssd1 vssd1 vccd1 vccd1 _20640_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__22954__D _22954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20571_ _15325_/X _15326_/X _20723_/A _17401_/A _20745_/A vssd1 vssd1 vccd1 vccd1
+ _20575_/B sky130_fd_sc_hd__o2111ai_4
XANTENNA__16307__A _20605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22310_ _22310_/A _22310_/B vssd1 vssd1 vccd1 vccd1 _22310_/X sky130_fd_sc_hd__and2_1
XFILLER_164_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22241_ _22241_/A _22241_/B vssd1 vssd1 vccd1 vccd1 _22243_/A sky130_fd_sc_hd__or2_1
XFILLER_180_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20275__A1 _20143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22172_ _22172_/A vssd1 vssd1 vccd1 vccd1 _22304_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11960__B1 _11935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21123_ _21072_/Y _21065_/X _21071_/Y _21104_/B vssd1 vssd1 vccd1 vccd1 _21130_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__15151__B1 _15182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21054_ _21054_/A _21054_/B vssd1 vssd1 vccd1 vccd1 _21055_/B sky130_fd_sc_hd__xnor2_1
XFILLER_99_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20578__A2 _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20005_ _20005_/A _20026_/B _20024_/B vssd1 vssd1 vccd1 vccd1 _20008_/A sky130_fd_sc_hd__and3_1
XFILLER_143_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16651__B1 _16431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19196__A2 _17635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21956_ _22042_/A vssd1 vssd1 vccd1 vccd1 _22037_/C sky130_fd_sc_hd__clkbuf_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _20907_/A vssd1 vssd1 vccd1 vccd1 _21037_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21887_ _21891_/A _21891_/B _21892_/B _21892_/C vssd1 vssd1 vccd1 vccd1 _21889_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12448__C _16256_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11640_ _11504_/X _11505_/X _11626_/X _11625_/X _11779_/B vssd1 vssd1 vccd1 vccd1
+ _11745_/B sky130_fd_sc_hd__o221a_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22864__D _22876_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20838_ _20902_/A _20833_/Y _20837_/Y vssd1 vssd1 vccd1 vccd1 _20839_/B sky130_fd_sc_hd__a21oi_1
XFILLER_74_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11571_ _19465_/A vssd1 vssd1 vccd1 vccd1 _19619_/B sky130_fd_sc_hd__buf_4
XFILLER_11_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20769_ _20566_/Y _20565_/Y _20768_/Y _20667_/Y vssd1 vssd1 vccd1 vccd1 _20772_/D
+ sky130_fd_sc_hd__o211ai_2
XFILLER_195_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _13300_/Y _13309_/Y _13577_/A _21220_/A vssd1 vssd1 vccd1 vccd1 _13314_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_161_1087 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22508_ _22749_/Q input56/X _22508_/S vssd1 vssd1 vccd1 vccd1 _22509_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14290_ _14288_/A _14288_/B _14288_/C vssd1 vssd1 vccd1 vccd1 _14290_/X sky130_fd_sc_hd__a21o_1
XFILLER_168_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13241_ _22847_/Q vssd1 vssd1 vccd1 vccd1 _13421_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22439_ _22719_/Q input59/X _22439_/S vssd1 vssd1 vccd1 vccd1 _22440_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18432__A _18432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13172_ _21448_/C _21588_/B vssd1 vssd1 vccd1 vccd1 _13172_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_input66_A wb_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11951__B1 _15714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ _18208_/A _12123_/B _12123_/C vssd1 vssd1 vccd1 vccd1 _12184_/A sky130_fd_sc_hd__nand3_1
X_17980_ _19941_/B vssd1 vssd1 vccd1 vccd1 _19983_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_124_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16931_ _16988_/A _16988_/B vssd1 vssd1 vccd1 vccd1 _16982_/A sky130_fd_sc_hd__nand2_1
X_12054_ _12054_/A _12054_/B _12055_/A _12055_/B vssd1 vssd1 vccd1 vccd1 _12054_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11703__B1 _11702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20569__A2 _20511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15791__A _20359_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19650_ _19650_/A _19650_/B _19650_/C _19650_/D vssd1 vssd1 vccd1 vccd1 _19656_/B
+ sky130_fd_sc_hd__nand4_1
X_16862_ _16531_/Y _16536_/Y _16861_/Y _16624_/B _16619_/C vssd1 vssd1 vccd1 vccd1
+ _16867_/A sky130_fd_sc_hd__a32oi_1
XANTENNA__18631__A1 _18810_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18092__C1 _12003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18631__B2 _18459_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_719 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18601_ _18601_/A _18601_/B vssd1 vssd1 vccd1 vccd1 _18601_/Y sky130_fd_sc_hd__nand2_1
X_15813_ _15631_/A _12493_/Y _15899_/B _11506_/A _11779_/C vssd1 vssd1 vccd1 vccd1
+ _15813_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19581_ _19581_/A vssd1 vssd1 vccd1 vccd1 _19581_/Y sky130_fd_sc_hd__inv_2
X_16793_ _16782_/X _16781_/Y _16787_/Y _16788_/X vssd1 vssd1 vccd1 vccd1 _16803_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15996__A2 _15546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18532_ _18665_/A vssd1 vssd1 vccd1 vccd1 _19194_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15744_ _15457_/A _15696_/Y _15304_/B vssd1 vssd1 vccd1 vccd1 _15744_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12956_ _12957_/B _12957_/C _12957_/A vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__a21o_1
XANTENNA__21017__B _21017_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_908 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _18365_/Y _18366_/Y _18367_/Y _18368_/Y vssd1 vssd1 vccd1 vccd1 _18463_/X
+ sky130_fd_sc_hd__o211a_1
X_11907_ _11904_/X _11905_/X _18953_/C vssd1 vssd1 vccd1 vccd1 _11907_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15675_ _15510_/B _15672_/Y _15678_/A _15677_/B _15677_/C vssd1 vssd1 vccd1 vccd1
+ _15676_/D sky130_fd_sc_hd__o2111ai_2
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16945__A1 _16940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ _12878_/X _12776_/X _16160_/C _20870_/C vssd1 vssd1 vccd1 vccd1 _12887_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__16945__B2 _16944_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20741__A2 _20730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17414_ _15941_/A _17388_/X _17235_/Y _17383_/Y _17412_/X vssd1 vssd1 vccd1 vccd1
+ _17414_/X sky130_fd_sc_hd__o311a_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14626_/A _14626_/B vssd1 vssd1 vccd1 vccd1 _14626_/Y sky130_fd_sc_hd__nand2_1
X_18394_ _18377_/Y _18396_/C _18385_/Y _18393_/Y vssd1 vssd1 vccd1 vccd1 _18394_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11838_ _11838_/A _12246_/A _12246_/B vssd1 vssd1 vccd1 vccd1 _11838_/Y sky130_fd_sc_hd__nand3_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14420__A2 _14418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17345_ _17341_/X _17338_/X _17337_/X vssd1 vssd1 vccd1 vccd1 _17345_/X sky130_fd_sc_hd__o21a_1
XANTENNA__20575__C _20637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14843_/A _14843_/B _14552_/X vssd1 vssd1 vccd1 vccd1 _14665_/A sky130_fd_sc_hd__a21o_1
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11769_ _11995_/A vssd1 vssd1 vccd1 vccd1 _11783_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_996 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ _22041_/B vssd1 vssd1 vccd1 vccd1 _22108_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_159_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17276_ _16944_/Y _17129_/Y _17131_/Y vssd1 vssd1 vccd1 vccd1 _17288_/B sky130_fd_sc_hd__o21ai_2
XFILLER_158_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14488_ _14684_/C vssd1 vssd1 vccd1 vccd1 _15006_/C sky130_fd_sc_hd__buf_2
XFILLER_173_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19015_ _14431_/A _15808_/A _15690_/X _19490_/C _19490_/D vssd1 vssd1 vccd1 vccd1
+ _19015_/Y sky130_fd_sc_hd__o2111ai_4
X_16227_ _16227_/A vssd1 vssd1 vccd1 vccd1 _16227_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_bq_clk_i clkbuf_3_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_bq_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15966__A _17643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13439_ _13434_/X _13436_/Y _13437_/X _13438_/Y vssd1 vssd1 vccd1 vccd1 _13440_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__21049__A3 _17839_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13931__A1 _14765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16158_ _17085_/C vssd1 vssd1 vccd1 vccd1 _16997_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_127_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15109_ _15149_/A _15152_/A _15073_/A _15073_/C _15108_/Y vssd1 vssd1 vccd1 vccd1
+ _15111_/A sky130_fd_sc_hd__a221oi_1
XANTENNA__13486__A _13659_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_1094 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16089_ _15917_/X _16026_/A _16030_/Y _16088_/X vssd1 vssd1 vccd1 vccd1 _16090_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_115_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16881__B1 _16879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19917_ _19917_/A _19917_/B vssd1 vssd1 vccd1 vccd1 _19922_/B sky130_fd_sc_hd__xor2_2
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_844 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17108__D _17672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19173__A _19320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17425__A2 _17422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19848_ _19848_/A _19848_/B vssd1 vssd1 vccd1 vccd1 _19850_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19779_ _19782_/A _19782_/B _19837_/A _19787_/A vssd1 vssd1 vccd1 vccd1 _19785_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_56_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19178__A2 _19167_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__A _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21810_ _21814_/A _21814_/D vssd1 vssd1 vccd1 vccd1 _21810_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22790_ _22791_/CLK _22790_/D vssd1 vssd1 vccd1 vccd1 _22790_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18386__B1 _18387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12549__B _15363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21741_ _22041_/A _21741_/B _22041_/C vssd1 vssd1 vccd1 vccd1 _21742_/B sky130_fd_sc_hd__nand3_2
XFILLER_24_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20732__A2 _20730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_446 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17421__A _17421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21672_ _21648_/X _21657_/Y _21664_/X _21671_/Y vssd1 vssd1 vccd1 vccd1 _21676_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20623_ _20623_/A _20623_/B vssd1 vssd1 vccd1 vccd1 _20623_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20554_ _20554_/A _20554_/B _20554_/C _20554_/D vssd1 vssd1 vccd1 vccd1 _20554_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_165_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20485_ _20465_/X _20470_/Y _20499_/D _20484_/Y vssd1 vssd1 vccd1 vccd1 _20485_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_118_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13099__C _14380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_498 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22224_ _22304_/A _22262_/A _22304_/C _22221_/C vssd1 vssd1 vccd1 vccd1 _22224_/Y
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__18846__D1 _19358_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22155_ _22155_/A vssd1 vssd1 vccd1 vccd1 _22336_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21106_ _21106_/A _21106_/B vssd1 vssd1 vccd1 vccd1 _22922_/D sky130_fd_sc_hd__xnor2_1
XFILLER_160_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22086_ _22086_/A _22086_/B vssd1 vssd1 vccd1 vccd1 _22145_/B sky130_fd_sc_hd__nand2_1
XFILLER_120_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21037_ _21037_/A _21067_/B _21067_/C _21037_/D vssd1 vssd1 vccd1 vccd1 _21039_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_847 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17315__B _17520_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19169__A2 _12167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20971__A2 _15355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12810_ _12810_/A _12810_/B _12810_/C vssd1 vssd1 vccd1 vccd1 _12852_/A sky130_fd_sc_hd__nand3_1
XFILLER_90_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11644__A _11644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13790_ _22874_/Q vssd1 vssd1 vccd1 vccd1 _14044_/B sky130_fd_sc_hd__buf_2
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12741_ _12741_/A _12741_/B _12741_/C vssd1 vssd1 vccd1 vccd1 _13007_/C sky130_fd_sc_hd__nand3_2
X_21939_ _21939_/A _21939_/B vssd1 vssd1 vccd1 vccd1 _21952_/C sky130_fd_sc_hd__nand2_1
XFILLER_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _15810_/A _15810_/B _15991_/B vssd1 vssd1 vccd1 vccd1 _15461_/B sky130_fd_sc_hd__and3_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12672_/A vssd1 vssd1 vccd1 vccd1 _12719_/A sky130_fd_sc_hd__buf_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_788 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14402__A2 _14370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14411_/A vssd1 vssd1 vccd1 vccd1 _14411_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11745_/A vssd1 vssd1 vccd1 vccd1 _11623_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15391_ _15665_/B _15665_/C vssd1 vssd1 vccd1 vccd1 _15392_/C sky130_fd_sc_hd__nand2_1
XFILLER_23_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_630 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17130_ _16039_/A _17634_/A _17129_/Y vssd1 vssd1 vccd1 vccd1 _17134_/A sky130_fd_sc_hd__o21ai_1
XFILLER_128_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14342_ _11980_/C _14338_/X _14339_/X _14331_/X _12413_/X vssd1 vssd1 vccd1 vccd1
+ _14342_/X sky130_fd_sc_hd__a32o_1
XFILLER_129_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11554_ _11554_/A _11554_/B _11554_/C vssd1 vssd1 vccd1 vccd1 _11839_/A sky130_fd_sc_hd__nand3_1
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17061_ _16652_/A _16652_/B _16644_/Y _16645_/X _16889_/C vssd1 vssd1 vccd1 vccd1
+ _17061_/X sky130_fd_sc_hd__a41o_1
XFILLER_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14273_ _14273_/A _14575_/B _14273_/C vssd1 vssd1 vccd1 vccd1 _14276_/B sky130_fd_sc_hd__and3_1
XFILLER_155_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11485_ _18115_/D _11980_/A _11980_/B vssd1 vssd1 vccd1 vccd1 _12157_/A sky130_fd_sc_hd__nand3b_1
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1111 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _16012_/A _16012_/B vssd1 vssd1 vccd1 vccd1 _16012_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13224_ _13504_/A vssd1 vssd1 vccd1 vccd1 _21383_/A sky130_fd_sc_hd__buf_2
XFILLER_183_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11819__A _11819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17655__A2 _19768_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16458__A3 _12938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ _22845_/Q vssd1 vssd1 vccd1 vccd1 _21351_/C sky130_fd_sc_hd__buf_2
XFILLER_112_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _18099_/A _18319_/B vssd1 vssd1 vccd1 vccd1 _12107_/B sky130_fd_sc_hd__nand2_1
X_17963_ _17226_/X _17227_/X _17959_/A _17959_/B vssd1 vssd1 vccd1 vccd1 _17963_/X
+ sky130_fd_sc_hd__o211a_1
X_13086_ _21213_/A _21312_/B _21214_/A vssd1 vssd1 vccd1 vccd1 _13087_/A sky130_fd_sc_hd__nand3_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19702_ _19899_/A _17388_/X _19697_/D _19697_/B vssd1 vssd1 vccd1 vccd1 _19703_/C
+ sky130_fd_sc_hd__o211ai_1
X_16914_ _16293_/X _16294_/X _15690_/X _11666_/X _20608_/B vssd1 vssd1 vccd1 vccd1
+ _16914_/Y sky130_fd_sc_hd__o2111ai_4
X_12037_ _12034_/Y _11815_/Y _12035_/Y _12036_/Y vssd1 vssd1 vccd1 vccd1 _12039_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_17894_ _17895_/A _17895_/B _17895_/C vssd1 vssd1 vccd1 vccd1 _17896_/A sky130_fd_sc_hd__a21o_1
XFILLER_93_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19633_ _19605_/Y _19610_/Y _19612_/X vssd1 vssd1 vccd1 vccd1 _19634_/B sky130_fd_sc_hd__a21o_1
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16845_ _16845_/A _17189_/B _16845_/C _16845_/D vssd1 vssd1 vccd1 vccd1 _16846_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16091__A1 _15936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19564_ _19556_/Y _19557_/X _19555_/C _19555_/D vssd1 vssd1 vccd1 vccd1 _19564_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_16776_ _16776_/A _16776_/B _16776_/C vssd1 vssd1 vccd1 vccd1 _16777_/A sky130_fd_sc_hd__nand3_1
XFILLER_20_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13988_ _13984_/Y _13986_/Y _13987_/X vssd1 vssd1 vccd1 vccd1 _13992_/B sky130_fd_sc_hd__a21o_1
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12101__B1 _12098_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18368__B1 _12018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12369__B _12378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15727_ _15727_/A _15727_/B vssd1 vssd1 vccd1 vccd1 _15825_/A sky130_fd_sc_hd__nor2_1
X_18515_ _18706_/B _18999_/A _18507_/C _18680_/D _18510_/A vssd1 vssd1 vccd1 vccd1
+ _18653_/A sky130_fd_sc_hd__a32o_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _20576_/B _12681_/A _12681_/B _15696_/D _12973_/A vssd1 vssd1 vccd1 vccd1
+ _12981_/B sky130_fd_sc_hd__a32o_1
X_19495_ _19359_/X _19500_/A _19494_/Y vssd1 vssd1 vccd1 vccd1 _19497_/A sky130_fd_sc_hd__o21ai_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17241__A _19047_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18446_ _18613_/A vssd1 vssd1 vccd1 vccd1 _18451_/B sky130_fd_sc_hd__clkbuf_2
X_15658_ _15616_/A _16397_/A _16062_/A _16361_/A vssd1 vssd1 vccd1 vccd1 _15658_/Y
+ sky130_fd_sc_hd__o211ai_2
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14609_ _14604_/Y _14605_/X _14600_/Y _14602_/Y vssd1 vssd1 vccd1 vccd1 _14611_/C
+ sky130_fd_sc_hd__o211ai_1
X_18377_ _18311_/X _18353_/Y _18356_/Y _18376_/Y vssd1 vssd1 vccd1 vccd1 _18377_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_18_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_900 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15589_ _15589_/A vssd1 vssd1 vccd1 vccd1 _15589_/X sky130_fd_sc_hd__buf_2
XFILLER_147_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17328_ _17486_/A _17486_/B _17486_/C vssd1 vssd1 vccd1 vccd1 _17330_/B sky130_fd_sc_hd__nand3_1
XFILLER_105_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12816__C _22818_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17259_ _17145_/B _17247_/X _17249_/Y _17258_/X vssd1 vssd1 vccd1 vccd1 _17260_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_147_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19168__A _19318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15696__A _18848_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20270_ _20115_/A _20115_/B _20115_/C _20147_/B vssd1 vssd1 vccd1 vccd1 _20270_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_127_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11729__A _16256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17119__C _21019_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15657__A1 _15358_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19615__B _19772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22880__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19334__C _19842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22041__B _22041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22911_ _22916_/CLK _22911_/D vssd1 vssd1 vccd1 vccd1 _22911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21880__B _22173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22842_ _22943_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 _22842_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_582 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22773_ _22805_/CLK _22773_/D vssd1 vssd1 vccd1 vccd1 _22773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21724_ _21724_/A _21724_/B _21724_/C _21724_/D vssd1 vssd1 vccd1 vccd1 _21724_/Y
+ sky130_fd_sc_hd__nand4_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20265__A2_N _20266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21655_ _21618_/Y _21624_/Y _21647_/Y vssd1 vssd1 vccd1 vccd1 _21662_/A sky130_fd_sc_hd__o21ai_1
XFILLER_149_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20469__A1 _12734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20606_ _12671_/A _15412_/A _20605_/Y vssd1 vssd1 vccd1 vccd1 _20606_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__12946__A2 _20584_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21586_ _21582_/A _21583_/D _13319_/A vssd1 vssd1 vccd1 vccd1 _21757_/D sky130_fd_sc_hd__a21oi_2
XFILLER_138_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12445__D _20694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_914 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20537_ _20393_/C _20536_/X _20393_/A vssd1 vssd1 vccd1 vccd1 _20538_/C sky130_fd_sc_hd__o21ai_1
XFILLER_193_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12159__B1 _15377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_936 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20468_ _12702_/A _16708_/A _20460_/A vssd1 vssd1 vccd1 vccd1 _20468_/X sky130_fd_sc_hd__o21a_1
X_11270_ _22786_/Q vssd1 vssd1 vccd1 vccd1 _11306_/A sky130_fd_sc_hd__buf_2
XFILLER_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19626__A3 _19793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11639__A _11639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12174__A3 _12167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22207_ _22206_/C _22206_/A _22682_/Q vssd1 vssd1 vccd1 vccd1 _22208_/B sky130_fd_sc_hd__a21o_1
XFILLER_165_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17637__A2 _17444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20399_ _20155_/X _20156_/X _20154_/A vssd1 vssd1 vccd1 vccd1 _20399_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__15648__A1 _15918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15648__B2 _15646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22138_ _22138_/A _22138_/B vssd1 vssd1 vccd1 vccd1 _22140_/A sky130_fd_sc_hd__nand2_1
XFILLER_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14960_ _14960_/A _14960_/B vssd1 vssd1 vccd1 vccd1 _14961_/B sky130_fd_sc_hd__nand2_1
XFILLER_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16230__A _17251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22069_ _22072_/A _22072_/B _22068_/C _22068_/D vssd1 vssd1 vccd1 vccd1 _22079_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22394__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13911_ _13814_/A _13814_/B _13923_/A vssd1 vssd1 vccd1 vccd1 _13911_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13573__B _21944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input29_A wb_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ _15058_/C _14722_/C _14722_/A _14955_/A _14892_/C vssd1 vssd1 vccd1 vccd1
+ _14893_/A sky130_fd_sc_hd__a32o_1
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16630_ _16630_/A _16630_/B vssd1 vssd1 vccd1 vccd1 _16706_/A sky130_fd_sc_hd__nor2_2
X_13842_ _13985_/A vssd1 vssd1 vccd1 vccd1 _14013_/A sky130_fd_sc_hd__buf_2
XFILLER_63_828 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15820__A1 _15727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16561_ _16561_/A _16561_/B _16561_/C vssd1 vssd1 vccd1 vccd1 _16751_/A sky130_fd_sc_hd__nand3_4
XFILLER_90_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13773_ _13773_/A vssd1 vssd1 vccd1 vccd1 _14383_/A sky130_fd_sc_hd__buf_2
XFILLER_15_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18300_ _18305_/A _18305_/D _18299_/X vssd1 vssd1 vccd1 vccd1 _18301_/C sky130_fd_sc_hd__a21o_1
X_15512_ _15517_/A _15512_/B _15512_/C vssd1 vssd1 vccd1 vccd1 _15512_/Y sky130_fd_sc_hd__nand3_2
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19280_ _19301_/A _19301_/D vssd1 vssd1 vccd1 vccd1 _19282_/C sky130_fd_sc_hd__nand2_1
X_12724_ _12737_/A _12737_/B _12709_/Y _12723_/Y vssd1 vssd1 vccd1 vccd1 _12724_/Y
+ sky130_fd_sc_hd__a31oi_2
X_16492_ _16506_/A _16762_/A _16489_/X _16496_/A vssd1 vssd1 vccd1 vccd1 _16493_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17573__A1 _17574_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18231_ _18224_/Y _18226_/Y _18230_/Y vssd1 vssd1 vccd1 vccd1 _18231_/Y sky130_fd_sc_hd__a21oi_2
X_15443_ _17129_/B vssd1 vssd1 vccd1 vccd1 _19351_/C sky130_fd_sc_hd__buf_4
XFILLER_130_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12655_ _16153_/A vssd1 vssd1 vccd1 vccd1 _16157_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_128_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19314__A2 _19838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18162_ _18162_/A _18162_/B vssd1 vssd1 vccd1 vccd1 _18163_/C sky130_fd_sc_hd__nand2_1
X_11606_ _11285_/A _11285_/B _15377_/A vssd1 vssd1 vccd1 vccd1 _11606_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15374_ _15389_/B _15382_/B _15912_/C _17281_/B vssd1 vssd1 vccd1 vccd1 _15374_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_30_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12586_ _12586_/A vssd1 vssd1 vccd1 vccd1 _15559_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_128_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17113_ _19619_/B _17116_/A _17116_/B _17530_/A vssd1 vssd1 vccd1 vccd1 _17311_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_129_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14325_ _11395_/A _14317_/X _14320_/X _14322_/X _13776_/A vssd1 vssd1 vccd1 vccd1
+ _14325_/X sky130_fd_sc_hd__a32o_2
XFILLER_184_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18093_ _18093_/A _18093_/B _18093_/C _18093_/D vssd1 vssd1 vccd1 vccd1 _18093_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11537_ _11537_/A vssd1 vssd1 vccd1 vccd1 _11552_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17044_ _17208_/B _17041_/X _17043_/X vssd1 vssd1 vccd1 vccd1 _17603_/A sky130_fd_sc_hd__a21oi_4
XFILLER_171_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14256_ _14256_/A _14256_/B _14256_/C vssd1 vssd1 vccd1 vccd1 _14281_/A sky130_fd_sc_hd__nand3_1
X_11468_ _15901_/A _15415_/C _11942_/A _15901_/B vssd1 vssd1 vccd1 vccd1 _11468_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_171_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13207_ _22722_/Q _13234_/A _13234_/B _21580_/A _13202_/A vssd1 vssd1 vccd1 vccd1
+ _13517_/C sky130_fd_sc_hd__o311ai_4
XFILLER_48_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14187_ _14188_/B _14188_/C _14188_/A vssd1 vssd1 vccd1 vccd1 _14198_/A sky130_fd_sc_hd__a21o_1
XFILLER_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11399_ _11942_/A _16308_/C _11936_/C _16563_/C vssd1 vssd1 vccd1 vccd1 _11399_/Y
+ sky130_fd_sc_hd__nand4_4
XANTENNA__16836__B1 _16825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15639__B2 _15319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12570__B1 _12493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _13330_/A _21480_/B _13138_/C vssd1 vssd1 vccd1 vccd1 _13139_/B sky130_fd_sc_hd__and3_1
XFILLER_174_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18995_ _18995_/A _18995_/B vssd1 vssd1 vccd1 vccd1 _18996_/A sky130_fd_sc_hd__nor2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17946_ _17946_/A _17946_/B vssd1 vssd1 vccd1 vccd1 _18020_/C sky130_fd_sc_hd__nand2_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _22728_/Q vssd1 vssd1 vccd1 vccd1 _13301_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19154__C _19154_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22385__A1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17877_ _19987_/A _21048_/B _21048_/C _17922_/A _19987_/D vssd1 vssd1 vccd1 vccd1
+ _17877_/X sky130_fd_sc_hd__o32a_1
XANTENNA__11676__A2 _16482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19616_ _11821_/X _19624_/A _19625_/A _19462_/Y _19461_/X vssd1 vssd1 vccd1 vccd1
+ _19616_/X sky130_fd_sc_hd__o311a_1
X_16828_ _16828_/A _16828_/B _16831_/C vssd1 vssd1 vccd1 vccd1 _16986_/B sky130_fd_sc_hd__nand3_1
XFILLER_26_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1010 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19547_ _19457_/Y _19389_/X _19529_/A _19540_/Y vssd1 vssd1 vccd1 vccd1 _19552_/C
+ sky130_fd_sc_hd__o211a_1
X_16759_ _16759_/A _17139_/A _17140_/A vssd1 vssd1 vccd1 vccd1 _16956_/A sky130_fd_sc_hd__nand3_1
XFILLER_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17013__B1 _17025_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19478_ _19475_/Y _19476_/X _19477_/X vssd1 vssd1 vccd1 vccd1 _19630_/A sky130_fd_sc_hd__o21ai_4
XFILLER_62_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18429_ _18427_/X _18428_/Y _18425_/Y _18274_/Y vssd1 vssd1 vccd1 vccd1 _18601_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_166_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21440_ _21440_/A _21440_/B vssd1 vssd1 vccd1 vccd1 _21440_/Y sky130_fd_sc_hd__nand2_4
XFILLER_194_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20856__D1 _17525_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15327__B1 _15776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21371_ _21372_/A _21372_/B _21372_/C vssd1 vssd1 vccd1 vccd1 _21371_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12051__B1_N _11762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20322_ _12680_/X _16563_/A _16563_/B _20608_/A _20481_/C vssd1 vssd1 vccd1 vccd1
+ _20446_/A sky130_fd_sc_hd__a32o_1
XFILLER_163_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19048__D _19490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20253_ _20242_/X _20244_/X _20249_/B _20245_/X _15991_/B vssd1 vssd1 vccd1 vccd1
+ _20262_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_89_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20184_ _20184_/A _20184_/B _20184_/C vssd1 vssd1 vccd1 vccd1 _20304_/B sky130_fd_sc_hd__nand3_1
XFILLER_170_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22376__A1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_920 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14489__B _14489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20387__B1 _20337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17252__B1 _20129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22825_ _22929_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 _22825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17004__B1 _16554_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18201__C1 _12050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22756_ _22761_/CLK _22756_/D vssd1 vssd1 vccd1 vccd1 _22756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21707_ _21930_/A _21707_/B vssd1 vssd1 vccd1 vccd1 _21707_/X sky130_fd_sc_hd__or2_1
XFILLER_185_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22687_ _22944_/CLK _22687_/D vssd1 vssd1 vccd1 vccd1 _22687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_527 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12440_ _20461_/C vssd1 vssd1 vccd1 vccd1 _20456_/C sky130_fd_sc_hd__clkbuf_4
X_21638_ _21638_/A _21638_/B _21638_/C vssd1 vssd1 vccd1 vccd1 _21640_/C sky130_fd_sc_hd__nand3_1
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12371_ _20089_/B vssd1 vssd1 vccd1 vccd1 _20605_/B sky130_fd_sc_hd__buf_2
XFILLER_165_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21569_ _21568_/B _21568_/C _21568_/A vssd1 vssd1 vccd1 vccd1 _21570_/B sky130_fd_sc_hd__a21o_1
XFILLER_181_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16225__A _16225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14110_ _14110_/A _14110_/B _14110_/C vssd1 vssd1 vccd1 vccd1 _14113_/B sky130_fd_sc_hd__and3_1
XFILLER_153_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11322_ _22954_/Q _22953_/Q vssd1 vssd1 vccd1 vccd1 _11712_/A sky130_fd_sc_hd__nor2_2
XFILLER_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1111 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15090_ _14990_/X _15026_/B _15026_/C _14951_/A _15023_/Y vssd1 vssd1 vccd1 vccd1
+ _15092_/C sky130_fd_sc_hd__a32o_1
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14041_ _14220_/D _22863_/D vssd1 vssd1 vccd1 vccd1 _14098_/A sky130_fd_sc_hd__nand2_2
XFILLER_181_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16879__B _16879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17800_ _17800_/A _17800_/B _17910_/A _17800_/D vssd1 vssd1 vccd1 vccd1 _17800_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_122_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13584__A _21595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18780_ _18770_/A _18779_/B _18779_/A vssd1 vssd1 vccd1 vccd1 _18780_/X sky130_fd_sc_hd__a21o_1
X_15992_ _15649_/X _17539_/D _16049_/A _16051_/C vssd1 vssd1 vccd1 vccd1 _16047_/C
+ sky130_fd_sc_hd__a22o_2
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12304__B1 _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17731_ _17731_/A vssd1 vssd1 vccd1 vccd1 _17928_/A sky130_fd_sc_hd__buf_2
X_14943_ _14945_/C _15080_/C vssd1 vssd1 vccd1 vccd1 _14943_/X sky130_fd_sc_hd__and2_1
XFILLER_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17662_ _17662_/A _17662_/B vssd1 vssd1 vccd1 vccd1 _17665_/B sky130_fd_sc_hd__nand2_1
XFILLER_169_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14874_ _14880_/C vssd1 vssd1 vccd1 vccd1 _14877_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19401_ _19229_/B _19229_/C _19229_/A _19400_/X vssd1 vssd1 vccd1 vccd1 _19401_/X
+ sky130_fd_sc_hd__a31o_1
X_16613_ _16351_/X _17431_/C _16613_/C _16613_/D vssd1 vssd1 vccd1 vccd1 _16613_/X
+ sky130_fd_sc_hd__and4b_1
X_13825_ _13826_/A _13826_/B _22756_/Q vssd1 vssd1 vccd1 vccd1 _14069_/A sky130_fd_sc_hd__a21o_2
XFILLER_78_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17593_ _17520_/X _17467_/X _17591_/X vssd1 vssd1 vccd1 vccd1 _17624_/B sky130_fd_sc_hd__a21oi_1
XFILLER_18_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20210__A _20210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12928__A _12928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19332_ _19521_/A _19512_/A _19512_/B vssd1 vssd1 vccd1 vccd1 _19332_/Y sky130_fd_sc_hd__nand3_1
X_16544_ _16155_/A _17391_/A _16506_/X _16507_/X _16496_/X vssd1 vssd1 vccd1 vccd1
+ _16544_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13756_ _22858_/D vssd1 vssd1 vccd1 vccd1 _14230_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17546__A1 _12234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_574 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17546__B2 _17424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _12938_/A _16489_/A _12973_/A _20576_/B vssd1 vssd1 vccd1 vccd1 _12708_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_188_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19263_ _19257_/X _19258_/Y _19259_/Y _19262_/Y vssd1 vssd1 vccd1 vccd1 _19272_/B
+ sky130_fd_sc_hd__o211ai_1
X_16475_ _16248_/X _16060_/A _16472_/Y _16474_/Y vssd1 vssd1 vccd1 vccd1 _16475_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13687_ _22672_/Q _21294_/B vssd1 vssd1 vccd1 vccd1 _13689_/A sky130_fd_sc_hd__or2_1
XANTENNA__18615__A _18810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15426_ _15426_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15430_/B sky130_fd_sc_hd__nand2_1
X_18214_ _18214_/A _18214_/B _18214_/C vssd1 vssd1 vccd1 vccd1 _18214_/X sky130_fd_sc_hd__and3_1
X_19194_ _19194_/A _19490_/A _19490_/B _19194_/D vssd1 vssd1 vccd1 vccd1 _19194_/Y
+ sky130_fd_sc_hd__nand4_2
X_12638_ _16498_/A _20853_/A _20972_/D _16498_/D vssd1 vssd1 vccd1 vccd1 _12742_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18145_ _18137_/Y _18139_/X _18896_/C _15988_/A _18141_/Y vssd1 vssd1 vccd1 vccd1
+ _18146_/C sky130_fd_sc_hd__o2111ai_1
X_15357_ _15357_/A _20355_/A _16304_/A _18985_/C vssd1 vssd1 vccd1 vccd1 _15382_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA__14780__A1 _14953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12386__A3 _16319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20302__B1 _13045_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ _12470_/X _12520_/A _12549_/A _15363_/C _16319_/C vssd1 vssd1 vccd1 vccd1
+ _12571_/A sky130_fd_sc_hd__o311ai_4
XANTENNA__12663__A _15746_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14308_ _14370_/A vssd1 vssd1 vccd1 vccd1 _14308_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12791__B1 _20241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18076_ _18080_/A _18076_/B vssd1 vssd1 vccd1 vccd1 _18079_/A sky130_fd_sc_hd__nand2_1
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15288_ _15288_/A _22884_/Q _15288_/C vssd1 vssd1 vccd1 vccd1 _15290_/A sky130_fd_sc_hd__and3_1
XFILLER_145_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15396__D _17128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17027_ _17027_/A _17027_/B _17027_/C vssd1 vssd1 vccd1 vccd1 _17028_/C sky130_fd_sc_hd__nand3_1
XANTENNA__11279__A _22799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14239_ _14239_/A _14239_/B vssd1 vssd1 vccd1 vccd1 _14239_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11897__A2 _11909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20081__A2 _13022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _18978_/A _18978_/B vssd1 vssd1 vccd1 vccd1 _19117_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _17929_/A _21011_/C _21011_/A vssd1 vssd1 vccd1 vccd1 _17932_/A sky130_fd_sc_hd__and3_1
XFILLER_113_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16037__A1 _15962_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20940_ _20934_/X _20935_/Y _20939_/Y vssd1 vssd1 vccd1 vccd1 _20941_/C sky130_fd_sc_hd__a21o_1
XANTENNA__22957__D _22957_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18982__B1 _19772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20871_ _20871_/A _20871_/B vssd1 vssd1 vccd1 vccd1 _20871_/Y sky130_fd_sc_hd__nand2_1
XFILLER_183_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16993__C1 _20854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22610_ _22656_/S vssd1 vssd1 vccd1 vccd1 _22619_/S sky130_fd_sc_hd__buf_2
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22530__A1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22541_ _14362_/X input37/X _22547_/S vssd1 vssd1 vccd1 vccd1 _22542_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22472_ _22472_/A vssd1 vssd1 vccd1 vccd1 _22732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18244__B _18258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13574__A2 _21848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21423_ _21423_/A _21560_/A _21560_/B _21559_/B vssd1 vssd1 vccd1 vccd1 _21423_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_108_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12573__A _22821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14491__C _14491_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21354_ _21509_/A _21509_/B _21386_/A _21386_/B vssd1 vssd1 vccd1 vccd1 _21355_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_30_47 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20305_ _20292_/X _20296_/Y _20549_/A _20314_/C vssd1 vssd1 vccd1 vccd1 _20305_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_190_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21285_ _21820_/A _21289_/B _21285_/C _21424_/A vssd1 vssd1 vccd1 vccd1 _21292_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22597__A1 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19462__A1 _12111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20236_ _20236_/A _20236_/B _20236_/C vssd1 vssd1 vccd1 vccd1 _20240_/B sky130_fd_sc_hd__nand3_2
XFILLER_131_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15079__A2 _13851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__A _18830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20072__A2 _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20167_ _20167_/A _20167_/B _20167_/C vssd1 vssd1 vccd1 vccd1 _20170_/B sky130_fd_sc_hd__nand3_1
XFILLER_130_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20098_ _20478_/C _20098_/B _20101_/A _20098_/D vssd1 vssd1 vccd1 vccd1 _20098_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19091__A _19091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _11940_/A vssd1 vssd1 vccd1 vccd1 _18107_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_45_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13851__B _13851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15787__B1 _17133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ _18984_/A _18984_/B _11664_/D _19000_/A _18288_/A vssd1 vssd1 vccd1 vccd1
+ _11871_/X sky130_fd_sc_hd__a32o_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15251__A2 _15233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ _13617_/A _13617_/B _13609_/Y vssd1 vssd1 vccd1 vccd1 _13611_/C sky130_fd_sc_hd__a21oi_1
XFILLER_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22808_ _22808_/CLK _22808_/D vssd1 vssd1 vccd1 vccd1 _22808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14889_/D _14590_/B _15056_/B _14595_/B vssd1 vssd1 vccd1 vccd1 _14605_/D
+ sky130_fd_sc_hd__nand4_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22656__S _22656_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22521__A1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ _13527_/Y _13530_/X _13524_/A _13526_/X vssd1 vssd1 vccd1 vccd1 _13543_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_544 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22739_ _22771_/CLK _22739_/D vssd1 vssd1 vccd1 vccd1 _22739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16260_ _15557_/Y _16256_/Y _17133_/A _16258_/Y _18848_/C vssd1 vssd1 vccd1 vccd1
+ _16263_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_9_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13472_ _13516_/D vssd1 vssd1 vccd1 vccd1 _13563_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15211_ _15217_/A _15114_/A _15160_/A _15186_/X vssd1 vssd1 vccd1 vccd1 _15227_/A
+ sky130_fd_sc_hd__a31oi_4
X_12423_ _15326_/A _15325_/A _16256_/C vssd1 vssd1 vccd1 vccd1 _12461_/A sky130_fd_sc_hd__o21ai_1
XFILLER_127_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16191_ _16191_/A vssd1 vssd1 vccd1 vccd1 _20734_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_138_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15142_ _15101_/B _15101_/A _14987_/C vssd1 vssd1 vccd1 vccd1 _15143_/B sky130_fd_sc_hd__o21ai_1
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12354_ _12369_/A _12361_/A vssd1 vssd1 vccd1 vccd1 _12377_/A sky130_fd_sc_hd__nand2_2
XFILLER_154_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11305_ _12148_/A vssd1 vssd1 vccd1 vccd1 _11420_/A sky130_fd_sc_hd__clkbuf_2
X_19950_ _19905_/A _19937_/B _19905_/C _19939_/Y _19949_/B vssd1 vssd1 vccd1 vccd1
+ _19951_/B sky130_fd_sc_hd__o311a_1
X_15073_ _15073_/A _15108_/A _15073_/C vssd1 vssd1 vccd1 vccd1 _15074_/C sky130_fd_sc_hd__and3_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12285_ _22694_/Q vssd1 vssd1 vccd1 vccd1 _12368_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_181_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18170__A _19329_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18901_ _18901_/A vssd1 vssd1 vccd1 vccd1 _19085_/A sky130_fd_sc_hd__clkbuf_2
X_14024_ _14026_/C _14026_/D vssd1 vssd1 vccd1 vccd1 _14024_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19881_ _19881_/A _19881_/B _19881_/C vssd1 vssd1 vccd1 vccd1 _19881_/X sky130_fd_sc_hd__and3_1
XFILLER_136_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11879__A2 _18258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16402__B _16402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18832_ _18824_/X _19080_/A _18827_/Y _18831_/Y vssd1 vssd1 vccd1 vccd1 _19112_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_121_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15475__C1 _15755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15750__A1_N _15755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19205__A1 _11859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18763_ _18763_/A _18763_/B vssd1 vssd1 vccd1 vccd1 _18764_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15975_ _15975_/A _15975_/B vssd1 vssd1 vccd1 vccd1 _15976_/C sky130_fd_sc_hd__nand2_1
XANTENNA__22941__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17216__B1 _17215_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17714_ _17721_/C _17721_/A _22900_/Q vssd1 vssd1 vccd1 vccd1 _17716_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__21012__B2 _17922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14926_ _14982_/A _14982_/C vssd1 vssd1 vccd1 vccd1 _14927_/B sky130_fd_sc_hd__and2_1
X_18694_ _11800_/X _19160_/A _18707_/A vssd1 vssd1 vccd1 vccd1 _18702_/A sky130_fd_sc_hd__o21ai_1
XFILLER_76_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17645_ _17652_/B _18830_/D _19768_/D _17645_/D vssd1 vssd1 vccd1 vccd1 _17645_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13761__B _13761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14857_ _14857_/A _14857_/B _15070_/A vssd1 vssd1 vccd1 vccd1 _14952_/B sky130_fd_sc_hd__and3_1
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19508__A2 _18629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13808_ _13808_/A _13881_/A vssd1 vssd1 vccd1 vccd1 _13808_/Y sky130_fd_sc_hd__nor2_2
XFILLER_56_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17576_ _17627_/A _17581_/B vssd1 vssd1 vccd1 vccd1 _17578_/A sky130_fd_sc_hd__nand2_1
X_14788_ _14793_/A _14793_/B _14862_/A _14685_/B vssd1 vssd1 vccd1 vccd1 _14788_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14450__B1 _14448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22512__A1 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16990__A2 _16822_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19315_ _18699_/A _18699_/B _11511_/X vssd1 vssd1 vccd1 vccd1 _19315_/X sky130_fd_sc_hd__a21o_1
X_16527_ _15545_/X _12922_/X _16476_/X _16515_/Y _16479_/X vssd1 vssd1 vccd1 vccd1
+ _16527_/X sky130_fd_sc_hd__o221a_1
XFILLER_143_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13739_ _13963_/B vssd1 vssd1 vccd1 vccd1 _13833_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11712__D _15482_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19246_ _19246_/A _19246_/B vssd1 vssd1 vccd1 vccd1 _19246_/Y sky130_fd_sc_hd__nand2_1
X_16458_ _18445_/A _18797_/B _12938_/A _15997_/C _16471_/A vssd1 vssd1 vccd1 vccd1
+ _16458_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_192_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15409_ _15409_/A vssd1 vssd1 vccd1 vccd1 _15412_/A sky130_fd_sc_hd__clkbuf_4
X_16389_ _16372_/X _16388_/Y _16636_/A _16378_/X vssd1 vssd1 vccd1 vccd1 _16393_/A
+ sky130_fd_sc_hd__o22ai_1
X_19177_ _17427_/X _19176_/X _19174_/A vssd1 vssd1 vccd1 vccd1 _19179_/A sky130_fd_sc_hd__o21ai_2
XFILLER_192_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11567__A1 _11561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18128_ _18128_/A _18128_/B _18128_/C vssd1 vssd1 vccd1 vccd1 _18129_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19692__A1 _17380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22028__B1 _21841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19176__A _19176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14505__A1 _14818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18059_ _18019_/Y _17999_/A _18042_/A vssd1 vssd1 vccd1 vccd1 _18059_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21070_ _21065_/X _21070_/B _22941_/Q vssd1 vssd1 vccd1 vccd1 _21074_/A sky130_fd_sc_hd__nand3b_1
XFILLER_125_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20115__A _20115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16258__A1 _16059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20021_ _20020_/B _20021_/B vssd1 vssd1 vccd1 vccd1 _20022_/B sky130_fd_sc_hd__and2b_1
XFILLER_101_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17424__A _17424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15870__C _17816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21972_ _21972_/A _21972_/B _21972_/C _21972_/D vssd1 vssd1 vccd1 vccd1 _22030_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20923_ _20923_/A _20923_/B _20923_/C vssd1 vssd1 vccd1 vccd1 _20936_/D sky130_fd_sc_hd__nand3_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16430__B2 _16397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20854_ _20854_/A _20854_/B _21011_/B vssd1 vssd1 vccd1 vccd1 _20854_/Y sky130_fd_sc_hd__nand3_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14441__B1 _22952_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20109__A3 _20098_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20785_ _20685_/A _15940_/A _20784_/Y vssd1 vssd1 vccd1 vccd1 _20787_/C sky130_fd_sc_hd__o21ai_2
XFILLER_168_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22524_ _22524_/A vssd1 vssd1 vccd1 vccd1 _22755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_655 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16733__A2 _16726_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22455_ _22512_/S vssd1 vssd1 vccd1 vccd1 _22464_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20817__A1 _20818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21406_ _21406_/A _21406_/B _21406_/C vssd1 vssd1 vccd1 vccd1 _21417_/B sky130_fd_sc_hd__nand3_2
XANTENNA__12622__A2_N _12602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22386_ _22386_/A vssd1 vssd1 vccd1 vccd1 _22694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21337_ _21336_/B _13098_/A _13301_/X vssd1 vssd1 vccd1 vccd1 _21338_/B sky130_fd_sc_hd__a21bo_1
XFILLER_190_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19435__A1 _19418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12070_ _12064_/X _11914_/Y _12069_/X _11918_/A vssd1 vssd1 vccd1 vccd1 _12070_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21268_ _21268_/A vssd1 vssd1 vccd1 vccd1 _21269_/A sky130_fd_sc_hd__buf_2
XANTENNA__22964__CLK _22964_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16249__A1 _16248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20219_ _20219_/A _20219_/B vssd1 vssd1 vccd1 vccd1 _20219_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21199_ _21609_/A vssd1 vssd1 vccd1 vccd1 _22229_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_bq_clk_i clkbuf_4_9_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _22949_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _15862_/A _15864_/D _15759_/Y vssd1 vssd1 vccd1 vccd1 _15761_/C sky130_fd_sc_hd__a21oi_1
XFILLER_46_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _16100_/D vssd1 vssd1 vccd1 vccd1 _16106_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17749__A1 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18946__B1 _18627_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input11_A wb_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _14716_/A _14716_/B _14711_/C _14711_/D vssd1 vssd1 vccd1 vccd1 _14714_/B
+ sky130_fd_sc_hd__nand4_1
X_11923_ _11923_/A _11923_/B vssd1 vssd1 vccd1 vccd1 _11924_/D sky130_fd_sc_hd__nand2_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15691_ _14431_/A _15808_/A _16498_/D _15690_/X vssd1 vssd1 vccd1 vccd1 _15691_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _17313_/A _19336_/A _17431_/B _17431_/D vssd1 vssd1 vccd1 vccd1 _17430_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14642_ _14505_/X _14640_/Y _14516_/C vssd1 vssd1 vccd1 vccd1 _14642_/Y sky130_fd_sc_hd__o21ai_1
X_11854_ _18810_/A vssd1 vssd1 vccd1 vccd1 _19418_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17361_ _17361_/A _17370_/A _17370_/B _17361_/D vssd1 vssd1 vccd1 vccd1 _17361_/Y
+ sky130_fd_sc_hd__nand4_2
X_14573_ _14573_/A _14573_/B vssd1 vssd1 vccd1 vccd1 _14688_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16709__C1 _20098_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ _12127_/A _18325_/A vssd1 vssd1 vccd1 vccd1 _12010_/A sky130_fd_sc_hd__nand2_2
XANTENNA__15004__D _15004_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19100_ _19117_/A _19117_/B _19117_/C vssd1 vssd1 vccd1 vccd1 _19303_/A sky130_fd_sc_hd__nand3_1
X_16312_ _16552_/A vssd1 vssd1 vccd1 vccd1 _16312_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13524_ _13524_/A vssd1 vssd1 vccd1 vccd1 _13524_/X sky130_fd_sc_hd__clkbuf_2
X_17292_ _19336_/A _17449_/A _17293_/B _20793_/C vssd1 vssd1 vccd1 vccd1 _17292_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_158_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17382__C1 _20928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16243_ _15536_/X _16240_/X _16228_/Y _16241_/Y _16242_/X vssd1 vssd1 vccd1 vccd1
+ _16498_/C sky130_fd_sc_hd__a32oi_2
XFILLER_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19031_ _19689_/A _19334_/B _19013_/B _19012_/X vssd1 vssd1 vccd1 vccd1 _19031_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15301__B _16257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13455_ _13455_/A _13455_/B _13455_/C vssd1 vssd1 vccd1 vccd1 _13455_/Y sky130_fd_sc_hd__nand3_1
XFILLER_127_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11549__A1 _11401_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_3_0_bq_clk_i_A clkbuf_4_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12406_ _20359_/B _12844_/A _12400_/X _20358_/A _12487_/B vssd1 vssd1 vccd1 vccd1
+ _12407_/B sky130_fd_sc_hd__o221ai_1
X_16174_ _16174_/A _16174_/B _16111_/A vssd1 vssd1 vccd1 vccd1 _16174_/X sky130_fd_sc_hd__or3b_1
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13386_ _21251_/A _21249_/A vssd1 vssd1 vccd1 vccd1 _13390_/B sky130_fd_sc_hd__nand2_1
XANTENNA__22415__A _22426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18331__D1 _19322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15125_ _15064_/C _15050_/C _15050_/A _15122_/X _15124_/Y vssd1 vssd1 vccd1 vccd1
+ _15128_/C sky130_fd_sc_hd__a311o_1
Xoutput108 _14336_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[4] sky130_fd_sc_hd__buf_2
X_12337_ _12822_/B vssd1 vssd1 vccd1 vccd1 _15631_/C sky130_fd_sc_hd__clkbuf_2
Xoutput119 _22667_/Q vssd1 vssd1 vccd1 vccd1 y[3] sky130_fd_sc_hd__buf_2
XFILLER_142_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12941__A _16489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19933_ _19973_/A _19975_/A _19891_/Y _19976_/C _19976_/A vssd1 vssd1 vccd1 vccd1
+ _19934_/B sky130_fd_sc_hd__o2111ai_1
X_15056_ _15056_/A _15056_/B vssd1 vssd1 vccd1 vccd1 _15057_/A sky130_fd_sc_hd__nand2_1
X_12268_ _22693_/Q vssd1 vssd1 vccd1 vccd1 _12273_/B sky130_fd_sc_hd__clkbuf_4
X_14007_ _14007_/A _14007_/B vssd1 vssd1 vccd1 vccd1 _14033_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11557__A _22959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19864_ _19864_/A _19864_/B vssd1 vssd1 vccd1 vccd1 _19865_/A sky130_fd_sc_hd__nand2_1
XFILLER_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12199_ _12046_/A _12208_/B _11727_/C vssd1 vssd1 vccd1 vccd1 _12212_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__13475__C _13475_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput90 _14390_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[17] sky130_fd_sc_hd__buf_2
X_18815_ _18814_/X _12204_/X _18830_/C _18828_/A vssd1 vssd1 vccd1 vccd1 _18818_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_68_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15999__B1 _17085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21692__C _21809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19795_ _17421_/X _17422_/X _18843_/A _18843_/B vssd1 vssd1 vccd1 vccd1 _19795_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13772__A _22871_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18746_ _18744_/Y _18745_/Y _18646_/C vssd1 vssd1 vccd1 vccd1 _18746_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15958_ _15937_/X _15942_/X _15947_/Y _15949_/A vssd1 vssd1 vccd1 vccd1 _15964_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14909_ _13833_/X _13736_/B _15082_/A _14963_/A _14908_/Y vssd1 vssd1 vccd1 vccd1
+ _14909_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18677_ _18677_/A _18677_/B _18677_/C vssd1 vssd1 vccd1 vccd1 _18678_/B sky130_fd_sc_hd__and3_1
X_15889_ _15887_/X _16155_/A _12968_/D _15888_/X vssd1 vssd1 vccd1 vccd1 _15889_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__20101__C _20101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17628_ _17628_/A vssd1 vssd1 vccd1 vccd1 _17628_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14423__B1 _14413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17559_ _17559_/A _17559_/B _17559_/C vssd1 vssd1 vccd1 vccd1 _17580_/A sky130_fd_sc_hd__nand3_2
XANTENNA__11338__A_N _11334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22837__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20570_ _20519_/C _20569_/Y _20519_/B vssd1 vssd1 vccd1 vccd1 _20745_/A sky130_fd_sc_hd__o21ai_2
XFILLER_177_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12835__B _20092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19229_ _19229_/A _19229_/B _19229_/C vssd1 vssd1 vccd1 vccd1 _19244_/A sky130_fd_sc_hd__nand3_1
XANTENNA__13529__A2 _13050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18803__A _19202_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22240_ _22240_/A _22240_/B _22240_/C vssd1 vssd1 vccd1 vccd1 _22241_/B sky130_fd_sc_hd__and3_1
XFILLER_145_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17023__A2_N _16732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21867__C _21938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22171_ _22171_/A _22171_/B vssd1 vssd1 vccd1 vccd1 _22173_/A sky130_fd_sc_hd__nand2_1
XFILLER_132_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11960__A1 _11751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21122_ _21122_/A _21122_/B vssd1 vssd1 vccd1 vccd1 _21122_/X sky130_fd_sc_hd__and2_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17428__B1 _11672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__A _15776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21053_ _21053_/A _21081_/D vssd1 vssd1 vccd1 vccd1 _21054_/B sky130_fd_sc_hd__xor2_1
XFILLER_141_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20578__A3 _17875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20004_ _20026_/A vssd1 vssd1 vccd1 vccd1 _20024_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input3_A wb_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19353__B _19353_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16651__A1 _15646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13682__A _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21955_ _21185_/X _21187_/X _21724_/B _22229_/A vssd1 vssd1 vccd1 vccd1 _22042_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20906_ _20828_/A _20906_/B _20906_/C vssd1 vssd1 vccd1 vccd1 _20906_/Y sky130_fd_sc_hd__nand3b_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14414__B1 _14413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21886_ _21886_/A _21886_/B vssd1 vssd1 vccd1 vccd1 _21892_/C sky130_fd_sc_hd__nand2_1
XFILLER_42_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ _20902_/A _20902_/B _22936_/Q vssd1 vssd1 vccd1 vccd1 _20837_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12448__D _20694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ _19318_/A vssd1 vssd1 vccd1 vccd1 _19465_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_20768_ _20768_/A _22934_/Q _20768_/C vssd1 vssd1 vccd1 vccd1 _20768_/Y sky130_fd_sc_hd__nand3_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22507_ _22507_/A vssd1 vssd1 vccd1 vccd1 _22748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20699_ _20699_/A vssd1 vssd1 vccd1 vccd1 _20797_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13240_ _13240_/A _13257_/A vssd1 vssd1 vccd1 vccd1 _13273_/B sky130_fd_sc_hd__nand2_1
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22438_ _22438_/A vssd1 vssd1 vccd1 vccd1 _22718_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14193__A2 _14494_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13171_ _22841_/Q vssd1 vssd1 vccd1 vccd1 _21588_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22369_ input68/X input67/X input34/X _22369_/D vssd1 vssd1 vccd1 vccd1 _22426_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_164_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11951__A1 _11859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12122_ _15694_/A _18848_/D _11956_/C _11943_/B _11938_/Y vssd1 vssd1 vccd1 vccd1
+ _12123_/C sky130_fd_sc_hd__a32o_2
XFILLER_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15142__A1 _15101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input59_A wb_dat_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16930_ _16930_/A _17341_/A _16930_/C vssd1 vssd1 vccd1 vccd1 _16988_/B sky130_fd_sc_hd__nand3_1
XFILLER_105_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ _12029_/Y _12039_/Y _12081_/A vssd1 vssd1 vccd1 vccd1 _12245_/B sky130_fd_sc_hd__a21o_1
XFILLER_117_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11703__A1 _11381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18631__A2 _18303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16861_ _16535_/A _16535_/B _16541_/X _16546_/Y _16534_/B vssd1 vssd1 vccd1 vccd1
+ _16861_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18600_ _18600_/A vssd1 vssd1 vccd1 vccd1 _19281_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15812_ _15824_/A _15824_/B _15812_/C _15812_/D vssd1 vssd1 vccd1 vccd1 _15886_/A
+ sky130_fd_sc_hd__nand4_1
X_19580_ _19580_/A vssd1 vssd1 vccd1 vccd1 _19580_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16792_ _16792_/A _16792_/B vssd1 vssd1 vccd1 vccd1 _16803_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18531_ _18531_/A vssd1 vssd1 vccd1 vccd1 _18664_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15743_ _15298_/Y _15309_/A _15304_/B _15457_/A vssd1 vssd1 vccd1 vccd1 _15743_/X
+ sky130_fd_sc_hd__o211a_1
X_12955_ _12937_/Y _12944_/X _12954_/Y vssd1 vssd1 vccd1 vccd1 _12957_/A sky130_fd_sc_hd__o21a_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20726__B1 _20449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21017__C _21017_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17198__A2 _17025_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _18305_/B vssd1 vssd1 vccd1 vccd1 _18953_/C sky130_fd_sc_hd__buf_4
XFILLER_33_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_712 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18462_ _18462_/A _18474_/B vssd1 vssd1 vccd1 vccd1 _18462_/Y sky130_fd_sc_hd__nand2_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15666_/A _15668_/X _15673_/B _15673_/C vssd1 vssd1 vccd1 vccd1 _15677_/C
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12886_ _12886_/A _12886_/B vssd1 vssd1 vccd1 vccd1 _12886_/X sky130_fd_sc_hd__or2_1
XANTENNA__16945__A2 _15723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17383_/Y _17385_/Y _17412_/X vssd1 vssd1 vccd1 vccd1 _17413_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11837_ _11831_/C _11837_/B _12084_/A vssd1 vssd1 vccd1 vccd1 _12246_/B sky130_fd_sc_hd__nand3b_1
XFILLER_33_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14625_ _14616_/Y _14614_/Y _15188_/A _13924_/X vssd1 vssd1 vccd1 vccd1 _14625_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_18393_ _18407_/A _18407_/B _18396_/C _18559_/A vssd1 vssd1 vccd1 vccd1 _18393_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_650 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _17340_/Y _17342_/X _17350_/A vssd1 vssd1 vccd1 vccd1 _17344_/Y sky130_fd_sc_hd__o21bai_1
X_14556_ _22672_/D _14987_/C _14554_/B _14555_/X vssd1 vssd1 vccd1 vccd1 _22673_/D
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__20575__D _20870_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11768_ _12127_/A vssd1 vssd1 vccd1 vccd1 _19197_/A sky130_fd_sc_hd__buf_2
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13507_ _21724_/B vssd1 vssd1 vccd1 vccd1 _22106_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19719__A _19788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17275_ _17464_/B vssd1 vssd1 vccd1 vccd1 _17275_/Y sky130_fd_sc_hd__inv_2
X_14487_ _14684_/A vssd1 vssd1 vccd1 vccd1 _15006_/A sky130_fd_sc_hd__buf_2
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11699_ _11644_/A _11645_/A _11645_/B _11553_/B _11552_/B vssd1 vssd1 vccd1 vccd1
+ _11699_/X sky130_fd_sc_hd__a32o_1
X_19014_ _19014_/A vssd1 vssd1 vccd1 vccd1 _19014_/X sky130_fd_sc_hd__clkbuf_2
X_16226_ _16226_/A _16226_/B _16226_/C vssd1 vssd1 vccd1 vccd1 _16227_/A sky130_fd_sc_hd__nor3_4
XFILLER_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13438_ _13438_/A _13438_/B vssd1 vssd1 vccd1 vccd1 _13438_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15966__B _16192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21687__C _21687_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16157_ _16157_/A _16157_/B _16157_/C _16157_/D vssd1 vssd1 vccd1 vccd1 _16157_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_127_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ _13213_/X _13364_/Y _21638_/B _13367_/Y _13572_/A vssd1 vssd1 vccd1 vccd1
+ _13385_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_177_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ _15108_/A vssd1 vssd1 vccd1 vccd1 _15108_/Y sky130_fd_sc_hd__inv_2
X_16088_ _15971_/A _15927_/Y _15886_/Y vssd1 vssd1 vccd1 vccd1 _16088_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11287__A _22954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19916_ _19916_/A _19916_/B vssd1 vssd1 vccd1 vccd1 _19917_/B sky130_fd_sc_hd__xor2_1
XANTENNA__14341__C1 _14340_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15039_ _15039_/A _15047_/B vssd1 vssd1 vccd1 vccd1 _15040_/B sky130_fd_sc_hd__or2b_1
XANTENNA__19454__A _19651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16881__B2 _16880_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19847_ _19353_/B _19353_/C _19985_/C _19846_/B _19846_/C vssd1 vssd1 vccd1 vccd1
+ _19850_/C sky130_fd_sc_hd__a32o_1
XANTENNA__19173__B _19358_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19778_ _19848_/B _19783_/B _19781_/B vssd1 vssd1 vccd1 vccd1 _19787_/A sky130_fd_sc_hd__a21o_1
XFILLER_113_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18729_ _18729_/A vssd1 vssd1 vccd1 vccd1 _18729_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11458__B1 _14429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21740_ _21868_/A vssd1 vssd1 vccd1 vccd1 _21740_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21224__A _21621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21671_ _21677_/A _21677_/B vssd1 vssd1 vccd1 vccd1 _21671_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12846__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16318__A _16318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20622_ _20602_/Y _20603_/X _20626_/A vssd1 vssd1 vccd1 vccd1 _20631_/A sky130_fd_sc_hd__o21bai_1
XFILLER_138_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20553_ _20553_/A _20553_/B vssd1 vssd1 vccd1 vccd1 _20554_/C sky130_fd_sc_hd__nand2_1
XFILLER_193_956 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20484_ _20499_/A _20499_/B vssd1 vssd1 vccd1 vccd1 _20484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22223_ _22223_/A vssd1 vssd1 vccd1 vccd1 _22304_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18846__C1 _19358_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20102__D1 _16261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22154_ _22154_/A vssd1 vssd1 vccd1 vccd1 _22938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16321__B1 _14369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11909__B _11909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21105_ _21074_/B _21124_/A _21074_/A vssd1 vssd1 vccd1 vccd1 _21106_/B sky130_fd_sc_hd__a21boi_1
XFILLER_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22085_ _22025_/Y _21932_/Y _22160_/A _22084_/Y vssd1 vssd1 vccd1 vccd1 _22090_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_102_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21036_ _21008_/X _21062_/A _21031_/X vssd1 vssd1 vccd1 vccd1 _21067_/B sky130_fd_sc_hd__a21o_1
XANTENNA__20303__A _20442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11449__B1 _15435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19023__C1 _18856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_712 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12740_ _12920_/C _12732_/Y _13002_/B vssd1 vssd1 vccd1 vccd1 _12741_/C sky130_fd_sc_hd__o21ai_1
X_21938_ _22182_/A _21938_/B _22182_/C vssd1 vssd1 vccd1 vccd1 _21939_/B sky130_fd_sc_hd__nand3_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12671_/A vssd1 vssd1 vccd1 vccd1 _12671_/X sky130_fd_sc_hd__buf_2
XFILLER_163_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21869_ _21742_/B _21871_/A _21972_/A vssd1 vssd1 vccd1 vccd1 _21880_/A sky130_fd_sc_hd__o21ai_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12756__A _15746_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14410_ _14410_/A vssd1 vssd1 vccd1 vccd1 _14410_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _12062_/A _11415_/A _18133_/A vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__o21ai_1
XFILLER_42_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15390_ _15664_/A _15665_/A _15388_/Y _15389_/X vssd1 vssd1 vccd1 vccd1 _15512_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ _12273_/B _14308_/X _14337_/X _13131_/X _14340_/X vssd1 vssd1 vccd1 vccd1
+ _14341_/X sky130_fd_sc_hd__a221o_1
XFILLER_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _11553_/A _11553_/B vssd1 vssd1 vccd1 vccd1 _11554_/C sky130_fd_sc_hd__nand2_1
XFILLER_184_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17060_ _17060_/A _17060_/B vssd1 vssd1 vccd1 vccd1 _17215_/D sky130_fd_sc_hd__nand2_2
XFILLER_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14272_ _14272_/A _14276_/D _14272_/C _14272_/D vssd1 vssd1 vccd1 vccd1 _14279_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_183_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16560__B1 _17281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11484_ _11615_/A vssd1 vssd1 vccd1 vccd1 _11980_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16011_ _16011_/A _16011_/B vssd1 vssd1 vccd1 vccd1 _16012_/B sky130_fd_sc_hd__and2_1
XFILLER_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13223_ _13384_/B _13385_/A _13384_/A vssd1 vssd1 vccd1 vccd1 _13223_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20644__C1 _20737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13154_ _13513_/B vssd1 vssd1 vccd1 vccd1 _21362_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_163_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12105_ _11771_/X _11770_/X _18313_/B _18674_/A vssd1 vssd1 vccd1 vccd1 _12108_/A
+ sky130_fd_sc_hd__o211ai_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _17959_/A _17920_/A _17953_/B vssd1 vssd1 vccd1 vccd1 _17962_/Y sky130_fd_sc_hd__a21oi_2
X_13085_ _21351_/A _21351_/B _21476_/C vssd1 vssd1 vccd1 vccd1 _13300_/A sky130_fd_sc_hd__nand3_4
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19701_ _19590_/X _19588_/A _19690_/X vssd1 vssd1 vccd1 vccd1 _19703_/B sky130_fd_sc_hd__a21o_1
X_16913_ _17110_/A vssd1 vssd1 vccd1 vccd1 _16913_/X sky130_fd_sc_hd__clkbuf_2
X_12036_ _12036_/A vssd1 vssd1 vccd1 vccd1 _12036_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17893_ _17893_/A _17893_/B vssd1 vssd1 vccd1 vccd1 _17895_/C sky130_fd_sc_hd__nand2_1
XFILLER_78_664 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19632_ _19611_/X _19613_/Y _19631_/Y vssd1 vssd1 vccd1 vccd1 _19635_/A sky130_fd_sc_hd__o21ai_2
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16844_ _16541_/X _16546_/Y _16534_/B _16843_/Y vssd1 vssd1 vccd1 vccd1 _16846_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__22682__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16091__A2 _20728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19563_ _19411_/X _19562_/Y _19559_/Y vssd1 vssd1 vccd1 vccd1 _19563_/Y sky130_fd_sc_hd__a21oi_1
X_16775_ _16494_/X _16760_/X _16954_/A _16774_/X vssd1 vssd1 vccd1 vccd1 _16776_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12101__A1 _12117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13987_ _13899_/A _13899_/B _14074_/A vssd1 vssd1 vccd1 vccd1 _13987_/X sky130_fd_sc_hd__a21o_1
XANTENNA__18368__B2 _16921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18514_ _16241_/A _11988_/X _15893_/A _18706_/B _18876_/B vssd1 vssd1 vccd1 vccd1
+ _18514_/Y sky130_fd_sc_hd__o2111ai_4
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ _15723_/X _15725_/Y _17108_/B _15649_/X _15959_/A vssd1 vssd1 vccd1 vccd1
+ _15727_/B sky130_fd_sc_hd__o2111a_2
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19494_ _15839_/A _18856_/A _19352_/A vssd1 vssd1 vccd1 vccd1 _19494_/Y sky130_fd_sc_hd__o21ai_2
X_12938_ _12938_/A vssd1 vssd1 vccd1 vccd1 _15774_/D sky130_fd_sc_hd__buf_2
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17241__B _20928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18445_ _18445_/A _18797_/B _18445_/C vssd1 vssd1 vccd1 vccd1 _18613_/A sky130_fd_sc_hd__nand3_1
X_15657_ _15358_/X _16737_/A _16431_/A vssd1 vssd1 vccd1 vccd1 _15657_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _12509_/A _12564_/B _12865_/Y vssd1 vssd1 vccd1 vccd1 _12872_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11570__A _19318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15042__A _15175_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14608_ _14580_/X _14601_/Y _14606_/Y _14607_/Y vssd1 vssd1 vccd1 vccd1 _14740_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18376_ _18396_/A _18396_/B vssd1 vssd1 vccd1 vccd1 _18376_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15588_ _16215_/A _16215_/B _16530_/C vssd1 vssd1 vccd1 vccd1 _15588_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17327_ _17472_/B vssd1 vssd1 vccd1 vccd1 _17486_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15977__A _16011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14539_ _14524_/Y _14534_/X _14537_/Y _14538_/Y vssd1 vssd1 vccd1 vccd1 _14547_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17258_ _12294_/A _12294_/B _15538_/X _15541_/X vssd1 vssd1 vccd1 vccd1 _17258_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15696__B _16912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19168__B _19461_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16209_ _16209_/A _16403_/A _16209_/C vssd1 vssd1 vccd1 vccd1 _16210_/D sky130_fd_sc_hd__nand3_1
XFILLER_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17189_ _17189_/A _17189_/B vssd1 vssd1 vccd1 vccd1 _17189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11376__C1 _11306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11915__A1 _16157_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11729__B _16256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15657__A2 _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19615__C _19615_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22910_ _22922_/CLK _22910_/D vssd1 vssd1 vccd1 vccd1 _22910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_612 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22841_ _22937_/CLK hold5/X vssd1 vssd1 vccd1 vccd1 _22841_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18359__A1 _12018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21880__C _22057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12279__C _15363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22772_ _22772_/CLK _22772_/D vssd1 vssd1 vccd1 vccd1 _22772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_594 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_907 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21723_ _21767_/A _21455_/X _21610_/A _21610_/B vssd1 vssd1 vccd1 vccd1 _21730_/B
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__11851__B1 _17313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16048__A _17539_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19308__B1 _11511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11480__A _12094_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14494__C _14494_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21654_ _21654_/A _21654_/B _21654_/C vssd1 vssd1 vccd1 vccd1 _21654_/X sky130_fd_sc_hd__and3_1
XANTENNA__20793__A _20793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20605_ _20605_/A _20605_/B _20675_/C vssd1 vssd1 vccd1 vccd1 _20605_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__20469__A2 _16611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15887__A _15887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21585_ _21588_/C vssd1 vssd1 vccd1 vccd1 _21937_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20536_ _20844_/A _16179_/X _20263_/B _20264_/A _20263_/A vssd1 vssd1 vccd1 vccd1
+ _20536_/X sky130_fd_sc_hd__o221a_1
XFILLER_153_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12159__A1 _12157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13356__B1 _13141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22615__A0 _22796_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20467_ _20464_/A _20464_/B _20462_/A _20587_/A vssd1 vssd1 vccd1 vccd1 _20495_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_4_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13200__A _21473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22206_ _22206_/A _22682_/Q _22206_/C vssd1 vssd1 vccd1 vccd1 _22208_/A sky130_fd_sc_hd__nand3_1
XFILLER_134_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20398_ _20398_/A vssd1 vssd1 vccd1 vccd1 _20398_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15648__A2 _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22137_ _22196_/A _22196_/B _22137_/C _22137_/D vssd1 vssd1 vccd1 vccd1 _22138_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22068_ _22072_/A _22072_/B _22068_/C _22068_/D vssd1 vssd1 vccd1 vccd1 _22079_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_59_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11655__A _22960_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21019_ _21019_/A _21019_/B _21050_/C vssd1 vssd1 vccd1 vccd1 _21020_/B sky130_fd_sc_hd__and3_1
X_13910_ _13904_/Y _13905_/Y _13909_/Y vssd1 vssd1 vccd1 vccd1 _13937_/A sky130_fd_sc_hd__o21ai_2
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14890_ _15107_/A _15107_/B _14808_/D _14889_/D _14808_/B vssd1 vssd1 vccd1 vccd1
+ _14892_/C sky130_fd_sc_hd__a32o_1
XFILLER_75_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13841_ _13892_/A _13821_/B _13892_/B _13869_/B vssd1 vssd1 vccd1 vccd1 _13985_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15820__A2 _15727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16560_ _16295_/Y _16550_/Y _17281_/B _16552_/Y _15711_/A vssd1 vssd1 vccd1 vccd1
+ _16561_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_16_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13772_ _22871_/Q vssd1 vssd1 vccd1 vccd1 _14503_/A sky130_fd_sc_hd__clkinv_2
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15511_ _15738_/A vssd1 vssd1 vccd1 vccd1 _15859_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12723_ _12933_/C _12933_/D vssd1 vssd1 vccd1 vccd1 _12723_/Y sky130_fd_sc_hd__nand2_1
X_16491_ _16494_/A _16491_/B vssd1 vssd1 vccd1 vccd1 _16496_/A sky130_fd_sc_hd__nand2_2
XFILLER_128_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17573__A2 _17574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18230_ _18227_/X _18229_/X _18272_/B vssd1 vssd1 vccd1 vccd1 _18230_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15442_ _16473_/B vssd1 vssd1 vccd1 vccd1 _17129_/B sky130_fd_sc_hd__buf_2
XFILLER_128_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12654_ _16067_/B vssd1 vssd1 vccd1 vccd1 _16153_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22394__S _22402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_940 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ _11605_/A vssd1 vssd1 vccd1 vccd1 _15377_/A sky130_fd_sc_hd__buf_2
XFILLER_156_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15797__A _15797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18161_ _12164_/Y _12168_/X _18165_/A vssd1 vssd1 vccd1 vccd1 _18162_/B sky130_fd_sc_hd__o21ai_1
X_12585_ _15466_/B vssd1 vssd1 vccd1 vccd1 _15559_/C sky130_fd_sc_hd__clkbuf_4
X_15373_ _20593_/B vssd1 vssd1 vccd1 vccd1 _17281_/B sky130_fd_sc_hd__buf_2
XFILLER_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_984 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17112_ _17116_/A _17116_/B _16015_/A _17732_/A vssd1 vssd1 vccd1 vccd1 _17311_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_129_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15336__A1 _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14324_ _12876_/X _14308_/X _14313_/X _13659_/C _14323_/X vssd1 vssd1 vccd1 vccd1
+ _14324_/X sky130_fd_sc_hd__a221o_1
X_11536_ _11536_/A _11536_/B _11536_/C vssd1 vssd1 vccd1 vccd1 _11537_/A sky130_fd_sc_hd__nand3_1
X_18092_ _11737_/X _11738_/X _11846_/B _12003_/A _15810_/A vssd1 vssd1 vccd1 vccd1
+ _18092_/Y sky130_fd_sc_hd__o2111ai_4
XANTENNA__11740__A1_N _11736_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19419__D _19455_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22606__A0 _11771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17043_ _16885_/B _16884_/X _17042_/Y vssd1 vssd1 vccd1 vccd1 _17043_/X sky130_fd_sc_hd__a21o_1
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14255_ _14255_/A _14255_/B _14255_/C vssd1 vssd1 vccd1 vccd1 _14256_/C sky130_fd_sc_hd__nand3_1
X_11467_ _15776_/B vssd1 vssd1 vccd1 vccd1 _15901_/B sky130_fd_sc_hd__buf_4
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13206_ _22720_/Q vssd1 vssd1 vccd1 vccd1 _13234_/B sky130_fd_sc_hd__buf_2
XANTENNA__18286__B1 _18203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14186_ _14274_/A _14561_/C _14119_/Y _14185_/X vssd1 vssd1 vccd1 vccd1 _14188_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_139_1141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11398_ _18876_/C vssd1 vssd1 vccd1 vccd1 _16563_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16836__A1 _19615_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _22843_/Q vssd1 vssd1 vccd1 vccd1 _21480_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18994_ _18495_/A _18495_/B _15981_/X vssd1 vssd1 vccd1 vccd1 _18995_/B sky130_fd_sc_hd__a21o_2
XFILLER_151_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _17945_/A _17945_/B vssd1 vssd1 vccd1 vccd1 _17946_/B sky130_fd_sc_hd__nand2_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _21188_/C vssd1 vssd1 vccd1 vccd1 _13073_/A sky130_fd_sc_hd__buf_2
X_12019_ _12018_/X _15888_/A _11425_/Y _18508_/A _12001_/Y vssd1 vssd1 vccd1 vccd1
+ _12019_/X sky130_fd_sc_hd__o221a_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17876_ _17876_/A vssd1 vssd1 vccd1 vccd1 _19987_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19615_ _19615_/A _19772_/B _19615_/C vssd1 vssd1 vccd1 vccd1 _19615_/X sky130_fd_sc_hd__and3_1
XFILLER_38_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16827_ _16828_/A _16828_/B _16831_/C vssd1 vssd1 vccd1 vccd1 _16986_/A sky130_fd_sc_hd__a21o_1
XFILLER_4_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19546_ _19650_/A _19540_/Y _19543_/Y vssd1 vssd1 vccd1 vccd1 _19552_/A sky130_fd_sc_hd__a21oi_1
XFILLER_81_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16758_ _16758_/A vssd1 vssd1 vccd1 vccd1 _16758_/X sky130_fd_sc_hd__buf_4
XFILLER_0_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15709_ _15748_/A _15709_/B _15709_/C vssd1 vssd1 vccd1 vccd1 _15709_/Y sky130_fd_sc_hd__nand3_2
X_19477_ _15580_/X _19839_/D _19323_/X _19330_/B vssd1 vssd1 vccd1 vccd1 _19477_/X
+ sky130_fd_sc_hd__o31a_1
X_16689_ _16690_/C _16690_/A _22891_/Q vssd1 vssd1 vccd1 vccd1 _16698_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1047 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18428_ _18232_/X _18233_/Y _18224_/Y vssd1 vssd1 vccd1 vccd1 _18428_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_167_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18359_ _12018_/X _16921_/X _18367_/A _18367_/B vssd1 vssd1 vccd1 vccd1 _18471_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_147_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15327__A1 _15325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21370_ _21522_/C _22849_/Q _21522_/A vssd1 vssd1 vccd1 vccd1 _21372_/C sky130_fd_sc_hd__and3_1
XFILLER_190_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19329__D _19329_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20321_ _20295_/Y _20181_/A _20319_/Y _20320_/Y vssd1 vssd1 vccd1 vccd1 _20549_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_174_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13020__A _16106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16034__C _16034_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_bq_clk_i clkbuf_3_5_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _22964_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_150_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20252_ _20246_/Y _20249_/Y _20251_/Y vssd1 vssd1 vccd1 vccd1 _20252_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_131_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_992 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17427__A _17427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20183_ _20183_/A _20183_/B vssd1 vssd1 vccd1 vccd1 _20184_/C sky130_fd_sc_hd__nand2_1
XFILLER_142_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20153__B1_N _20125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_932 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16055__A2 _15983_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18258__A _18258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22824_ _22850_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 _22824_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18201__B1 _17632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22755_ _22757_/CLK _22755_/D vssd1 vssd1 vccd1 vccd1 _22755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16209__C _16209_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21706_ _21706_/A _21832_/A vssd1 vssd1 vccd1 vccd1 _21711_/A sky130_fd_sc_hd__nand2_1
XFILLER_158_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22686_ _22943_/CLK _22686_/D vssd1 vssd1 vccd1 vccd1 _22686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21637_ _21352_/X _21607_/X _21499_/X vssd1 vssd1 vccd1 vccd1 _21640_/B sky130_fd_sc_hd__a21o_1
XFILLER_100_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19162__D1 _19156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15318__A1 _15482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ _16323_/A _16323_/B _12403_/D _16293_/A vssd1 vssd1 vccd1 vccd1 _20089_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21568_ _21568_/A _21568_/B _21568_/C vssd1 vssd1 vccd1 vccd1 _21570_/A sky130_fd_sc_hd__nand3_1
XFILLER_126_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11321_ _18338_/C vssd1 vssd1 vccd1 vccd1 _18875_/D sky130_fd_sc_hd__buf_2
XFILLER_181_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20519_ _20519_/A _20519_/B _20519_/C vssd1 vssd1 vccd1 vccd1 _20623_/B sky130_fd_sc_hd__and3_1
XFILLER_125_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21499_ _21338_/A _21338_/B _13504_/A vssd1 vssd1 vccd1 vccd1 _21499_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14040_ _14273_/A vssd1 vssd1 vccd1 vccd1 _14220_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_158_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16879__C _17840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16241__A _16241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input41_A wb_dat_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15991_ _16129_/A _15991_/B _16129_/C _15991_/D vssd1 vssd1 vccd1 vccd1 _16051_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12304__A1 _12387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17730_ _17730_/A vssd1 vssd1 vccd1 vccd1 _17873_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14942_ _14942_/A _14942_/B _14942_/C vssd1 vssd1 vccd1 vccd1 _15080_/C sky130_fd_sc_hd__or3_1
XFILLER_76_932 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21575__B1 _21421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17661_ _17661_/A _17661_/B vssd1 vssd1 vccd1 vccd1 _17662_/B sky130_fd_sc_hd__nor2_1
X_14873_ _14793_/B _14998_/C _14575_/B _14933_/A _14872_/Y vssd1 vssd1 vccd1 vccd1
+ _14880_/C sky130_fd_sc_hd__o2111ai_2
XANTENNA__18168__A _19199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20783__D1 _17385_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19400_ _19400_/A _19400_/B vssd1 vssd1 vccd1 vccd1 _19400_/X sky130_fd_sc_hd__and2_1
XANTENNA__18991__A1 _11541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16612_ _11541_/X _17435_/A _15645_/X vssd1 vssd1 vccd1 vccd1 _16613_/D sky130_fd_sc_hd__o21ai_4
X_13824_ _13820_/X _13821_/Y _13831_/A _13823_/Y vssd1 vssd1 vccd1 vccd1 _13824_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_91_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17592_ _17467_/X _17520_/X _17624_/A _17625_/A _17591_/X vssd1 vssd1 vccd1 vccd1
+ _17597_/B sky130_fd_sc_hd__a221o_1
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20210__B _20210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19331_ _19174_/B _19334_/A _19167_/Y _19016_/Y vssd1 vssd1 vccd1 vccd1 _19512_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16543_ _16758_/A vssd1 vssd1 vccd1 vccd1 _17391_/A sky130_fd_sc_hd__clkbuf_4
X_13755_ _13968_/C vssd1 vssd1 vccd1 vccd1 _14191_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17546__A2 _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19262_ _19148_/X _19150_/Y _19260_/X _19261_/Y vssd1 vssd1 vccd1 vccd1 _19262_/Y
+ sky130_fd_sc_hd__o22ai_1
X_12706_ _16759_/A vssd1 vssd1 vccd1 vccd1 _16489_/A sky130_fd_sc_hd__buf_2
X_16474_ _16474_/A _16782_/A vssd1 vssd1 vccd1 vccd1 _16474_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__20550__A1 _20442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13686_ _21426_/A vssd1 vssd1 vccd1 vccd1 _21294_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18615__B _19353_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18213_ _18232_/A _18232_/B _18232_/C vssd1 vssd1 vccd1 vccd1 _18226_/C sky130_fd_sc_hd__nand3_2
XANTENNA__13568__B1 _21498_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15425_ _15331_/Y _15329_/X _15344_/X vssd1 vssd1 vccd1 vccd1 _15426_/A sky130_fd_sc_hd__o21ai_1
X_19193_ _19504_/A _19694_/B _19052_/A _19055_/Y _19062_/B vssd1 vssd1 vccd1 vccd1
+ _19201_/A sky130_fd_sc_hd__a32oi_4
X_12637_ _16486_/C vssd1 vssd1 vccd1 vccd1 _16498_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_86_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22870__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18144_ _12131_/Y _12134_/B _12126_/X _12128_/X vssd1 vssd1 vccd1 vccd1 _18146_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_141_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12568_ _15299_/D vssd1 vssd1 vccd1 vccd1 _12681_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__20302__A1 _12754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15356_ _20477_/A vssd1 vssd1 vccd1 vccd1 _16304_/A sky130_fd_sc_hd__buf_4
XFILLER_184_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11519_ _11968_/B vssd1 vssd1 vccd1 vccd1 _18339_/C sky130_fd_sc_hd__clkbuf_2
X_14307_ _22369_/D vssd1 vssd1 vccd1 vccd1 _14370_/A sky130_fd_sc_hd__buf_2
XANTENNA__12791__B2 _12929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18075_ _22907_/Q _18075_/B _18082_/B vssd1 vssd1 vccd1 vccd1 _18076_/B sky130_fd_sc_hd__nand3b_1
XFILLER_176_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_594 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15287_ _22881_/Q _22882_/Q _22883_/Q _15287_/D vssd1 vssd1 vccd1 vccd1 _15288_/A
+ sky130_fd_sc_hd__or4_2
X_12499_ _12479_/B _12543_/A _20255_/B _15455_/A vssd1 vssd1 vccd1 vccd1 _12503_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_17026_ _17027_/A _17027_/B _17024_/X _17025_/X vssd1 vssd1 vccd1 vccd1 _17028_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_144_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14238_ _14238_/A _14238_/B vssd1 vssd1 vccd1 vccd1 _14239_/A sky130_fd_sc_hd__nand2_1
XFILLER_160_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20066__B1 _20065_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14169_ _14169_/A _14169_/B _14169_/C vssd1 vssd1 vccd1 vccd1 _14169_/X sky130_fd_sc_hd__and3_1
XFILLER_112_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _18977_/A _18977_/B vssd1 vssd1 vccd1 vccd1 _18978_/B sky130_fd_sc_hd__nand2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11295__A _11295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17928_ _17928_/A _19941_/B _19899_/B _17928_/D vssd1 vssd1 vccd1 vccd1 _17928_/X
+ sky130_fd_sc_hd__or4_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20369__A1 _20250_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16037__A2 _15959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17859_ _17858_/Y _17778_/Y _17787_/A _17787_/B vssd1 vssd1 vccd1 vccd1 _17860_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14599__A2 _13873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20870_ _20870_/A _20870_/B _20870_/C vssd1 vssd1 vccd1 vccd1 _20877_/A sky130_fd_sc_hd__and3_1
XFILLER_54_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19529_ _19529_/A vssd1 vssd1 vccd1 vccd1 _19650_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17314__A2_N _19482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19931__B1 _22923_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12557__C _16486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22540_ _22540_/A vssd1 vssd1 vccd1 vccd1 _22762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22471_ _21307_/B input38/X _22475_/S vssd1 vssd1 vccd1 vccd1 _22472_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15230__A _15230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21422_ _21422_/A _21422_/B vssd1 vssd1 vccd1 vccd1 _21559_/B sky130_fd_sc_hd__nand2_2
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21353_ _13326_/Y _21352_/X _21220_/X _21349_/X _21460_/A vssd1 vssd1 vccd1 vccd1
+ _21509_/B sky130_fd_sc_hd__o311a_1
XFILLER_163_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20304_ _20304_/A _20304_/B vssd1 vssd1 vccd1 vccd1 _20304_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21284_ _21423_/A _21424_/C vssd1 vssd1 vccd1 vccd1 _21289_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20235_ _20236_/A _20236_/B _20236_/C vssd1 vssd1 vccd1 vccd1 _20240_/A sky130_fd_sc_hd__a21o_1
XFILLER_104_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19462__A2 _19160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11742__C1 _11438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11917__B _16106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20166_ _20293_/B _20161_/B _20162_/A vssd1 vssd1 vccd1 vccd1 _20170_/A sky130_fd_sc_hd__o21ai_1
XFILLER_77_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16996__A _16996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21557__B1 _21838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20097_ _12577_/X _12576_/X _12687_/B _12578_/A vssd1 vssd1 vccd1 vccd1 _20098_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15405__A _15893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15787__A1 _16192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ _16563_/C vssd1 vssd1 vccd1 vccd1 _19000_/A sky130_fd_sc_hd__buf_4
XFILLER_73_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15787__B2 _15991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22807_ _22807_/CLK _22807_/D vssd1 vssd1 vccd1 vccd1 _22807_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20999_ _20999_/A _20999_/B _22939_/Q vssd1 vssd1 vccd1 vccd1 _21076_/B sky130_fd_sc_hd__nand3_1
XANTENNA__18716__A _18716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22893__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12467__C _22821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13540_ _13460_/A _13460_/B _13537_/A vssd1 vssd1 vccd1 vccd1 _13543_/A sky130_fd_sc_hd__o21ai_1
X_22738_ _22738_/CLK _22738_/D vssd1 vssd1 vccd1 vccd1 _22738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11371__C _15357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14963__B _14963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _13447_/X _13446_/X _13169_/X vssd1 vssd1 vccd1 vccd1 _13471_/Y sky130_fd_sc_hd__a21oi_1
X_22669_ _22964_/CLK _22669_/D vssd1 vssd1 vccd1 vccd1 _22669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15210_ _15210_/A _15210_/B vssd1 vssd1 vccd1 vccd1 _15210_/X sky130_fd_sc_hd__or2_1
X_12422_ _12447_/A vssd1 vssd1 vccd1 vccd1 _16256_/C sky130_fd_sc_hd__buf_2
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16190_ _16190_/A _16190_/B vssd1 vssd1 vccd1 vccd1 _16195_/A sky130_fd_sc_hd__nand2_1
XFILLER_154_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15141_ _15100_/A _15135_/X _15136_/Y _15173_/B vssd1 vssd1 vccd1 vccd1 _15175_/B
+ sky130_fd_sc_hd__a31o_2
X_12353_ _12802_/A vssd1 vssd1 vccd1 vccd1 _15633_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_127_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11304_ _11764_/A vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15072_ _15108_/A _15073_/C _15073_/A vssd1 vssd1 vccd1 vccd1 _15074_/B sky130_fd_sc_hd__a21oi_1
X_12284_ _12284_/A vssd1 vssd1 vccd1 vccd1 _12402_/A sky130_fd_sc_hd__buf_2
XFILLER_84_1010 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18900_ _18900_/A vssd1 vssd1 vccd1 vccd1 _18908_/B sky130_fd_sc_hd__clkbuf_2
X_14023_ _22873_/Q _13709_/A _13954_/A _13954_/B vssd1 vssd1 vccd1 vccd1 _14026_/D
+ sky130_fd_sc_hd__a22o_1
X_19880_ _19880_/A _19880_/B _19880_/C _19880_/D vssd1 vssd1 vccd1 vccd1 _19880_/Y
+ sky130_fd_sc_hd__nand4_2
X_18831_ _18825_/A _19079_/A _18829_/X _18830_/X vssd1 vssd1 vccd1 vccd1 _18831_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_150_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15475__B1 _12672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18762_ _18762_/A _18762_/B _18762_/C vssd1 vssd1 vccd1 vccd1 _18770_/A sky130_fd_sc_hd__nand3_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19205__A2 _11861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15974_ _15504_/X _15427_/X _15900_/A _15813_/Y _15778_/Y vssd1 vssd1 vccd1 vccd1
+ _15976_/B sky130_fd_sc_hd__o221ai_1
XFILLER_67_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__C _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17713_ _17713_/A _17713_/B vssd1 vssd1 vccd1 vccd1 _17721_/A sky130_fd_sc_hd__nand2_1
XANTENNA__21012__A2 _21048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17216__B2 _17373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14925_ _14756_/B _14839_/Y _14838_/B _14840_/Y vssd1 vssd1 vccd1 vccd1 _14982_/C
+ sky130_fd_sc_hd__o211ai_1
X_18693_ _18695_/A _18877_/A _18692_/Y vssd1 vssd1 vccd1 vccd1 _18707_/A sky130_fd_sc_hd__o21ai_1
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20221__A _20355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17644_ _17535_/Y _17533_/X _17643_/X vssd1 vssd1 vccd1 vccd1 _17654_/A sky130_fd_sc_hd__a21oi_1
XFILLER_1_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14856_ _15010_/A vssd1 vssd1 vccd1 vccd1 _15070_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13807_ _13807_/A _14270_/A _14892_/A vssd1 vssd1 vccd1 vccd1 _13807_/Y sky130_fd_sc_hd__nand3_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17575_ _17573_/Y _17575_/B _17575_/C vssd1 vssd1 vccd1 vccd1 _17581_/B sky130_fd_sc_hd__nand3b_2
XFILLER_56_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14787_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14862_/A sky130_fd_sc_hd__buf_2
XFILLER_17_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11999_ _12170_/A _12171_/A _15633_/A vssd1 vssd1 vccd1 vccd1 _12001_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_670 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19314_ _16098_/X _19838_/A _19156_/D _19156_/Y _19311_/Y vssd1 vssd1 vccd1 vccd1
+ _19340_/B sky130_fd_sc_hd__o311a_2
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16526_ _16472_/Y _16474_/Y _16513_/X vssd1 vssd1 vccd1 vccd1 _16526_/X sky130_fd_sc_hd__o21a_1
XANTENNA__17530__A _17530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13738_ _13738_/A vssd1 vssd1 vccd1 vccd1 _13963_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__16727__B1 _16582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19245_ _19400_/A _19400_/B vssd1 vssd1 vccd1 vccd1 _19245_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16457_ _15522_/A _15521_/A _15523_/A vssd1 vssd1 vccd1 vccd1 _16471_/A sky130_fd_sc_hd__a21oi_2
XFILLER_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13669_ _13665_/Y _13660_/X _13667_/X _13668_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_32_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12674__A _12742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15408_ _15397_/Y _15513_/B _15513_/A vssd1 vssd1 vccd1 vccd1 _15700_/B sky130_fd_sc_hd__nand3b_2
X_19176_ _19176_/A vssd1 vssd1 vccd1 vccd1 _19176_/X sky130_fd_sc_hd__buf_2
XFILLER_192_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16388_ _16388_/A vssd1 vssd1 vccd1 vccd1 _16388_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11567__A2 _11563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13961__B1 _14112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18127_ _18679_/C _18127_/B vssd1 vssd1 vccd1 vccd1 _18128_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15339_ _15339_/A _15339_/B _15339_/C vssd1 vssd1 vccd1 vccd1 _15664_/A sky130_fd_sc_hd__nand3_2
XFILLER_118_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19692__A2 _17381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18058_ _18058_/A vssd1 vssd1 vccd1 vccd1 _22966_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15702__A1 _15978_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14505__A2 _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12516__A1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17009_ _16990_/Y _16991_/Y _17006_/Y _17008_/Y vssd1 vssd1 vccd1 vccd1 _17009_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20115__B _20115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20020_ _20021_/B _20020_/B vssd1 vssd1 vccd1 vccd1 _20022_/A sky130_fd_sc_hd__and2b_1
XANTENNA__17455__A1 _17457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16258__A2 _16274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21227__A _21848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21971_ _21767_/X _21970_/X _21740_/X _22045_/A vssd1 vssd1 vccd1 vccd1 _21972_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_132_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15870__D _17039_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_475 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11753__A _16447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20922_ _20923_/B _20923_/C _20923_/A vssd1 vssd1 vccd1 vccd1 _20922_/X sky130_fd_sc_hd__a21o_1
XFILLER_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20853_ _20853_/A vssd1 vssd1 vccd1 vccd1 _21011_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14441__A1 _18259_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17440__A _17440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16718__B1 _16712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20784_ _20676_/B _20780_/Y _20782_/Y vssd1 vssd1 vccd1 vccd1 _20784_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22523_ _13725_/A input60/X _22525_/S vssd1 vssd1 vccd1 vccd1 _22524_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17930__A2 _17880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22454_ _22454_/A vssd1 vssd1 vccd1 vccd1 _22724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21405_ _21403_/Y _21404_/Y _21390_/Y _21401_/Y vssd1 vssd1 vccd1 vccd1 _21406_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_182_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20817__A2 _20818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22385_ _12413_/X input63/X _22391_/S vssd1 vssd1 vccd1 vccd1 _22386_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21336_ _13301_/X _21336_/B _21336_/C vssd1 vssd1 vccd1 vccd1 _21338_/A sky130_fd_sc_hd__nand3b_2
XFILLER_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18891__B1 _19587_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21267_ _21265_/Y _21266_/Y _21263_/Y _21257_/Y vssd1 vssd1 vccd1 vccd1 _21267_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16249__A2 _16179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20218_ _20218_/A _20457_/A vssd1 vssd1 vccd1 vccd1 _20224_/A sky130_fd_sc_hd__nand2_2
X_21198_ _13662_/A _21606_/A _21970_/A _21195_/Y _21197_/Y vssd1 vssd1 vccd1 vccd1
+ _21198_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_106_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20149_ _20154_/A _20154_/B _20149_/C _20149_/D vssd1 vssd1 vccd1 vccd1 _20150_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_103_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _15893_/C vssd1 vssd1 vccd1 vccd1 _16100_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_58_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12759__A _12988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18946__A1 _18953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11663__A _19322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14710_ _14710_/A _14716_/C vssd1 vssd1 vccd1 vccd1 _14714_/A sky130_fd_sc_hd__nand2_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11922_ _11922_/A _11922_/B _11922_/C vssd1 vssd1 vccd1 vccd1 _11923_/B sky130_fd_sc_hd__nand3_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _16257_/B vssd1 vssd1 vccd1 vccd1 _15690_/X sky130_fd_sc_hd__buf_6
XFILLER_18_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _14505_/X _14640_/Y _14512_/A _14044_/B _14516_/C vssd1 vssd1 vccd1 vccd1
+ _14646_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _18107_/A vssd1 vssd1 vccd1 vccd1 _18810_/A sky130_fd_sc_hd__buf_2
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _17060_/A _17060_/B _16665_/A vssd1 vssd1 vccd1 vccd1 _17361_/D sky130_fd_sc_hd__a21oi_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16709__B1 _16715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11784_ _12130_/A vssd1 vssd1 vccd1 vccd1 _18325_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__20505__A1 _15631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14572_ _14571_/X _14775_/A _14362_/X vssd1 vssd1 vccd1 vccd1 _14573_/B sky130_fd_sc_hd__o21ai_1
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16311_ _15888_/A _15792_/C _15792_/A _15938_/A _15887_/A vssd1 vssd1 vccd1 vccd1
+ _16311_/X sky130_fd_sc_hd__o32a_1
XFILLER_159_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _13523_/A _13523_/B _13523_/C vssd1 vssd1 vccd1 vccd1 _13524_/A sky130_fd_sc_hd__nand3_1
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17291_ _17464_/B _17464_/A vssd1 vssd1 vccd1 vccd1 _17291_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17382__B1 _20928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19030_ _19504_/A vssd1 vssd1 vccd1 vccd1 _19689_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16242_ _16242_/A _16242_/B vssd1 vssd1 vccd1 vccd1 _16242_/X sky130_fd_sc_hd__and2_1
XFILLER_186_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13454_ _13516_/D _13454_/B vssd1 vssd1 vccd1 vccd1 _13455_/C sky130_fd_sc_hd__nand2_1
XFILLER_167_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19123__A1 _18812_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11549__A2 _11895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ _16294_/A _16293_/A _12687_/B _16302_/A vssd1 vssd1 vccd1 vccd1 _20358_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_173_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16173_ _16169_/C _16118_/C _16172_/Y _16141_/X vssd1 vssd1 vccd1 vccd1 _16173_/Y
+ sky130_fd_sc_hd__o22ai_1
X_13385_ _13385_/A _13385_/B _13385_/C _13385_/D vssd1 vssd1 vccd1 vccd1 _21249_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18331__C1 _19322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ _15146_/A _15121_/X _15123_/X vssd1 vssd1 vccd1 vccd1 _15124_/Y sky130_fd_sc_hd__a21oi_1
Xoutput109 _14341_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[5] sky130_fd_sc_hd__buf_2
X_12336_ _22695_/Q _22694_/Q vssd1 vssd1 vccd1 vccd1 _12822_/B sky130_fd_sc_hd__nor2_2
XFILLER_126_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12941__B _15696_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19932_ _19976_/A _19891_/Y _19976_/C _19973_/A _19975_/A vssd1 vssd1 vccd1 vccd1
+ _19971_/B sky130_fd_sc_hd__a311o_1
XFILLER_114_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15055_ _15055_/A _15128_/A vssd1 vssd1 vccd1 vccd1 _15074_/A sky130_fd_sc_hd__nand2_1
X_12267_ _12824_/A _12303_/A vssd1 vssd1 vccd1 vccd1 _12387_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17437__A1 _17442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14006_ _14006_/A _14006_/B _14006_/C vssd1 vssd1 vccd1 vccd1 _14035_/A sky130_fd_sc_hd__nand3_1
X_19863_ _19796_/B _19794_/B _19859_/Y _19860_/Y vssd1 vssd1 vccd1 vccd1 _19863_/Y
+ sky130_fd_sc_hd__a211oi_4
X_12198_ _16226_/C _12208_/B _16242_/A _15486_/C vssd1 vssd1 vccd1 vccd1 _12202_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__15448__B1 _16106_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput91 _14393_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[18] sky130_fd_sc_hd__buf_2
X_18814_ _18814_/A vssd1 vssd1 vccd1 vccd1 _18814_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17525__A _19772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19794_ _19790_/Y _19794_/B _19794_/C vssd1 vssd1 vccd1 vccd1 _19860_/A sky130_fd_sc_hd__nand3b_2
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18745_ _18933_/C vssd1 vssd1 vccd1 vccd1 _18745_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15957_ _16035_/C _15957_/B _15957_/C vssd1 vssd1 vccd1 vccd1 _16422_/A sky130_fd_sc_hd__nand3b_2
XFILLER_37_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12669__A _12669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14671__A1 _13930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ _14905_/X _14907_/Y _14816_/B vssd1 vssd1 vccd1 vccd1 _14908_/Y sky130_fd_sc_hd__o21ai_1
X_18676_ _18698_/B _18676_/B _18841_/C vssd1 vssd1 vccd1 vccd1 _18857_/A sky130_fd_sc_hd__nand3_2
X_15888_ _15888_/A vssd1 vssd1 vccd1 vccd1 _15888_/X sky130_fd_sc_hd__buf_4
XFILLER_91_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17627_ _17627_/A vssd1 vssd1 vccd1 vccd1 _17627_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14839_ _14839_/A _14839_/B vssd1 vssd1 vccd1 vccd1 _14839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17558_ _17390_/Y _17556_/X _17557_/Y vssd1 vssd1 vccd1 vccd1 _17559_/C sky130_fd_sc_hd__o21ai_1
XFILLER_108_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16509_ _16506_/X _16507_/X _16496_/A vssd1 vssd1 vccd1 vccd1 _16509_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_177_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17489_ _17490_/A _17490_/B _17490_/C vssd1 vssd1 vccd1 vccd1 _17491_/A sky130_fd_sc_hd__a21o_1
XFILLER_108_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19228_ _19206_/Y _19211_/X _19227_/Y _19208_/A vssd1 vssd1 vccd1 vccd1 _19229_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_149_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12198__C1 _15486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18803__B _19353_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19159_ _19386_/A vssd1 vssd1 vccd1 vccd1 _19530_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17676__A1 _15840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22170_ _22170_/A _22170_/B vssd1 vssd1 vccd1 vccd1 _22194_/A sky130_fd_sc_hd__nand2_1
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11960__A2 _11703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21121_ _21119_/A _21119_/B _22943_/Q vssd1 vssd1 vccd1 vccd1 _21127_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__20680__B1 _12721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11748__A _11762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19417__A2 _19203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17428__A1 _14432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18625__B1 _17647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21052_ _21090_/B _21052_/B vssd1 vssd1 vccd1 vccd1 _21081_/D sky130_fd_sc_hd__nand2_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20003_ _20001_/Y _20002_/Y _19999_/Y vssd1 vssd1 vccd1 vccd1 _20026_/A sky130_fd_sc_hd__o21bai_1
XFILLER_143_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17435__A _17435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19353__C _19353_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16651__A2 _15645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21954_ _22036_/A _22064_/A vssd1 vssd1 vccd1 vccd1 _21977_/A sky130_fd_sc_hd__nand2_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20905_ _20905_/A _20905_/B vssd1 vssd1 vccd1 vccd1 _22917_/D sky130_fd_sc_hd__xor2_2
XFILLER_27_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21885_ _21762_/B _21884_/X _21760_/B vssd1 vssd1 vccd1 vccd1 _21886_/A sky130_fd_sc_hd__o21a_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _20834_/X _20835_/X _20994_/A _20840_/A _20840_/B vssd1 vssd1 vccd1 vccd1
+ _20902_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_70_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20767_ _20776_/A _22935_/Q _20776_/C vssd1 vssd1 vccd1 vccd1 _20772_/C sky130_fd_sc_hd__nand3_1
XFILLER_195_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22506_ _22748_/Q input55/X _22508_/S vssd1 vssd1 vccd1 vccd1 _22507_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20698_ _20695_/A _20695_/B _20696_/Y _20697_/Y vssd1 vssd1 vccd1 vccd1 _20699_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_11_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22437_ _22718_/Q input58/X _22439_/S vssd1 vssd1 vccd1 vccd1 _22438_/A sky130_fd_sc_hd__mux2_1
XANTENNA__21420__A _21421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13170_ _13099_/B _21336_/C _13095_/X vssd1 vssd1 vccd1 vccd1 _13170_/Y sky130_fd_sc_hd__a21oi_1
X_22368_ _22368_/A _22368_/B vssd1 vssd1 vccd1 vccd1 _22948_/D sky130_fd_sc_hd__nor2_1
XFILLER_191_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15775__D _17085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ _18648_/B vssd1 vssd1 vccd1 vccd1 _18848_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__11658__A _11712_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11951__A2 _11861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21319_ _13662_/A _21958_/A _21466_/A _21466_/B _21467_/A vssd1 vssd1 vccd1 vccd1
+ _21320_/C sky130_fd_sc_hd__o221ai_2
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22299_ _22299_/A vssd1 vssd1 vccd1 vccd1 _22941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12052_ _12052_/A _12240_/B vssd1 vssd1 vccd1 vccd1 _12081_/A sky130_fd_sc_hd__xor2_2
XFILLER_117_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14350__B1 _14337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11703__A2 _12111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20663__A2_N _20827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16860_ _16860_/A _16860_/B _16860_/C vssd1 vssd1 vccd1 vccd1 _16873_/C sky130_fd_sc_hd__nand3_2
XFILLER_104_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18631__A3 _18303_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14688__B _14785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15811_ _15823_/A vssd1 vssd1 vccd1 vccd1 _15812_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16791_ _16778_/A _16779_/A _19358_/A _19358_/B vssd1 vssd1 vccd1 vccd1 _16792_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18530_ _18156_/A _11702_/X _19316_/A _18330_/A vssd1 vssd1 vccd1 vccd1 _18531_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_93_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19041__B1 _17393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15742_ _19587_/A vssd1 vssd1 vccd1 vccd1 _19772_/D sky130_fd_sc_hd__buf_4
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _12954_/A _12954_/B _12954_/C vssd1 vssd1 vccd1 vccd1 _12954_/Y sky130_fd_sc_hd__nand3_1
XFILLER_93_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18461_ _18464_/A _18461_/B vssd1 vssd1 vccd1 vccd1 _18474_/B sky130_fd_sc_hd__nor2_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _11905_/A vssd1 vssd1 vccd1 vccd1 _11905_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _15673_/A _15673_/B _15673_/C vssd1 vssd1 vccd1 vccd1 _15677_/B sky130_fd_sc_hd__nand3_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output110_A _14343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ _16157_/C _20452_/C vssd1 vssd1 vccd1 vccd1 _12886_/A sky130_fd_sc_hd__nand2_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18176__A _18279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17412_ _12234_/X _12237_/X _15355_/A _15355_/B vssd1 vssd1 vccd1 vccd1 _17412_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14624_/A vssd1 vssd1 vccd1 vccd1 _15188_/A sky130_fd_sc_hd__buf_2
X_18392_ _18397_/B vssd1 vssd1 vccd1 vccd1 _18559_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _11837_/B _12084_/A _11831_/C vssd1 vssd1 vccd1 vccd1 _12246_/A sky130_fd_sc_hd__a21bo_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21297__B1_N _21423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17198_/X _17197_/Y _17193_/Y _17186_/X vssd1 vssd1 vccd1 vccd1 _17350_/A
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_14_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14555_ _14843_/A _14552_/X _14843_/B vssd1 vssd1 vccd1 vccd1 _14555_/X sky130_fd_sc_hd__o21a_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _18319_/A _11772_/A _18319_/B vssd1 vssd1 vccd1 vccd1 _12127_/A sky130_fd_sc_hd__a21o_1
XFILLER_158_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13506_ _13506_/A _13506_/B _13506_/C vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__nor3_4
X_17274_ _17120_/B _17116_/B _17116_/A vssd1 vssd1 vccd1 vccd1 _17464_/B sky130_fd_sc_hd__a21bo_2
XFILLER_147_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14486_ _14486_/A vssd1 vssd1 vccd1 vccd1 _14626_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__19719__B _19719_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22426__A _22426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11698_ _11698_/A _11698_/B _11698_/C vssd1 vssd1 vccd1 vccd1 _11698_/X sky130_fd_sc_hd__and3_1
X_19013_ _19504_/A _19013_/B _19013_/C vssd1 vssd1 vccd1 vccd1 _19013_/X sky130_fd_sc_hd__and3_1
X_16225_ _16225_/A vssd1 vssd1 vccd1 vccd1 _16225_/X sky130_fd_sc_hd__clkbuf_4
X_13437_ _13428_/A _13428_/B _21383_/A _13361_/X vssd1 vssd1 vccd1 vccd1 _13437_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17107__B1 _16944_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12952__A _16772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15966__C _17039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16156_ _15936_/A _20429_/B _16107_/X vssd1 vssd1 vccd1 vccd1 _16157_/A sky130_fd_sc_hd__o21ai_1
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20111__C1 _20593_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13368_ _13370_/A vssd1 vssd1 vccd1 vccd1 _13572_/A sky130_fd_sc_hd__buf_2
XANTENNA__13931__A3 _14765_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11568__A _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ _15107_/A _15107_/B _15107_/C vssd1 vssd1 vccd1 vccd1 _15112_/A sky130_fd_sc_hd__and3_1
X_12319_ _12368_/D vssd1 vssd1 vccd1 vccd1 _12319_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_181_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16087_ _16072_/X _16084_/Y _16085_/Y _16086_/Y vssd1 vssd1 vccd1 vccd1 _16090_/A
+ sky130_fd_sc_hd__o211a_1
X_13299_ _21495_/A _21588_/B _13311_/C vssd1 vssd1 vccd1 vccd1 _13300_/B sky130_fd_sc_hd__nand3_1
XFILLER_47_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19915_ _19861_/Y _19859_/Y _19860_/Y vssd1 vssd1 vccd1 vccd1 _19916_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__14341__B1 _14337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ _15098_/A _15047_/C vssd1 vssd1 vccd1 vccd1 _15040_/A sky130_fd_sc_hd__nand2_2
XANTENNA__19454__B _19896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19846_ _19985_/C _19846_/B _19846_/C _19901_/A vssd1 vssd1 vccd1 vccd1 _19850_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19173__C _19358_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20965__B2 _17928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16633__A2 _16630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19777_ _19848_/B _19783_/B _19781_/B vssd1 vssd1 vccd1 vccd1 _19837_/A sky130_fd_sc_hd__nand3_1
X_16989_ _16989_/A _16989_/B _16989_/C vssd1 vssd1 vccd1 vccd1 _17027_/B sky130_fd_sc_hd__nand3_2
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12104__C1 _12098_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15841__B1 _12765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19470__A _19792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18728_ _18522_/Y _18916_/B _18726_/Y _18727_/X vssd1 vssd1 vccd1 vccd1 _18729_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18386__A2 _18387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18659_ _18865_/A _18659_/B _19507_/D _18659_/D vssd1 vssd1 vccd1 vccd1 _18661_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21670_ _21689_/A _13162_/C _13162_/A _21669_/Y vssd1 vssd1 vccd1 vccd1 _21677_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_52_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22954__CLK _22959_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20621_ _20621_/A _20621_/B vssd1 vssd1 vccd1 vccd1 _20626_/A sky130_fd_sc_hd__nand2_1
XFILLER_178_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18814__A _18814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20552_ _20195_/Y _20065_/Y _20189_/B _20189_/C vssd1 vssd1 vccd1 vccd1 _20554_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__21878__C _21878_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_968 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20483_ _12832_/Y _20481_/Y _20593_/D _20482_/Y _20678_/A vssd1 vssd1 vccd1 vccd1
+ _20499_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_121_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22222_ _22304_/A _22223_/A _22308_/A vssd1 vssd1 vccd1 vccd1 _22222_/X sky130_fd_sc_hd__and3_1
XFILLER_118_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22153_ _22151_/X _22153_/B vssd1 vssd1 vccd1 vccd1 _22154_/A sky130_fd_sc_hd__and2b_1
XANTENNA__16321__A1 _16435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11909__C _11909_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21104_ _21102_/Y _21104_/B vssd1 vssd1 vccd1 vccd1 _21106_/A sky130_fd_sc_hd__and2b_1
X_22084_ _22084_/A vssd1 vssd1 vccd1 vccd1 _22084_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13693__A _14199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21035_ _21037_/D _21037_/A _21032_/Y _21034_/Y vssd1 vssd1 vccd1 vccd1 _21039_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_102_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11697__A1 _11693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_654 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20708__A1 _20110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11644__C _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21415__A _21415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21937_ _21937_/A vssd1 vssd1 vccd1 vccd1 _22182_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15413__A _20092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14399__B1 _14370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12758_/A vssd1 vssd1 vccd1 vccd1 _12968_/B sky130_fd_sc_hd__buf_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21868_ _21868_/A _21940_/A vssd1 vssd1 vccd1 vccd1 _21972_/A sky130_fd_sc_hd__nand2_2
XANTENNA__15060__A1 _14818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11660__B _15435_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11621_ _18328_/C _12154_/C _18328_/B vssd1 vssd1 vccd1 vccd1 _18133_/A sky130_fd_sc_hd__nand3_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20819_ _20812_/Y _20816_/Y _20818_/X vssd1 vssd1 vccd1 vccd1 _20822_/B sky130_fd_sc_hd__a21o_1
X_21799_ _21799_/A _21799_/B vssd1 vssd1 vccd1 vccd1 _21803_/A sky130_fd_sc_hd__nand2_1
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14340_ _11430_/C _14338_/X _14339_/X _14334_/X _13815_/X vssd1 vssd1 vccd1 vccd1
+ _14340_/X sky130_fd_sc_hd__a32o_1
XANTENNA__21684__A2 _22229_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ _11552_/A _11552_/B vssd1 vssd1 vccd1 vccd1 _11553_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14271_ _14231_/A _14231_/B _14575_/B _14861_/C _14212_/D vssd1 vssd1 vccd1 vccd1
+ _14272_/D sky130_fd_sc_hd__a32o_1
X_11483_ _12148_/A _11764_/B _12146_/A vssd1 vssd1 vccd1 vccd1 _11615_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12772__A _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16010_ _16010_/A _16010_/B vssd1 vssd1 vccd1 vccd1 _16012_/A sky130_fd_sc_hd__nand2_1
XANTENNA_input71_A x[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13222_ _13475_/C _13475_/A _13475_/B vssd1 vssd1 vccd1 vccd1 _13396_/B sky130_fd_sc_hd__a21bo_1
XFILLER_136_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20644__B1 _20631_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13153_ _21495_/B vssd1 vssd1 vccd1 vccd1 _21212_/C sky130_fd_sc_hd__buf_2
XFILLER_83_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12104_ _11381_/X _11731_/A _11702_/X _12096_/Y _12098_/Y vssd1 vssd1 vccd1 vccd1
+ _12110_/B sky130_fd_sc_hd__o221ai_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ _17907_/A _17907_/B _17958_/B _17920_/Y vssd1 vssd1 vccd1 vccd1 _17961_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__16863__A2 _16853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13084_ _22842_/Q vssd1 vssd1 vccd1 vccd1 _21476_/C sky130_fd_sc_hd__buf_2
XFILLER_3_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14699__A _22764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_610 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19700_ _19697_/D _19697_/B _19699_/X vssd1 vssd1 vccd1 vccd1 _19703_/A sky130_fd_sc_hd__a21o_1
XFILLER_151_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16912_ _16912_/A _20608_/B _20608_/C vssd1 vssd1 vccd1 vccd1 _17110_/A sky130_fd_sc_hd__nand3_2
X_12035_ _12035_/A _12035_/B vssd1 vssd1 vccd1 vccd1 _12035_/Y sky130_fd_sc_hd__nand2_1
X_17892_ _17890_/A _17890_/B _17891_/A vssd1 vssd1 vccd1 vccd1 _17893_/B sky130_fd_sc_hd__a21o_1
XANTENNA__21309__B _21476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22827__CLK _22929_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19631_ _19634_/C _19724_/A vssd1 vssd1 vccd1 vccd1 _19631_/Y sky130_fd_sc_hd__nand2_1
X_16843_ _16843_/A _16843_/B vssd1 vssd1 vccd1 vccd1 _16843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19562_ _19419_/X _19418_/X _19555_/A vssd1 vssd1 vccd1 vccd1 _19562_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_168_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16774_ _12571_/A _12571_/B _15538_/X _15541_/X vssd1 vssd1 vccd1 vccd1 _16774_/X
+ sky130_fd_sc_hd__a22o_1
X_13986_ _13986_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18513_ _18508_/Y _18511_/Y _18512_/X vssd1 vssd1 vccd1 vccd1 _18526_/A sky130_fd_sc_hd__o21bai_2
XFILLER_19_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15725_ _12378_/B _15631_/X _15991_/D _19154_/C _20870_/A vssd1 vssd1 vccd1 vccd1
+ _15725_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_20_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19493_ _17381_/A _17380_/A _19490_/D _19490_/C _19351_/B vssd1 vssd1 vccd1 vccd1
+ _19500_/A sky130_fd_sc_hd__o2111ai_4
X_12937_ _12937_/A _12958_/C vssd1 vssd1 vccd1 vccd1 _12937_/Y sky130_fd_sc_hd__nand2_1
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12947__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18444_ _18443_/Y _18406_/Y _18399_/Y vssd1 vssd1 vccd1 vccd1 _18564_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__15323__A _17532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15656_ _15621_/X _15630_/X _15652_/X _15653_/Y vssd1 vssd1 vccd1 vccd1 _15662_/A
+ sky130_fd_sc_hd__o22ai_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21044__B _21044_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17241__C _20928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12868_ _12868_/A vssd1 vssd1 vccd1 vccd1 _12868_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15051__B2 _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14607_ _14611_/A _14607_/B vssd1 vssd1 vccd1 vccd1 _14607_/Y sky130_fd_sc_hd__nand2_1
X_11819_ _11819_/A vssd1 vssd1 vccd1 vccd1 _11820_/A sky130_fd_sc_hd__clkbuf_4
X_18375_ _18387_/A _18387_/B _18387_/C vssd1 vssd1 vccd1 vccd1 _18396_/B sky130_fd_sc_hd__nand3_1
XFILLER_15_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15587_ _15587_/A vssd1 vssd1 vccd1 vccd1 _16530_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12526_/X _20508_/A _16498_/A _12540_/X vssd1 vssd1 vccd1 vccd1 _12799_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_762 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17326_ _17333_/C _17333_/D vssd1 vssd1 vccd1 vccd1 _17472_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17879__A1 _17731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14538_ _14099_/B _14096_/C _14099_/C vssd1 vssd1 vccd1 vccd1 _14538_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__17879__B2 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257_ _17257_/A _17257_/B vssd1 vssd1 vccd1 vccd1 _17260_/B sky130_fd_sc_hd__nand2_1
X_14469_ _13986_/B _14568_/A _14143_/X _14467_/X _14468_/Y vssd1 vssd1 vccd1 vccd1
+ _14472_/B sky130_fd_sc_hd__o221ai_1
XFILLER_88_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19168__C _19168_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15696__C _15997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16208_ _16208_/A _16402_/B vssd1 vssd1 vccd1 vccd1 _16210_/C sky130_fd_sc_hd__nand2_1
XFILLER_146_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12168__A2 _15887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17188_ _17188_/A _17188_/B vssd1 vssd1 vccd1 vccd1 _17188_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11298__A _22786_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ _16169_/A _16169_/B _16174_/A vssd1 vssd1 vccd1 vccd1 _16143_/C sky130_fd_sc_hd__and3_1
XFILLER_6_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18056__A1 _22905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21219__B _21944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19829_ _19890_/A _19890_/B _19891_/A _19891_/D vssd1 vssd1 vccd1 vccd1 _19831_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_624 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14617__A1 _15058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22840_ _22933_/CLK _22852_/Q vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18359__A2 _16921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22771_ _22771_/CLK _22771_/D vssd1 vssd1 vccd1 vccd1 _22771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15233__A _15233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11851__A1 _15978_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21722_ _21801_/A _21801_/B vssd1 vssd1 vccd1 vccd1 _21799_/B sky130_fd_sc_hd__xnor2_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11851__B2 _12050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20571__C1 _17401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12575__A2_N _20101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21653_ _21658_/A _21658_/B _21658_/C _21652_/Y vssd1 vssd1 vccd1 vccd1 _21653_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20793__B _20793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20604_ _20482_/Y _20486_/X _20479_/Y vssd1 vssd1 vccd1 vccd1 _20613_/A sky130_fd_sc_hd__a21oi_1
XFILLER_149_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21584_ _21584_/A _22734_/Q _21584_/C vssd1 vssd1 vccd1 vccd1 _21588_/C sky130_fd_sc_hd__nand3_1
XFILLER_166_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20535_ _20531_/B _20535_/B _20535_/C vssd1 vssd1 vccd1 vccd1 _20538_/B sky130_fd_sc_hd__nand3b_1
XFILLER_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12159__A2 _12158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22615__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13356__B2 _13166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20466_ _20582_/A _20466_/B _20582_/C vssd1 vssd1 vccd1 vccd1 _20495_/B sky130_fd_sc_hd__and3_1
XFILLER_174_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18295__A1 _18636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22205_ _21700_/X _21701_/X _22212_/A _22212_/B _22258_/B vssd1 vssd1 vccd1 vccd1
+ _22206_/C sky130_fd_sc_hd__o221ai_4
XFILLER_145_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17100__A1_N _17310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20397_ _20397_/A _20397_/B vssd1 vssd1 vccd1 vccd1 _20397_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22136_ _22196_/A _22196_/B _22137_/C _22137_/D vssd1 vssd1 vccd1 vccd1 _22138_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22067_ _22131_/A _22131_/B _22132_/B _22135_/A vssd1 vssd1 vccd1 vccd1 _22068_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21018_ _21044_/C _21018_/B vssd1 vssd1 vccd1 vccd1 _21020_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__19795__A1 _17421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19822__B _22921_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15805__B1 _15298_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13840_ _22760_/Q vssd1 vssd1 vccd1 vccd1 _13892_/B sky130_fd_sc_hd__inv_2
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13771_ _22872_/Q vssd1 vssd1 vccd1 vccd1 _14502_/A sky130_fd_sc_hd__inv_2
X_22969_ input67/X vssd1 vssd1 vccd1 vccd1 _22969_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15510_ _15756_/B _15510_/B _15510_/C vssd1 vssd1 vccd1 vccd1 _15738_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__11671__A _16257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15143__A _15175_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12722_ _12716_/X _12718_/X _12968_/D _12721_/X _12682_/X vssd1 vssd1 vccd1 vccd1
+ _12933_/D sky130_fd_sc_hd__o221ai_4
X_16490_ _12772_/A _12774_/A _16225_/A _16227_/A _17251_/A vssd1 vssd1 vccd1 vccd1
+ _16494_/A sky130_fd_sc_hd__o221ai_4
XFILLER_128_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15441_ _17234_/A vssd1 vssd1 vccd1 vccd1 _18197_/C sky130_fd_sc_hd__buf_4
XFILLER_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _16498_/D vssd1 vssd1 vccd1 vccd1 _16067_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_169_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15584__A2 _14430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_790 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _11627_/A vssd1 vssd1 vccd1 vccd1 _18328_/A sky130_fd_sc_hd__buf_2
X_18160_ _18383_/A _18383_/B _18155_/Y _18159_/X vssd1 vssd1 vccd1 vccd1 _18163_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15372_ _20456_/B vssd1 vssd1 vccd1 vccd1 _20593_/B sky130_fd_sc_hd__buf_2
XFILLER_8_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12584_ _12584_/A _12630_/B vssd1 vssd1 vccd1 vccd1 _12584_/Y sky130_fd_sc_hd__nand2_1
X_17111_ _17111_/A vssd1 vssd1 vccd1 vccd1 _17732_/A sky130_fd_sc_hd__buf_2
XFILLER_129_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14323_ _18953_/C _14317_/X _14320_/X _14322_/X _14220_/D vssd1 vssd1 vccd1 vccd1
+ _14323_/X sky130_fd_sc_hd__a32o_2
XFILLER_156_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18091_ _11738_/X _11737_/X _15458_/A _18093_/A _18093_/B vssd1 vssd1 vccd1 vccd1
+ _18091_/Y sky130_fd_sc_hd__o2111ai_4
X_11535_ _11578_/A _11581_/A _11542_/A _11541_/A _11529_/Y vssd1 vssd1 vccd1 vccd1
+ _11536_/C sky130_fd_sc_hd__o221ai_1
XFILLER_183_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15336__A2 _15718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17042_ _17042_/A vssd1 vssd1 vccd1 vccd1 _17042_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22606__A1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14254_ _14220_/D _15154_/B _14226_/A _14250_/Y _14253_/Y vssd1 vssd1 vccd1 vccd1
+ _14254_/X sky130_fd_sc_hd__a32o_1
XFILLER_125_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11466_ _11324_/X _11325_/A _11311_/Y _11988_/A vssd1 vssd1 vccd1 vccd1 _15776_/B
+ sky130_fd_sc_hd__a31o_4
XANTENNA__11358__B1 _11334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13205_ _22721_/Q vssd1 vssd1 vccd1 vccd1 _13234_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1011 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11397_ _11968_/B vssd1 vssd1 vccd1 vccd1 _18876_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_99_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14185_ _13930_/A _13930_/B _14181_/Y _14259_/A _14074_/A vssd1 vssd1 vccd1 vccd1
+ _14185_/X sky130_fd_sc_hd__a221o_2
XFILLER_139_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16297__B1 _15981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16836__A2 _20806_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ _13105_/Y _13180_/B _13120_/Y vssd1 vssd1 vccd1 vccd1 _13136_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _18980_/X _18982_/X _19185_/A _19187_/C vssd1 vssd1 vccd1 vccd1 _19086_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11846__A _12003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17944_ _17891_/B _17891_/A _17896_/A vssd1 vssd1 vccd1 vccd1 _17945_/B sky130_fd_sc_hd__o21a_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13067_ _13067_/A _13067_/B _21469_/B _13112_/C vssd1 vssd1 vccd1 vccd1 _21188_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_140_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12018_ _12018_/A vssd1 vssd1 vccd1 vccd1 _12018_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17875_ _17875_/A vssd1 vssd1 vccd1 vccd1 _21048_/C sky130_fd_sc_hd__buf_2
XFILLER_93_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18629__A _18629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17533__A _20870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19614_ _19614_/A _19614_/B _19614_/C vssd1 vssd1 vccd1 vccd1 _19615_/A sky130_fd_sc_hd__and3_2
XFILLER_66_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16826_ _16451_/B _16825_/X _16452_/X vssd1 vssd1 vccd1 vccd1 _16831_/C sky130_fd_sc_hd__o21ai_2
XFILLER_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11284__C _11860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19545_ _19545_/A _19545_/B _19545_/C vssd1 vssd1 vccd1 vccd1 _19545_/Y sky130_fd_sc_hd__nand3_2
X_16757_ _16541_/X _16546_/Y _16521_/Y vssd1 vssd1 vccd1 vccd1 _16906_/A sky130_fd_sc_hd__o21ai_1
XFILLER_59_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13969_ _13904_/Y _14073_/A _13968_/Y vssd1 vssd1 vccd1 vccd1 _14002_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12677__A _16932_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15708_ _15397_/Y _15513_/Y _15700_/C _15706_/A vssd1 vssd1 vccd1 vccd1 _15709_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14595__C _15056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16688_ _16424_/Y _16667_/A _16686_/Y vssd1 vssd1 vccd1 vccd1 _16690_/A sky130_fd_sc_hd__a21o_1
X_19476_ _19476_/A _19476_/B _19476_/C vssd1 vssd1 vccd1 vccd1 _19476_/X sky130_fd_sc_hd__and3_1
XFILLER_34_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15024__A1 _15213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18427_ _12241_/B _12241_/A _18227_/X _18229_/X vssd1 vssd1 vccd1 vccd1 _18427_/X
+ sky130_fd_sc_hd__o2bb2a_2
X_15639_ _15333_/Y _15638_/X _15632_/Y _15319_/B vssd1 vssd1 vccd1 vccd1 _15639_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__15988__A _15988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14892__A _14892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18358_ _18156_/A _12111_/A _18093_/Y vssd1 vssd1 vccd1 vccd1 _18367_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__20305__C1 _20314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21304__A_N _13112_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19171__C1 _19170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_760 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17309_ _17334_/B vssd1 vssd1 vccd1 vccd1 _17486_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20856__B1 _20913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18289_ _12116_/A _16248_/X _18200_/Y vssd1 vssd1 vccd1 vccd1 _18289_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__15327__A2 _15326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20320_ _20293_/A _20293_/B _20298_/A _20298_/B vssd1 vssd1 vccd1 vccd1 _20320_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_190_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20251_ _20096_/Y _20250_/X _20110_/Y vssd1 vssd1 vccd1 vccd1 _20251_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__20084__A1 _12734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20182_ _20182_/A _20182_/B vssd1 vssd1 vccd1 vccd1 _20183_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14489__D _15006_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17443__A _17443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14786__B _14786_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18258__B _18258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22823_ _22929_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 _22823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16059__A _16059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22754_ _22791_/CLK _22754_/D vssd1 vssd1 vccd1 vccd1 _22754_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21705_ _21704_/C _21704_/A _22676_/Q vssd1 vssd1 vccd1 vccd1 _21832_/A sky130_fd_sc_hd__a21o_1
XFILLER_80_682 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22685_ _22943_/CLK _22685_/D vssd1 vssd1 vccd1 vccd1 _22685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15113__D _15154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21636_ _21654_/A _21654_/B vssd1 vssd1 vccd1 vccd1 _21636_/X sky130_fd_sc_hd__and2_1
XFILLER_139_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19162__C1 _16554_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15318__A2 _11988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21567_ _21574_/A _21820_/A _21707_/B vssd1 vssd1 vccd1 vccd1 _21568_/C sky130_fd_sc_hd__a21o_1
XANTENNA__17712__B1 _17502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22672__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13211__A _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11320_ _11790_/C vssd1 vssd1 vccd1 vccd1 _18338_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20518_ _20519_/A _20519_/B _20519_/C vssd1 vssd1 vccd1 vccd1 _20623_/A sky130_fd_sc_hd__a21oi_2
X_21498_ _21850_/A _21498_/B _21615_/A _21498_/D vssd1 vssd1 vccd1 vccd1 _21640_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_180_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20449_ _20449_/A _20449_/B _20449_/C vssd1 vssd1 vccd1 vccd1 _20449_/Y sky130_fd_sc_hd__nor3_2
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20075__A1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11666__A _16257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22119_ _22119_/A _22119_/B _22119_/C vssd1 vssd1 vccd1 vccd1 _22128_/A sky130_fd_sc_hd__nand3_1
XFILLER_95_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15990_ _12273_/B _16324_/C _12279_/B _11911_/A vssd1 vssd1 vccd1 vccd1 _16129_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_125_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input34_A wb_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ _15056_/A _15056_/B _15004_/D _15010_/A _14953_/A vssd1 vssd1 vccd1 vccd1
+ _14945_/C sky130_fd_sc_hd__a32o_1
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21575__A1 _21551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17660_ _17660_/A _17660_/B vssd1 vssd1 vccd1 vccd1 _17662_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14872_ _14872_/A _14932_/A vssd1 vssd1 vccd1 vccd1 _14872_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16611_ _16611_/A vssd1 vssd1 vccd1 vccd1 _17435_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__18991__A2 _19313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ _13820_/A _13845_/B _13799_/X vssd1 vssd1 vccd1 vccd1 _13823_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_169_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17591_ _17591_/A _17591_/B _20936_/C _19482_/A vssd1 vssd1 vccd1 vccd1 _17591_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16542_ _16530_/C _16231_/X _16509_/Y _16489_/X vssd1 vssd1 vccd1 vccd1 _16542_/Y
+ sky130_fd_sc_hd__a22oi_2
X_19330_ _19330_/A _19330_/B _19330_/C vssd1 vssd1 vccd1 vccd1 _19512_/A sky130_fd_sc_hd__nand3_4
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13754_ _13975_/D vssd1 vssd1 vccd1 vccd1 _13968_/C sky130_fd_sc_hd__buf_2
XFILLER_44_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19261_ _19251_/Y _19248_/Y _19249_/Y vssd1 vssd1 vccd1 vccd1 _19261_/Y sky130_fd_sc_hd__a21oi_2
X_12705_ _12968_/A _12716_/A _12967_/A _12727_/A vssd1 vssd1 vccd1 vccd1 _12705_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16473_ _16473_/A _16473_/B _17141_/A vssd1 vssd1 vccd1 vccd1 _16782_/A sky130_fd_sc_hd__nand3_1
XFILLER_31_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13685_ _21424_/A _21285_/C vssd1 vssd1 vccd1 vccd1 _21426_/A sky130_fd_sc_hd__nand2_1
X_18212_ _18212_/A _18277_/A _18276_/B vssd1 vssd1 vccd1 vccd1 _18232_/C sky130_fd_sc_hd__nand3_1
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15424_ _15403_/X _15731_/B _15423_/Y vssd1 vssd1 vccd1 vccd1 _15430_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__13568__A1 _21741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18615__C _19353_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19192_ _19010_/X _19237_/B _19237_/C _19237_/D vssd1 vssd1 vccd1 vccd1 _19192_/Y
+ sky130_fd_sc_hd__a22oi_4
X_12636_ _20675_/C vssd1 vssd1 vccd1 vccd1 _20972_/D sky130_fd_sc_hd__buf_2
XFILLER_15_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18143_ _11541_/A _12167_/X _18150_/A vssd1 vssd1 vccd1 vccd1 _18146_/A sky130_fd_sc_hd__o21ai_1
XFILLER_8_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15355_ _15355_/A _15355_/B vssd1 vssd1 vccd1 vccd1 _20477_/A sky130_fd_sc_hd__nand2_2
XFILLER_8_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12567_ _12567_/A vssd1 vssd1 vccd1 vccd1 _15299_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_129_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20302__A2 _12894_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14306_ _22586_/D input26/X _14310_/A vssd1 vssd1 vccd1 vccd1 _22369_/D sky130_fd_sc_hd__nor3b_2
X_18074_ _18075_/B _18082_/B _22907_/Q vssd1 vssd1 vccd1 vccd1 _18080_/A sky130_fd_sc_hd__a21bo_1
X_11518_ _18348_/A vssd1 vssd1 vccd1 vccd1 _15624_/A sky130_fd_sc_hd__buf_4
X_15286_ _22883_/Q _15286_/B vssd1 vssd1 vccd1 vccd1 _22871_/D sky130_fd_sc_hd__xor2_1
X_12498_ _12704_/A vssd1 vssd1 vccd1 vccd1 _15455_/A sky130_fd_sc_hd__buf_2
XFILLER_89_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17025_ _17025_/A _17025_/B _17025_/C vssd1 vssd1 vccd1 vccd1 _17025_/X sky130_fd_sc_hd__and3_1
XFILLER_109_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14237_ _14237_/A _14237_/B _14237_/C vssd1 vssd1 vccd1 vccd1 _14237_/X sky130_fd_sc_hd__and3_1
X_11449_ _11720_/A _11438_/B _15435_/B vssd1 vssd1 vccd1 vccd1 _11778_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__22055__A2 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20066__A1 _13041_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ _14165_/X _14166_/Y _14089_/Y _14167_/X vssd1 vssd1 vccd1 vccd1 _14172_/B
+ sky130_fd_sc_hd__o22ai_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13119_ _21448_/A _13168_/C vssd1 vssd1 vccd1 vccd1 _13120_/A sky130_fd_sc_hd__nand2_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _18935_/A _18932_/Y _18938_/Y _18937_/Y vssd1 vssd1 vccd1 vccd1 _19122_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _14099_/A _14099_/B _14099_/C vssd1 vssd1 vccd1 vccd1 _14099_/Y sky130_fd_sc_hd__nand3_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11295__B _11295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _17927_/A vssd1 vssd1 vccd1 vccd1 _19899_/B sky130_fd_sc_hd__clkbuf_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20369__A2 _20611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17858_ _17858_/A vssd1 vssd1 vccd1 vccd1 _17858_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18982__A2 _18889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16809_ _19461_/A _16809_/B _17133_/A _19317_/D vssd1 vssd1 vccd1 vccd1 _16810_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13256__B1 _21584_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17789_ _17507_/A _17726_/Y _17788_/X _17959_/C vssd1 vssd1 vccd1 vccd1 _17793_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16993__A1 _11904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19528_ _19528_/A _19528_/B _19528_/C vssd1 vssd1 vccd1 vccd1 _19529_/A sky130_fd_sc_hd__nand3_1
XANTENNA__11806__A1 _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19459_ _19390_/Y _19458_/Y _19392_/B vssd1 vssd1 vccd1 vccd1 _19528_/A sky130_fd_sc_hd__o21ai_1
XFILLER_179_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22470_ _22470_/A vssd1 vssd1 vccd1 vccd1 _22731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20129__A _20129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21421_ _21421_/A vssd1 vssd1 vccd1 vccd1 _21560_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21352_ _21496_/A vssd1 vssd1 vccd1 vccd1 _21352_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20303_ _20442_/A _20444_/A _20442_/B vssd1 vssd1 vccd1 vccd1 _20553_/A sky130_fd_sc_hd__nand3_4
XFILLER_163_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21283_ _21422_/B vssd1 vssd1 vccd1 vccd1 _21424_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20234_ _20234_/A vssd1 vssd1 vccd1 vccd1 _20397_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13685__B _21285_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20165_ _20165_/A _20165_/B _20165_/C vssd1 vssd1 vccd1 vccd1 _20165_/Y sky130_fd_sc_hd__nand3_2
XFILLER_162_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11917__C _18629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20096_ _20096_/A _20096_/B vssd1 vssd1 vccd1 vccd1 _20096_/Y sky130_fd_sc_hd__nand2_2
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15405__B _15776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15787__A2 _12689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22806_ _22807_/CLK _22806_/D vssd1 vssd1 vccd1 vccd1 _22806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15251__A4 _15205_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ _20999_/A _20999_/B _22939_/Q vssd1 vssd1 vccd1 vccd1 _21076_/A sky130_fd_sc_hd__a21o_1
XANTENNA__18716__B _19358_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21423__A _21423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22737_ _22768_/CLK _22737_/D vssd1 vssd1 vccd1 vccd1 _22737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _13470_/A vssd1 vssd1 vccd1 vccd1 _13470_/Y sky130_fd_sc_hd__inv_2
X_22668_ _22964_/CLK _22668_/D vssd1 vssd1 vccd1 vccd1 _22668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ _12421_/A _12822_/A _16319_/C _12550_/A vssd1 vssd1 vccd1 vccd1 _15326_/A
+ sky130_fd_sc_hd__and4_2
XANTENNA__18489__A1 _12009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21619_ _21508_/A _21508_/B _21485_/A vssd1 vssd1 vccd1 vccd1 _21624_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__19686__B1 _17391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22599_ _22656_/S vssd1 vssd1 vccd1 vccd1 _22608_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_166_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15140_ _15097_/A _15100_/A _15139_/Y vssd1 vssd1 vccd1 vccd1 _15173_/B sky130_fd_sc_hd__a21boi_1
X_12352_ _12341_/A _12324_/X _12361_/A vssd1 vssd1 vccd1 vccd1 _12802_/A sky130_fd_sc_hd__a21o_1
XFILLER_138_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11981__B1 _11372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11303_ _22784_/Q _22785_/Q vssd1 vssd1 vccd1 vccd1 _11764_/A sky130_fd_sc_hd__nor2_1
X_15071_ _15154_/A _15154_/B _15152_/A _15186_/A _15080_/A vssd1 vssd1 vccd1 vccd1
+ _15073_/A sky130_fd_sc_hd__a41o_1
X_12283_ _22693_/Q _22692_/Q _22691_/Q vssd1 vssd1 vccd1 vccd1 _12284_/A sky130_fd_sc_hd__nor3_1
XFILLER_5_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13183__C1 _21473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14022_ _14022_/A _14022_/B _14022_/C vssd1 vssd1 vccd1 vccd1 _14052_/C sky130_fd_sc_hd__nand3_1
XFILLER_84_1022 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17067__B _22895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18830_ _18830_/A _18830_/B _18830_/C _18830_/D vssd1 vssd1 vccd1 vccd1 _18830_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_45_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15475__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14278__A2 _14834_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14203__C _14785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18761_ _18761_/A _18761_/B vssd1 vssd1 vccd1 vccd1 _18762_/C sky130_fd_sc_hd__nand2_1
X_15973_ _15972_/X _16100_/D _17312_/A _15900_/Y _16006_/B vssd1 vssd1 vccd1 vccd1
+ _15976_/A sky130_fd_sc_hd__a32oi_1
XFILLER_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17712_ _17708_/Y _17790_/C _17502_/X _17607_/X vssd1 vssd1 vccd1 vccd1 _17713_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14924_ _14924_/A _14982_/B vssd1 vssd1 vccd1 vccd1 _14927_/A sky130_fd_sc_hd__or2b_2
XANTENNA__21012__A3 _21048_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18692_ _18890_/A _18690_/Y _18691_/Y vssd1 vssd1 vccd1 vccd1 _18692_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__14500__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17643_ _17643_/A _18830_/D _19768_/D _20745_/C vssd1 vssd1 vccd1 vccd1 _17643_/X
+ sky130_fd_sc_hd__and4_1
X_14855_ _14942_/A _14854_/X _13904_/Y _14942_/B vssd1 vssd1 vccd1 vccd1 _14881_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_64_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13806_ _14118_/B vssd1 vssd1 vccd1 vccd1 _14270_/A sky130_fd_sc_hd__buf_2
X_17574_ _17574_/A _17574_/B _17574_/C vssd1 vssd1 vccd1 vccd1 _17575_/C sky130_fd_sc_hd__nand3_1
X_14786_ _14786_/A _14786_/B _14786_/C vssd1 vssd1 vccd1 vccd1 _14872_/A sky130_fd_sc_hd__nand3_1
X_11998_ _16241_/A _11988_/X _15893_/A _12135_/A _12135_/B vssd1 vssd1 vccd1 vccd1
+ _18508_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_63_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14450__A2 _11334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16525_ _16493_/A _16493_/B _16508_/X _16510_/Y _16524_/Y vssd1 vssd1 vccd1 vccd1
+ _16529_/B sky130_fd_sc_hd__o221ai_1
X_19313_ _19313_/A vssd1 vssd1 vccd1 vccd1 _19838_/A sky130_fd_sc_hd__clkbuf_4
X_13737_ _13750_/A vssd1 vssd1 vccd1 vccd1 _13737_/X sky130_fd_sc_hd__buf_2
XFILLER_44_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16727__A1 _11295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16727__B2 _16584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15331__A _15893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19244_ _19244_/A vssd1 vssd1 vccd1 vccd1 _19244_/Y sky130_fd_sc_hd__inv_2
X_16456_ _17129_/B vssd1 vssd1 vccd1 vccd1 _18797_/B sky130_fd_sc_hd__clkbuf_4
X_13668_ _13647_/A _13640_/B _13666_/X _13641_/Y vssd1 vssd1 vccd1 vccd1 _13668_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15407_ _15731_/B _15403_/X _15404_/X _15406_/X vssd1 vssd1 vccd1 vccd1 _15513_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19175_ _18158_/X _18995_/B _19171_/Y _19174_/Y vssd1 vssd1 vccd1 vccd1 _19190_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15050__B _15050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13946__D1 _15058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ _12619_/A vssd1 vssd1 vccd1 vccd1 _12745_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16387_ _15339_/B _15339_/C _15339_/A _15668_/X _16213_/Y vssd1 vssd1 vccd1 vccd1
+ _16388_/A sky130_fd_sc_hd__a311o_1
X_13599_ _13526_/X _13567_/Y _13598_/Y vssd1 vssd1 vccd1 vccd1 _13599_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_191_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18126_ _18126_/A _18841_/B _18677_/B vssd1 vssd1 vccd1 vccd1 _18129_/A sky130_fd_sc_hd__nand3_1
X_15338_ _15327_/Y _15333_/Y _16720_/C _15336_/Y _16809_/B vssd1 vssd1 vccd1 vccd1
+ _15339_/C sky130_fd_sc_hd__o2111ai_4
XANTENNA__13961__A1 _13833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18057_ _18057_/A _18057_/B vssd1 vssd1 vccd1 vccd1 _18058_/A sky130_fd_sc_hd__and2_1
X_15269_ _15269_/A vssd1 vssd1 vccd1 vccd1 _22687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15702__A2 _17525_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20039__A1 _18778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17008_ _17006_/B _17006_/C _15936_/X _17728_/A vssd1 vssd1 vccd1 vccd1 _17008_/Y
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_126_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12516__A2 _12525_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11724__B1 _19320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17455__A2 _17523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18652__A1 _15981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14113__C _14963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16663__B1 _22893_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18959_ _19138_/B _19138_/C vssd1 vssd1 vccd1 vccd1 _19279_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21970_ _21970_/A vssd1 vssd1 vccd1 vccd1 _21970_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1032 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20921_ _20782_/B _20854_/Y _20860_/B vssd1 vssd1 vccd1 vccd1 _20923_/A sky130_fd_sc_hd__o21ai_1
XFILLER_6_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20852_ _12671_/X _17444_/A _20782_/B _20787_/B vssd1 vssd1 vccd1 vccd1 _20864_/B
+ sky130_fd_sc_hd__o31a_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20783_ _20676_/B _20780_/Y _20913_/A _20782_/Y _17385_/C vssd1 vssd1 vccd1 vccd1
+ _20787_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22522_ _22522_/A vssd1 vssd1 vccd1 vccd1 _22754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22453_ _13161_/C input61/X _22453_/S vssd1 vssd1 vccd1 vccd1 _22454_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20278__A1 _12761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21404_ _21404_/A _21404_/B vssd1 vssd1 vccd1 vccd1 _21404_/Y sky130_fd_sc_hd__nand2_1
XFILLER_194_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13952__B2 _22872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22384_ _22384_/A vssd1 vssd1 vccd1 vccd1 _22693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18891__A1 _11636_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21335_ _21351_/B vssd1 vssd1 vccd1 vccd1 _21725_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21266_ _21266_/A _21266_/B vssd1 vssd1 vccd1 vccd1 _21266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20217_ _20217_/A vssd1 vssd1 vccd1 vccd1 _20457_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11647__C _11647_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21197_ _21202_/A _21301_/A vssd1 vssd1 vccd1 vccd1 _21197_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20450__A1 _20449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20148_ _12864_/B _12862_/B _12843_/X _12851_/Y vssd1 vssd1 vccd1 vccd1 _20150_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__17615__B _17719_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _12970_/A vssd1 vssd1 vccd1 vccd1 _15893_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__22860__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20079_ _20177_/A vssd1 vssd1 vccd1 vccd1 _20728_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20202__A1 _20115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18946__A2 _20012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11921_ _11922_/A _11922_/B _11922_/C vssd1 vssd1 vccd1 vccd1 _11923_/A sky130_fd_sc_hd__a21o_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17631__A _17631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14640_ _14515_/B _14515_/C _14515_/A vssd1 vssd1 vccd1 vccd1 _14640_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _11566_/X _11845_/X _11846_/Y _11851_/X vssd1 vssd1 vccd1 vccd1 _11922_/C
+ sky130_fd_sc_hd__o31ai_4
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14571_/A vssd1 vssd1 vccd1 vccd1 _14571_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_159_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16709__A1 _11904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ _11783_/A _18319_/B _11783_/C vssd1 vssd1 vccd1 vccd1 _12130_/A sky130_fd_sc_hd__nand3_1
XANTENNA__20505__A2 _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16310_ _16301_/Y _16305_/Y _16309_/Y vssd1 vssd1 vccd1 vccd1 _16310_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_25_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13522_ _13517_/X _13528_/A _13452_/A _13521_/Y vssd1 vssd1 vccd1 vccd1 _13523_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_17290_ _17290_/A _17290_/B _17290_/C vssd1 vssd1 vccd1 vccd1 _17464_/A sky130_fd_sc_hd__nand3_2
XFILLER_15_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17382__A1 _17380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16241_ _16241_/A _16481_/B _16241_/C _16241_/D vssd1 vssd1 vccd1 vccd1 _16241_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13453_ _21177_/A _21750_/C _13461_/B _13461_/A vssd1 vssd1 vccd1 vccd1 _13454_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_174_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15379__A1_N _15389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14990__A _15186_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19123__A2 _19113_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12404_ _12404_/A vssd1 vssd1 vccd1 vccd1 _16302_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16172_ _16124_/X _12876_/X _16122_/Y _16126_/Y vssd1 vssd1 vccd1 vccd1 _16172_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_103_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13384_ _13384_/A _13384_/B vssd1 vssd1 vccd1 vccd1 _13385_/D sky130_fd_sc_hd__nand2_1
XANTENNA__18331__B1 _15901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15123_ _15119_/D _15152_/A _15059_/Y _15113_/X vssd1 vssd1 vccd1 vccd1 _15123_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12335_ _12335_/A vssd1 vssd1 vccd1 vccd1 _16318_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18882__A1 _12009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19931_ _19970_/C _19970_/A _22923_/Q vssd1 vssd1 vccd1 vccd1 _19975_/A sky130_fd_sc_hd__a21oi_2
XFILLER_173_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15054_ _14998_/X _15001_/C _15052_/X vssd1 vssd1 vccd1 vccd1 _15128_/A sky130_fd_sc_hd__a21o_1
X_12266_ _22703_/Q vssd1 vssd1 vccd1 vccd1 _12303_/A sky130_fd_sc_hd__clkbuf_2
X_14005_ _13916_/Y _14021_/C _14021_/D vssd1 vssd1 vccd1 vccd1 _14006_/C sky130_fd_sc_hd__a21boi_1
XANTENNA__18634__A1 _18619_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17437__A2 _17440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19862_ _19859_/Y _19860_/Y _19861_/Y vssd1 vssd1 vccd1 vccd1 _19862_/X sky130_fd_sc_hd__o21a_1
XANTENNA__17806__A _20975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12197_ _22963_/Q vssd1 vssd1 vccd1 vccd1 _15486_/C sky130_fd_sc_hd__clkinv_2
XANTENNA__15448__A1 _18197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16645__B1 _16644_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15448__B2 _19694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput81 _22969_/X vssd1 vssd1 vccd1 vccd1 wb_ack_o sky130_fd_sc_hd__buf_2
X_18813_ _18828_/A _18830_/C _18812_/Y vssd1 vssd1 vccd1 vccd1 _18818_/A sky130_fd_sc_hd__a21o_1
XFILLER_150_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput92 _14395_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_110_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19793_ _19793_/A _19901_/C _19793_/C vssd1 vssd1 vccd1 vccd1 _19794_/C sky130_fd_sc_hd__and3_1
XANTENNA__17525__B _17739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13459__B1 _21621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11854__A _18810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15326__A _15326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14868__C _14868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14120__A1 _14122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18744_ _18933_/A _18933_/B vssd1 vssd1 vccd1 vccd1 _18744_/Y sky130_fd_sc_hd__nand2_1
X_15956_ _16034_/A _16210_/A _15955_/X vssd1 vssd1 vccd1 vccd1 _15957_/C sky130_fd_sc_hd__a21o_1
XFILLER_110_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14671__A2 _13930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ _14815_/C _14815_/B _14815_/A vssd1 vssd1 vccd1 vccd1 _14907_/Y sky130_fd_sc_hd__a21oi_1
X_15887_ _15887_/A vssd1 vssd1 vccd1 vccd1 _15887_/X sky130_fd_sc_hd__buf_4
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12682__A1 _12689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18675_ _22798_/Q vssd1 vssd1 vccd1 vccd1 _18841_/C sky130_fd_sc_hd__inv_2
XFILLER_37_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17626_ _17626_/A _17626_/B vssd1 vssd1 vccd1 vccd1 _17626_/X sky130_fd_sc_hd__or2_1
X_14838_ _14982_/A _14838_/B vssd1 vssd1 vccd1 vccd1 _14842_/A sky130_fd_sc_hd__nand2_2
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17557_ _17413_/Y _17414_/X _17410_/X vssd1 vssd1 vccd1 vccd1 _17557_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14769_ _14769_/A _14917_/B vssd1 vssd1 vccd1 vccd1 _14826_/A sky130_fd_sc_hd__xor2_1
XFILLER_189_451 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12685__A _16498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ _12716_/X _16758_/A _16506_/X _16507_/X _16496_/X vssd1 vssd1 vccd1 vccd1
+ _16508_/X sky130_fd_sc_hd__o221a_1
XFILLER_60_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17488_ _17483_/Y _17484_/X _17491_/C vssd1 vssd1 vccd1 vccd1 _17514_/A sky130_fd_sc_hd__o21bai_2
XFILLER_60_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19227_ _19227_/A _19227_/B _19227_/C vssd1 vssd1 vccd1 vccd1 _19227_/Y sky130_fd_sc_hd__nand3_1
XFILLER_165_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16439_ _16439_/A _16439_/B vssd1 vssd1 vccd1 vccd1 _16439_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16581__C1 _22702_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19114__A2 _18023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18803__C _19353_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19158_ _19155_/Y _19156_/Y _19185_/C _18990_/A vssd1 vssd1 vccd1 vccd1 _19386_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18322__B1 _19194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18109_ _18109_/A _18109_/B _18109_/C vssd1 vssd1 vccd1 vccd1 _18278_/A sky130_fd_sc_hd__nand3_4
XFILLER_173_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19089_ _19089_/A vssd1 vssd1 vccd1 vccd1 _19106_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16884__B1 _16880_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21120_ _21120_/A vssd1 vssd1 vccd1 vccd1 _21150_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__20680__A1 _17423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21051_ _21050_/C _21017_/A _21017_/B _21090_/A _21050_/B vssd1 vssd1 vccd1 vccd1
+ _21052_/B sky130_fd_sc_hd__a32o_1
XANTENNA__18625__A1 _19043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17428__A2 _15808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18625__B2 _18636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22883__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20002_ _19962_/A _19962_/B _19962_/C vssd1 vssd1 vccd1 vccd1 _20002_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_115_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14111__A1 _14112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19050__A1 _18371_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21953_ _21951_/Y _21952_/X _21758_/C _21882_/A vssd1 vssd1 vccd1 vccd1 _22064_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__12673__A1 _12968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12673__B2 _12719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ _20832_/Y _20902_/Y _20773_/B _20903_/Y vssd1 vssd1 vccd1 vccd1 _20905_/B
+ sky130_fd_sc_hd__a22oi_4
X_21884_ _21874_/C _21596_/B _21753_/B _21753_/C vssd1 vssd1 vccd1 vccd1 _21884_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20835_ _20835_/A vssd1 vssd1 vccd1 vccd1 _20835_/X sky130_fd_sc_hd__buf_2
XFILLER_168_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16067__A _19470_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21696__B1 _21838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20766_ _20776_/C _20776_/A _22935_/Q vssd1 vssd1 vccd1 vccd1 _20772_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22505_ _22505_/A vssd1 vssd1 vccd1 vccd1 _22747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15375__B1 _15367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20697_ _20697_/A _20697_/B _20697_/C vssd1 vssd1 vccd1 vccd1 _20697_/Y sky130_fd_sc_hd__nor3_1
XFILLER_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13925__A1 _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22436_ _22436_/A vssd1 vssd1 vccd1 vccd1 _22717_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__21420__B _21560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22367_ _22368_/A _22368_/B vssd1 vssd1 vccd1 vccd1 _22947_/D sky130_fd_sc_hd__nor2_1
XFILLER_136_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ _18208_/A _12123_/B _12115_/X _12119_/X vssd1 vssd1 vccd1 vccd1 _12189_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__20671__A1 _15940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21318_ _21318_/A vssd1 vssd1 vccd1 vccd1 _21958_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22298_ _22298_/A _22325_/B vssd1 vssd1 vccd1 vccd1 _22299_/A sky130_fd_sc_hd__and2_1
XFILLER_7_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ _11932_/C _11762_/B _11762_/A vssd1 vssd1 vccd1 vccd1 _12240_/B sky130_fd_sc_hd__a21boi_2
XANTENNA__14350__A1 _22761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14350__B2 _13304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21249_ _21249_/A _21249_/B vssd1 vssd1 vccd1 vccd1 _21251_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20974__A2 _21017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15810_ _15810_/A _15810_/B _15810_/C vssd1 vssd1 vccd1 vccd1 _15823_/A sky130_fd_sc_hd__and3_1
X_16790_ _16972_/A _16971_/A _16784_/X _16789_/X vssd1 vssd1 vccd1 vccd1 _16796_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15741_ _15864_/A _15709_/Y _15734_/X vssd1 vssd1 vccd1 vccd1 _15854_/A sky130_fd_sc_hd__a21o_1
XFILLER_86_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19041__A1 _18795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20187__B1 _13045_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12664__A1 _16160_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ _12981_/D _16100_/A _12981_/B _12941_/X vssd1 vssd1 vccd1 vccd1 _12954_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__19041__B2 _12116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_530 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _11904_/A vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__clkbuf_4
X_18460_ _12204_/X _17400_/X _17817_/A _11566_/X vssd1 vssd1 vccd1 vccd1 _18461_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ _15672_/A _15672_/B vssd1 vssd1 vccd1 vccd1 _15672_/Y sky130_fd_sc_hd__nand2_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12755_/B _12755_/C _12755_/A _12898_/B _12898_/C vssd1 vssd1 vccd1 vccd1
+ _12889_/B sky130_fd_sc_hd__a32oi_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16260__D1 _18848_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18176__B _18278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17411_ _17550_/A _17550_/B _17399_/Y _17410_/X vssd1 vssd1 vccd1 vccd1 _17416_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14623_ _14506_/Y _14612_/X _14892_/D _14614_/Y _14510_/A vssd1 vssd1 vccd1 vccd1
+ _14623_/X sky130_fd_sc_hd__o2111a_1
X_18391_ _18389_/X _18390_/X _18353_/Y _18356_/Y vssd1 vssd1 vccd1 vccd1 _18397_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _11696_/C _11692_/Y _12247_/C vssd1 vssd1 vccd1 vccd1 _11838_/A sky130_fd_sc_hd__o21ai_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14810__C1 _13823_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17341_/X _17338_/X _17330_/Y _17337_/X vssd1 vssd1 vccd1 vccd1 _17342_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14554_/A _14554_/B vssd1 vssd1 vccd1 vccd1 _14843_/B sky130_fd_sc_hd__xnor2_2
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _22792_/Q vssd1 vssd1 vccd1 vccd1 _18319_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13505_ _21351_/C _13370_/A _13579_/A _21212_/C vssd1 vssd1 vccd1 vccd1 _13506_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19288__A _22916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17273_ _17273_/A vssd1 vssd1 vccd1 vccd1 _17307_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14485_ _14684_/A _13968_/C _14684_/C _14484_/Y vssd1 vssd1 vccd1 vccd1 _14486_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18192__A _18192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11697_ _11693_/X _11565_/Y _12059_/B vssd1 vssd1 vccd1 vccd1 _12247_/C sky130_fd_sc_hd__o21ai_2
XFILLER_158_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16224_ _16242_/A _16242_/B vssd1 vssd1 vccd1 vccd1 _16225_/A sky130_fd_sc_hd__nand2_4
X_19012_ _19687_/D _19351_/A _19012_/C _19012_/D vssd1 vssd1 vccd1 vccd1 _19012_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_174_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13436_ _21522_/C _21498_/B _21522_/A _21739_/B vssd1 vssd1 vccd1 vccd1 _13436_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_127_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18304__B1 _18459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15966__D _17401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16155_ _16155_/A vssd1 vssd1 vccd1 vccd1 _20429_/B sky130_fd_sc_hd__clkbuf_2
X_13367_ _13423_/A _13434_/A _13366_/Y vssd1 vssd1 vccd1 vccd1 _13367_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_154_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _15086_/B _15078_/B _15078_/A vssd1 vssd1 vccd1 vccd1 _15132_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__20662__A1 _20548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12318_ _12428_/B vssd1 vssd1 vccd1 vccd1 _12596_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11568__B _11568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16086_ _16093_/A _16093_/B _16017_/X _15824_/C vssd1 vssd1 vccd1 vccd1 _16086_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_142_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13298_ _13302_/A _13295_/X _21188_/B _13097_/A vssd1 vssd1 vccd1 vccd1 _13311_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_170_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19914_ _19914_/A _19914_/B vssd1 vssd1 vccd1 vccd1 _19916_/A sky130_fd_sc_hd__nor2_2
XFILLER_170_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14341__A1 _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15037_ _15035_/A _15035_/B _15035_/C vssd1 vssd1 vccd1 vccd1 _15047_/C sky130_fd_sc_hd__a21o_1
X_12249_ _12249_/A _12249_/B vssd1 vssd1 vccd1 vccd1 _12251_/B sky130_fd_sc_hd__nand2_1
XANTENNA__20414__A1 _20843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19845_ _19844_/B _20012_/B _20012_/C _19900_/A _19844_/D vssd1 vssd1 vccd1 vccd1
+ _19846_/C sky130_fd_sc_hd__a32o_1
XFILLER_123_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20965__A2 _15941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15056__A _15056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19776_ _19699_/X _19697_/B _19697_/D vssd1 vssd1 vccd1 vccd1 _19781_/B sky130_fd_sc_hd__a21boi_1
XFILLER_7_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16988_ _16988_/A _16988_/B _17188_/A _17188_/B vssd1 vssd1 vccd1 vccd1 _16989_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12104__B1 _11702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15841__B2 _15840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18727_ _18915_/A _18526_/D _18916_/A vssd1 vssd1 vccd1 vccd1 _18727_/X sky130_fd_sc_hd__a21o_1
XANTENNA__19470__B _19470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15939_ _15939_/A vssd1 vssd1 vccd1 vccd1 _15940_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18658_ _18797_/C vssd1 vssd1 vccd1 vccd1 _19507_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_276 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17609_ _17226_/A _17227_/A _17853_/A _17507_/A vssd1 vssd1 vccd1 vccd1 _17713_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18589_ _18589_/A vssd1 vssd1 vccd1 vccd1 _19293_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_3_2_0_bq_clk_i_A clkbuf_3_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20620_ _20620_/A _20620_/B _20620_/C vssd1 vssd1 vccd1 vccd1 _20621_/B sky130_fd_sc_hd__nand3_1
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14119__B _14564_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20551_ _20445_/Y _20550_/Y _20547_/X vssd1 vssd1 vccd1 vccd1 _20551_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_177_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16615__A _16617_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18533__C _19317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20482_ _20482_/A _20482_/B vssd1 vssd1 vccd1 vccd1 _20482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22221_ _22221_/A _22221_/B _22221_/C vssd1 vssd1 vccd1 vccd1 _22308_/A sky130_fd_sc_hd__and3_1
XANTENNA__18846__A1 _11704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20102__B1 _20250_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18830__A _18830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22152_ _22290_/C _22290_/D _22290_/A _22290_/B _22094_/A vssd1 vssd1 vccd1 vccd1
+ _22153_/B sky130_fd_sc_hd__a221o_1
XFILLER_161_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22352__A _22352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14332__A1 _11860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21103_ _21122_/B _22942_/Q _21122_/A vssd1 vssd1 vccd1 vccd1 _21104_/B sky130_fd_sc_hd__nand3_1
XFILLER_161_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14332__B2 _12493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22083_ _22090_/A vssd1 vssd1 vccd1 vccd1 _22142_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21034_ _21067_/C vssd1 vssd1 vccd1 vccd1 _21034_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11697__A2 _11565_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11449__A2 _11438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17034__B1 _16740_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21936_ _21936_/A vssd1 vssd1 vccd1 vccd1 _22182_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_563 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21867_ _21876_/A _21877_/A _21938_/B vssd1 vssd1 vccd1 vccd1 _21940_/A sky130_fd_sc_hd__nand3_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11620_ _11974_/C vssd1 vssd1 vccd1 vccd1 _18328_/B sky130_fd_sc_hd__buf_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11660__C _16482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20818_ _20818_/A _20818_/B vssd1 vssd1 vccd1 vccd1 _20818_/X sky130_fd_sc_hd__or2_1
XFILLER_169_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21798_ _21899_/A _21802_/C vssd1 vssd1 vccd1 vccd1 _21799_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18534__B1 _17421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11551_ _11552_/A _11551_/B _11551_/C _11552_/B vssd1 vssd1 vccd1 vccd1 _11554_/B
+ sky130_fd_sc_hd__nand4_1
X_20749_ _20650_/A _20648_/A _20650_/B vssd1 vssd1 vccd1 vccd1 _20751_/B sky130_fd_sc_hd__a21boi_2
XFILLER_196_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21684__A3 _21399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14270_ _14270_/A vssd1 vssd1 vccd1 vccd1 _14575_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_156_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11482_ _22789_/Q _22788_/Q vssd1 vssd1 vccd1 vccd1 _12146_/A sky130_fd_sc_hd__nor2_2
XFILLER_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13221_ _13221_/A _13221_/B _13221_/C vssd1 vssd1 vccd1 vccd1 _13475_/B sky130_fd_sc_hd__nand3_2
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18298__C1 _18305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22419_ _22419_/A vssd1 vssd1 vccd1 vccd1 _22709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13152_ _22844_/Q vssd1 vssd1 vccd1 vccd1 _21495_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_input64_A wb_dat_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ _11625_/X _11626_/X _16912_/A _12099_/Y vssd1 vssd1 vccd1 vccd1 _12110_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14323__A1 _18953_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17960_ _17960_/A _18002_/C _18002_/A _17960_/D vssd1 vssd1 vccd1 vccd1 _17967_/C
+ sky130_fd_sc_hd__nand4_2
X_13083_ _21351_/A _21351_/B _21312_/B vssd1 vssd1 vccd1 vccd1 _13316_/A sky130_fd_sc_hd__nand3_2
XANTENNA__14323__B2 _14220_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16911_ _16911_/A vssd1 vssd1 vccd1 vccd1 _16911_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12034_ _12034_/A _12034_/B vssd1 vssd1 vccd1 vccd1 _12034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_622 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17891_ _17891_/A _17891_/B vssd1 vssd1 vccd1 vccd1 _17893_/A sky130_fd_sc_hd__nand2_1
XFILLER_120_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19630_ _19630_/A _19630_/B _19630_/C _19630_/D vssd1 vssd1 vccd1 vccd1 _19724_/A
+ sky130_fd_sc_hd__nand4_4
X_16842_ _16842_/A _16842_/B _16842_/C vssd1 vssd1 vccd1 vccd1 _16843_/B sky130_fd_sc_hd__nand3_1
XFILLER_78_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19561_ _19561_/A _19561_/B _19577_/A _19577_/B vssd1 vssd1 vccd1 vccd1 _19669_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16773_ _16773_/A _16773_/B vssd1 vssd1 vccd1 vccd1 _16776_/B sky130_fd_sc_hd__nand2_1
X_13985_ _13985_/A _13985_/B _14200_/A vssd1 vssd1 vccd1 vccd1 _13986_/B sky130_fd_sc_hd__nand3_2
XFILLER_93_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18512_ _18512_/A _18512_/B _18512_/C vssd1 vssd1 vccd1 vccd1 _18512_/X sky130_fd_sc_hd__or3_1
XFILLER_19_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15724_ _16450_/B vssd1 vssd1 vccd1 vccd1 _20870_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15604__A _22700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12936_ _12988_/A _12721_/X _12934_/X _12935_/Y vssd1 vssd1 vccd1 vccd1 _12937_/A
+ sky130_fd_sc_hd__o22ai_2
X_19492_ _19352_/X _19490_/Y _19491_/Y vssd1 vssd1 vccd1 vccd1 _19492_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21325__B _21595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18443_ _18443_/A _18443_/B vssd1 vssd1 vccd1 vccd1 _18443_/Y sky130_fd_sc_hd__nand2_2
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15323__B _18690_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15655_ _15601_/Y _15602_/X _15644_/Y _15654_/Y vssd1 vssd1 vccd1 vccd1 _15673_/B
+ sky130_fd_sc_hd__o211ai_4
X_12867_ _12867_/A _12867_/B _12867_/C vssd1 vssd1 vccd1 vccd1 _12868_/A sky130_fd_sc_hd__nand3_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16784__C1 _19694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11818_ _11818_/A vssd1 vssd1 vccd1 vccd1 _18778_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14606_ _14600_/Y _14602_/Y _14604_/Y _14605_/X vssd1 vssd1 vccd1 vccd1 _14606_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_57_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15586_ _16770_/A _16771_/A _15586_/C vssd1 vssd1 vccd1 vccd1 _15587_/A sky130_fd_sc_hd__and3_1
X_18374_ _18090_/Y _18091_/Y _18370_/X vssd1 vssd1 vccd1 vccd1 _18387_/C sky130_fd_sc_hd__a21oi_2
XFILLER_57_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _20134_/C vssd1 vssd1 vccd1 vccd1 _20508_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _17324_/B _17324_/C _17341_/B vssd1 vssd1 vccd1 vccd1 _17333_/D sky130_fd_sc_hd__a21o_1
X_14537_ _14524_/Y _14535_/X _14536_/Y vssd1 vssd1 vccd1 vccd1 _14537_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_187_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11749_ _11749_/A vssd1 vssd1 vccd1 vccd1 _17421_/A sky130_fd_sc_hd__buf_2
XANTENNA__19449__C _22917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16435__A _18259_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17256_ _17138_/X _17142_/X _17149_/B _17145_/Y vssd1 vssd1 vccd1 vccd1 _17260_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_14468_ _14468_/A _14468_/B vssd1 vssd1 vccd1 vccd1 _14468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15696__D _15696_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16207_ _15952_/A _15952_/B _15952_/C _16034_/C vssd1 vssd1 vccd1 vccd1 _16210_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12168__A3 _12167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13419_ _13419_/A _13419_/B vssd1 vssd1 vccd1 vccd1 _13494_/B sky130_fd_sc_hd__xor2_2
X_17187_ _16908_/X _16909_/X _16982_/Y _16983_/X vssd1 vssd1 vccd1 vccd1 _17187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12022__C1 _12006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14399_ _22804_/Q _14397_/X _14398_/X _14370_/A _22708_/Q vssd1 vssd1 vccd1 vccd1
+ _14399_/X sky130_fd_sc_hd__a32o_1
XFILLER_143_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16138_ _16069_/X _16068_/Y _16055_/Y _16064_/Y _16070_/Y vssd1 vssd1 vccd1 vccd1
+ _16169_/A sky130_fd_sc_hd__a311o_1
XANTENNA__19465__B _19614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16069_ _19470_/D _16110_/B _16106_/D vssd1 vssd1 vccd1 vccd1 _16069_/X sky130_fd_sc_hd__and3_2
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12325__B1 _12320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19828_ _19757_/A _19757_/B _19827_/Y vssd1 vssd1 vccd1 vccd1 _19891_/A sky130_fd_sc_hd__o21bai_1
XANTENNA__19481__A _19481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12203__A _19587_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14078__B1 _14079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14617__A2 _14765_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19759_ _19759_/A _19759_/B vssd1 vssd1 vccd1 vccd1 _22900_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__22921__CLK _22922_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17016__B1 _16726_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22770_ _22802_/CLK _22770_/D vssd1 vssd1 vccd1 vccd1 _22770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21721_ _21721_/A _21721_/B vssd1 vssd1 vccd1 vccd1 _21801_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11851__A2 _12003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20571__B1 _20723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21652_ _21651_/X _21805_/D _21515_/Y vssd1 vssd1 vccd1 vccd1 _21652_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_178_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20603_ _20629_/C _20603_/B _20603_/C vssd1 vssd1 vccd1 vccd1 _20603_/X sky130_fd_sc_hd__and3_1
XANTENNA__20793__C _20793_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_700 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21583_ _13073_/A _21583_/B _21583_/C _21583_/D vssd1 vssd1 vccd1 vccd1 _21584_/A
+ sky130_fd_sc_hd__nand4b_1
XANTENNA__14791__C _22765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13688__B _22672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20534_ _20534_/A _20568_/B _20568_/A vssd1 vssd1 vccd1 vccd1 _20535_/C sky130_fd_sc_hd__nand3_1
XFILLER_177_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20465_ _13022_/C _16745_/A _20587_/A _20587_/B _20581_/A vssd1 vssd1 vccd1 vccd1
+ _20465_/X sky130_fd_sc_hd__o221a_1
XFILLER_193_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22204_ _22336_/A _22157_/Y _22212_/C vssd1 vssd1 vccd1 vccd1 _22206_/A sky130_fd_sc_hd__o21ai_1
XFILLER_152_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18295__A2 _17526_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20396_ _20396_/A _20396_/B vssd1 vssd1 vccd1 vccd1 _20427_/A sky130_fd_sc_hd__nand2_1
XFILLER_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22135_ _22135_/A _22135_/B _22170_/B _22135_/D vssd1 vssd1 vccd1 vccd1 _22137_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12316__B1 _12320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11936__B _18093_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22066_ _22131_/A _22196_/B _22132_/B _22135_/A vssd1 vssd1 vccd1 vccd1 _22068_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_82_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19795__A2 _17422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21017_ _21017_/A _21017_/B _21017_/C vssd1 vssd1 vccd1 vccd1 _21018_/B sky130_fd_sc_hd__and3_1
XFILLER_181_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12113__A _16274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15805__A1 _12988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_bq_clk_i clkbuf_3_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_bq_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_114_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15281__A2 _15271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ _14181_/A _14506_/B _14181_/C _14203_/B _14107_/A vssd1 vssd1 vccd1 vccd1
+ _13781_/A sky130_fd_sc_hd__a32o_1
X_22968_ _22968_/CLK _22968_/D vssd1 vssd1 vccd1 vccd1 _22968_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12721_ _12721_/A vssd1 vssd1 vccd1 vccd1 _12721_/X sky130_fd_sc_hd__clkbuf_4
X_21919_ _21836_/Y _21916_/Y _21918_/Y vssd1 vssd1 vccd1 vccd1 _21931_/A sky130_fd_sc_hd__a21oi_2
XFILLER_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22899_ _22951_/CLK _22899_/D vssd1 vssd1 vccd1 vccd1 _22899_/Q sky130_fd_sc_hd__dfxtp_2
X_15440_ _15440_/A vssd1 vssd1 vccd1 vccd1 _17234_/A sky130_fd_sc_hd__buf_2
X_12652_ _12898_/A _12898_/B vssd1 vssd1 vccd1 vccd1 _12666_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ _12003_/C vssd1 vssd1 vccd1 vccd1 _11627_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15371_ _17423_/A _17424_/A vssd1 vssd1 vccd1 vccd1 _20456_/B sky130_fd_sc_hd__nand2_1
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12583_ _12583_/A _12630_/A _12583_/C vssd1 vssd1 vccd1 vccd1 _12630_/B sky130_fd_sc_hd__nand3_2
XANTENNA__16368__A2_N _16627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17110_ _17110_/A _17110_/B vssd1 vssd1 vccd1 vccd1 _17116_/B sky130_fd_sc_hd__nand2_2
X_14322_ _14413_/A vssd1 vssd1 vccd1 vccd1 _14322_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11534_ _12008_/A vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__clkbuf_4
X_18090_ _18116_/A _11430_/B _11846_/B _11666_/X _15690_/X vssd1 vssd1 vccd1 vccd1
+ _18090_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_184_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17041_ _17040_/A _17208_/A _17040_/C vssd1 vssd1 vccd1 vccd1 _17041_/X sky130_fd_sc_hd__a21o_1
XFILLER_144_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11399__A _11942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14253_ _14253_/A _14253_/B _14253_/C _14253_/D vssd1 vssd1 vccd1 vccd1 _14253_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_171_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11465_ _15776_/A vssd1 vssd1 vccd1 vccd1 _15901_/A sky130_fd_sc_hd__buf_4
XFILLER_184_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11358__A1 _15484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1080 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _13517_/A vssd1 vssd1 vccd1 vccd1 _21398_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14184_ _14184_/A _14184_/B _14184_/C vssd1 vssd1 vccd1 vccd1 _14259_/A sky130_fd_sc_hd__nand3_4
XFILLER_136_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11396_ _18259_/A _11395_/X _11384_/A vssd1 vssd1 vccd1 vccd1 _11942_/A sky130_fd_sc_hd__o21bai_4
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16297__A1 _12403_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13135_ _21367_/A _21367_/B _21315_/B vssd1 vssd1 vccd1 vccd1 _13180_/B sky130_fd_sc_hd__and3_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16836__A3 _16452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18992_ _19156_/D _18984_/Y _18986_/Y _18991_/Y _18881_/X vssd1 vssd1 vccd1 vccd1
+ _19187_/C sky130_fd_sc_hd__o2111ai_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14503__A _14503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _17893_/B _17896_/A _17945_/A vssd1 vssd1 vccd1 vccd1 _17946_/A sky130_fd_sc_hd__a21o_1
XFILLER_97_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _22727_/Q _22726_/Q vssd1 vssd1 vccd1 vccd1 _21469_/B sky130_fd_sc_hd__nor2_2
XFILLER_105_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22944__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14222__B _14494_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12017_ _12017_/A _18367_/C _17312_/A vssd1 vssd1 vccd1 vccd1 _12017_/X sky130_fd_sc_hd__and3_1
XANTENNA__17814__A _19769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17874_ _17874_/A vssd1 vssd1 vccd1 vccd1 _21048_/B sky130_fd_sc_hd__buf_2
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11530__A1 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18994__B1 _15981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19613_ _19605_/Y _19610_/Y _19612_/X vssd1 vssd1 vccd1 vccd1 _19613_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18629__B _18629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16825_ _19614_/A _18849_/D _17539_/D _17407_/A vssd1 vssd1 vccd1 vccd1 _16825_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17533__B _20870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11862__A _16106_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15272__A2 _15271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19544_ _19650_/A _19540_/Y _19543_/Y vssd1 vssd1 vccd1 vccd1 _19545_/C sky130_fd_sc_hd__a21o_1
XANTENNA__15334__A _16313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18348__C _18483_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16756_ _16866_/C _16866_/D vssd1 vssd1 vccd1 vccd1 _16847_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13968_ _14565_/A _14566_/A _13968_/C vssd1 vssd1 vccd1 vccd1 _13968_/Y sky130_fd_sc_hd__nand3_2
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15707_ _15707_/A _15707_/B vssd1 vssd1 vccd1 vccd1 _15709_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19475_ _19476_/C _19476_/A _19476_/B vssd1 vssd1 vccd1 vccd1 _19475_/Y sky130_fd_sc_hd__a21oi_2
X_12919_ _13002_/A _13002_/B _12920_/C vssd1 vssd1 vccd1 vccd1 _12963_/A sky130_fd_sc_hd__a21o_1
X_16687_ _16669_/A _16670_/A _16686_/Y _16424_/Y vssd1 vssd1 vccd1 vccd1 _16690_/C
+ sky130_fd_sc_hd__o211ai_1
X_13899_ _13899_/A _13899_/B vssd1 vssd1 vccd1 vccd1 _13996_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16221__A1 _12929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18426_ _18772_/C _18274_/Y _18425_/Y vssd1 vssd1 vccd1 vccd1 _18601_/A sky130_fd_sc_hd__a21o_1
XFILLER_22_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15638_ _15638_/A vssd1 vssd1 vccd1 vccd1 _15638_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15988__B _15988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22167__A _22167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18357_ _18663_/A _19322_/A _18797_/C _19318_/A vssd1 vssd1 vccd1 vccd1 _18367_/A
+ sky130_fd_sc_hd__nand4_4
XANTENNA__12693__A _15394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15569_ _15569_/A vssd1 vssd1 vccd1 vccd1 _16039_/A sky130_fd_sc_hd__buf_4
XANTENNA__19171__B1 _19334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17308_ _17475_/A _17475_/B _17475_/C vssd1 vssd1 vccd1 vccd1 _17334_/B sky130_fd_sc_hd__nand3_1
XFILLER_148_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18288_ _18288_/A _19199_/B _19199_/C vssd1 vssd1 vccd1 vccd1 _18296_/B sky130_fd_sc_hd__and3_2
XFILLER_119_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17239_ _17129_/Y _17237_/Y _17238_/X vssd1 vssd1 vccd1 vccd1 _17239_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20250_ _20502_/A _20502_/B _20250_/C vssd1 vssd1 vccd1 vccd1 _20250_/X sky130_fd_sc_hd__and3_1
XANTENNA__19474__A1 _19838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20084__A2 _16708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20181_ _20181_/A _20181_/B vssd1 vssd1 vccd1 vccd1 _20184_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19226__A1 _18131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16460__A1 _11935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22822_ _22929_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 _22822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22753_ _22757_/CLK _22753_/D vssd1 vssd1 vccd1 vccd1 _22753_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16748__C1 _16723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21704_ _21704_/A _22676_/Q _21704_/C vssd1 vssd1 vccd1 vccd1 _21706_/A sky130_fd_sc_hd__nand3_1
XFILLER_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13026__A1 _16157_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22684_ _22943_/CLK _22684_/D vssd1 vssd1 vccd1 vccd1 _22684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_514 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21635_ _21716_/A _21716_/B _21635_/C _21635_/D vssd1 vssd1 vccd1 vccd1 _21654_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19162__B1 _19792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22817__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20309__B _20553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20847__A1 _20793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20847__B2 _20793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21566_ _21566_/A _21566_/B vssd1 vssd1 vccd1 vccd1 _21707_/B sky130_fd_sc_hd__nand2_1
XFILLER_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20517_ _20514_/X _15934_/A _20244_/X _20328_/D vssd1 vssd1 vccd1 vccd1 _20519_/C
+ sky130_fd_sc_hd__o31a_2
XFILLER_5_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21497_ _21383_/A _21220_/X _21493_/Y _21610_/A _21716_/A vssd1 vssd1 vccd1 vccd1
+ _21501_/A sky130_fd_sc_hd__o221ai_4
XFILLER_181_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20448_ _20335_/B _20335_/C _20447_/Y vssd1 vssd1 vccd1 vccd1 _20449_/C sky130_fd_sc_hd__a21oi_2
XFILLER_107_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20075__A2 _12525_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15419__A _16058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13865__C _14808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20379_ _20204_/X _20205_/Y _20229_/Y _20232_/Y vssd1 vssd1 vccd1 vccd1 _20379_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22118_ _22037_/C _22105_/X _22044_/X _22171_/B _22173_/D vssd1 vssd1 vccd1 vccd1
+ _22119_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17634__A _17634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22049_ _22045_/Y _22048_/Y _22044_/X _22039_/Y vssd1 vssd1 vccd1 vccd1 _22049_/X
+ sky130_fd_sc_hd__o211a_1
X_14940_ _14862_/A _14996_/D _14877_/C _14939_/Y vssd1 vssd1 vccd1 vccd1 _15001_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_85_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21575__A2 _21551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input27_A wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14871_ _14871_/A _14871_/B vssd1 vssd1 vccd1 vccd1 _14933_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12778__A _12968_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20783__B1 _20913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16610_ _16996_/A vssd1 vssd1 vccd1 vccd1 _17431_/C sky130_fd_sc_hd__buf_2
XFILLER_91_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13822_ _22866_/Q vssd1 vssd1 vccd1 vccd1 _13831_/A sky130_fd_sc_hd__inv_2
X_17590_ _17586_/Y _17590_/B _17590_/C vssd1 vssd1 vccd1 vccd1 _17625_/A sky130_fd_sc_hd__nand3b_2
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21327__A2 _13633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ _16493_/A _16493_/B _16508_/X _16510_/Y _16524_/Y vssd1 vssd1 vccd1 vccd1
+ _16541_/X sky130_fd_sc_hd__o221a_1
XFILLER_141_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13753_ _22865_/Q vssd1 vssd1 vccd1 vccd1 _13975_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16739__C1 _16723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18597__A1_N _12250_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ _12704_/A vssd1 vssd1 vccd1 vccd1 _12727_/A sky130_fd_sc_hd__clkbuf_4
X_19260_ _19192_/Y _19238_/Y _19248_/Y _19249_/Y vssd1 vssd1 vccd1 vccd1 _19260_/X
+ sky130_fd_sc_hd__o211a_1
X_16472_ _19351_/B _18797_/B _20129_/B _16772_/A _17631_/A vssd1 vssd1 vccd1 vccd1
+ _16472_/Y sky130_fd_sc_hd__a32oi_4
X_13684_ _13558_/C _13557_/X _13679_/X _13612_/Y _13683_/Y vssd1 vssd1 vccd1 vccd1
+ _21285_/C sky130_fd_sc_hd__o221ai_4
X_18211_ _18214_/B _18214_/C _18214_/A _12230_/C _18228_/A vssd1 vssd1 vccd1 vccd1
+ _18232_/B sky130_fd_sc_hd__a32oi_4
XFILLER_70_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15423_ _18716_/A _15774_/B _20129_/A _15774_/C vssd1 vssd1 vccd1 vccd1 _15423_/Y
+ sky130_fd_sc_hd__nand4_1
X_12635_ _20130_/C vssd1 vssd1 vccd1 vccd1 _20675_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_176_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19191_ _19240_/A _19240_/B _19343_/B _19343_/C vssd1 vssd1 vccd1 vccd1 _19237_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_19_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19153__B1 _18514_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11579__A1 _15357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18142_ _18137_/Y _18139_/X _18141_/Y vssd1 vssd1 vccd1 vccd1 _18150_/A sky130_fd_sc_hd__o21ai_1
X_15354_ _15370_/A _16322_/A vssd1 vssd1 vccd1 vccd1 _15355_/B sky130_fd_sc_hd__nand2_4
X_12566_ _15299_/C vssd1 vssd1 vccd1 vccd1 _12681_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11517_ _11796_/A vssd1 vssd1 vccd1 vccd1 _18348_/A sky130_fd_sc_hd__clkbuf_1
X_14305_ _14305_/A _14305_/B _14305_/C _14305_/D vssd1 vssd1 vccd1 vccd1 _14310_/A
+ sky130_fd_sc_hd__nor4_1
X_18073_ _18082_/C _18069_/C _18066_/X _18072_/Y vssd1 vssd1 vccd1 vccd1 _18082_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_15285_ _22881_/Q _22882_/Q _15287_/D _22876_/D vssd1 vssd1 vccd1 vccd1 _15286_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_144_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _12497_/A vssd1 vssd1 vccd1 vccd1 _12704_/A sky130_fd_sc_hd__buf_2
XFILLER_8_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17024_ _17009_/X _17011_/Y _17023_/X _16742_/Y vssd1 vssd1 vccd1 vccd1 _17024_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14236_ _14236_/A _14236_/B _14236_/C vssd1 vssd1 vccd1 vccd1 _14246_/A sky130_fd_sc_hd__nand3_1
XFILLER_176_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11448_ _11448_/A vssd1 vssd1 vccd1 vccd1 _11778_/A sky130_fd_sc_hd__buf_2
XFILLER_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20066__A2 _20064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14167_ _14167_/A _14167_/B _14167_/C vssd1 vssd1 vccd1 vccd1 _14167_/X sky130_fd_sc_hd__and3_1
XANTENNA__20507__A2_N _20511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11379_ _11394_/A _11378_/X _11299_/X vssd1 vssd1 vccd1 vccd1 _11380_/B sky130_fd_sc_hd__o21ai_4
XFILLER_153_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11751__A1 _17421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13118_ _13099_/B _13098_/A _13095_/A _13126_/A vssd1 vssd1 vccd1 vccd1 _13168_/C
+ sky130_fd_sc_hd__a31oi_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18975_ _18945_/A _18945_/B _18945_/C vssd1 vssd1 vccd1 vccd1 _18975_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_113_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14098_ _14098_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14099_/A sky130_fd_sc_hd__xnor2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _19839_/C vssd1 vssd1 vccd1 vccd1 _19941_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13049_ _22843_/Q vssd1 vssd1 vccd1 vccd1 _13176_/A sky130_fd_sc_hd__inv_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17857_ _17857_/A _17857_/B vssd1 vssd1 vccd1 vccd1 _17861_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16808_ _16275_/A _15933_/A _16911_/A vssd1 vssd1 vccd1 vccd1 _16810_/C sky130_fd_sc_hd__o21ai_4
XFILLER_94_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18982__A3 _18890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14453__B1 _14448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17788_ _17799_/A _17799_/B vssd1 vssd1 vccd1 vccd1 _17788_/X sky130_fd_sc_hd__and2_1
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15650__C1 _16361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19527_ _19536_/A _19536_/B _19524_/X _19526_/Y vssd1 vssd1 vccd1 vccd1 _19528_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16739_ _16736_/Y _16738_/X _16732_/Y _16723_/X vssd1 vssd1 vccd1 vccd1 _16739_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11806__A2 _11809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18195__A1 _11634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19458_ _19458_/A _19458_/B vssd1 vssd1 vccd1 vccd1 _19458_/Y sky130_fd_sc_hd__nand2_1
X_18409_ _18183_/Y _18395_/X _18408_/X _18393_/Y vssd1 vssd1 vccd1 vccd1 _18409_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_22_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ _19457_/A _19389_/B _19389_/C vssd1 vssd1 vccd1 vccd1 _19389_/X sky130_fd_sc_hd__and3_1
XANTENNA__20129__B _20129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21420_ _21421_/A _21560_/B vssd1 vssd1 vccd1 vccd1 _21420_/X sky130_fd_sc_hd__and2_1
XFILLER_148_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15705__B1 _15700_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21351_ _21351_/A _21351_/B _21351_/C vssd1 vssd1 vccd1 vccd1 _21496_/A sky130_fd_sc_hd__nand3_1
XFILLER_175_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20302_ _12754_/X _12894_/Y _13045_/Y _20314_/C vssd1 vssd1 vccd1 vccd1 _20442_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21282_ _21282_/A _21282_/B _21419_/B vssd1 vssd1 vccd1 vccd1 _21422_/B sky130_fd_sc_hd__nand3_4
XFILLER_190_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22451__A0 _13202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20233_ _20204_/X _20205_/Y _20229_/Y _20232_/Y vssd1 vssd1 vccd1 vccd1 _20234_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_115_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20164_ _12868_/X _20163_/X _20169_/A vssd1 vssd1 vccd1 vccd1 _20165_/C sky130_fd_sc_hd__a21boi_4
XANTENNA__11917__D _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16681__A1 _17502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13982__A _22868_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20095_ _20101_/A _20101_/B _20357_/B vssd1 vssd1 vccd1 vccd1 _20096_/B sky130_fd_sc_hd__nand3_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15405__C _15799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22805_ _22805_/CLK _22805_/D vssd1 vssd1 vccd1 vccd1 _22805_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20997_ _21066_/A _21067_/A _21006_/B _21006_/A vssd1 vssd1 vccd1 vccd1 _20999_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18716__C _19358_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22736_ _22768_/CLK _22736_/D vssd1 vssd1 vccd1 vccd1 _22736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1085 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17933__A1 _19941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22667_ _22959_/CLK _22667_/D vssd1 vssd1 vccd1 vccd1 _22667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14318__A input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12420_ _15335_/A vssd1 vssd1 vccd1 vccd1 _12420_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21618_ _21846_/A _21763_/A _21763_/B vssd1 vssd1 vccd1 vccd1 _21618_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_187_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19686__B2 _18718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22598_ _22598_/A vssd1 vssd1 vccd1 vccd1 _22788_/D sky130_fd_sc_hd__clkbuf_1
X_12351_ _12428_/B vssd1 vssd1 vccd1 vccd1 _12734_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21549_ _21553_/B _21553_/C vssd1 vssd1 vccd1 vccd1 _21551_/A sky130_fd_sc_hd__nand2_2
XFILLER_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ _11302_/A vssd1 vssd1 vccd1 vccd1 _11377_/A sky130_fd_sc_hd__buf_2
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15070_ _15070_/A vssd1 vssd1 vccd1 vccd1 _15186_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13876__B _14722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12282_ _12340_/A vssd1 vssd1 vccd1 vccd1 _16319_/A sky130_fd_sc_hd__buf_2
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ _14021_/A _14021_/B _14021_/C _14021_/D vssd1 vssd1 vccd1 vccd1 _14022_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_135_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17364__A _22897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15475__A2 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14278__A3 _14834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18760_ _18572_/X _18571_/X _18575_/B vssd1 vssd1 vccd1 vccd1 _18761_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__14203__D _14786_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15972_ _16241_/A _11988_/X _12772_/X _12774_/X _15901_/A vssd1 vssd1 vccd1 vccd1
+ _15972_/X sky130_fd_sc_hd__o221a_4
XFILLER_103_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20502__B _20502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17711_ _17605_/B _17605_/A _17781_/C _17781_/B vssd1 vssd1 vccd1 vccd1 _17790_/C
+ sky130_fd_sc_hd__o211ai_2
X_14923_ _14923_/A _14923_/B vssd1 vssd1 vccd1 vccd1 _14982_/B sky130_fd_sc_hd__nand2_1
X_18691_ _18691_/A _18691_/B _18691_/C vssd1 vssd1 vccd1 vccd1 _18691_/Y sky130_fd_sc_hd__nand3_1
XFILLER_48_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20221__C _20456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17642_ _19687_/C vssd1 vssd1 vccd1 vccd1 _19768_/D sky130_fd_sc_hd__buf_2
XFILLER_152_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14854_ _14854_/A vssd1 vssd1 vccd1 vccd1 _14854_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16975__A2 _16944_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15632__C1 _15633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13805_ _22866_/Q vssd1 vssd1 vccd1 vccd1 _14118_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_189_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17811__B _20936_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17573_ _17574_/C _17574_/B _17574_/A vssd1 vssd1 vccd1 vccd1 _17573_/Y sky130_fd_sc_hd__a21oi_1
X_11997_ _18140_/A vssd1 vssd1 vccd1 vccd1 _12135_/B sky130_fd_sc_hd__clkbuf_2
X_14785_ _14785_/A _14785_/B _14786_/C vssd1 vssd1 vccd1 vccd1 _14793_/B sky130_fd_sc_hd__nand3_1
XANTENNA__16708__A _16708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19312_ _19000_/Y _19156_/Y _19311_/Y vssd1 vssd1 vccd1 vccd1 _19340_/A sky130_fd_sc_hd__a21oi_4
XFILLER_72_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16524_ _16524_/A _16524_/B vssd1 vssd1 vccd1 vccd1 _16524_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__15612__A _16611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13736_ _13869_/B _13736_/B _13736_/C vssd1 vssd1 vccd1 vccd1 _13750_/A sky130_fd_sc_hd__nand3_1
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16727__A2 _11295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21720__A2 _21522_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19243_ _19239_/X _19242_/Y _19396_/C vssd1 vssd1 vccd1 vccd1 _19248_/A sky130_fd_sc_hd__o21ai_1
XFILLER_189_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16455_ _15530_/A _15531_/A _15450_/A vssd1 vssd1 vccd1 vccd1 _16455_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15331__B _15901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_7_0_bq_clk_i_A clkbuf_3_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ _13666_/X _13641_/Y _13640_/Y vssd1 vssd1 vccd1 vccd1 _13667_/X sky130_fd_sc_hd__o21ba_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15406_ _15406_/A vssd1 vssd1 vccd1 vccd1 _15406_/X sky130_fd_sc_hd__buf_2
X_19174_ _19174_/A _19174_/B vssd1 vssd1 vccd1 vccd1 _19174_/Y sky130_fd_sc_hd__nand2_1
X_12618_ _12618_/A _12618_/B _12618_/C vssd1 vssd1 vccd1 vccd1 _12619_/A sky130_fd_sc_hd__nand3_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _16386_/A _16386_/B _16386_/C vssd1 vssd1 vccd1 vccd1 _16431_/C sky130_fd_sc_hd__nand3_1
X_13598_ _13627_/C _13589_/X _13627_/B vssd1 vssd1 vccd1 vccd1 _13598_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18125_ _18363_/A vssd1 vssd1 vccd1 vccd1 _18125_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17539__A _17645_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15337_ _20611_/A vssd1 vssd1 vccd1 vccd1 _16809_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__13961__A2 _13736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12549_ _12549_/A _15363_/C vssd1 vssd1 vccd1 vccd1 _12550_/B sky130_fd_sc_hd__nand2_1
XFILLER_184_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17152__A2 _16758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_595 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18056_ _22905_/Q _18055_/X _18051_/Y _18077_/A _18053_/Y vssd1 vssd1 vccd1 vccd1
+ _18057_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16360__B1 _16400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ _22816_/D _15265_/X _15268_/S vssd1 vssd1 vccd1 vccd1 _15269_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17007_ _17007_/A vssd1 vssd1 vccd1 vccd1 _17728_/A sky130_fd_sc_hd__buf_4
XANTENNA__19754__A _22920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18637__C1 _18953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14219_ _15004_/D vssd1 vssd1 vccd1 vccd1 _15118_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15199_ _15210_/A _15199_/B vssd1 vssd1 vccd1 vccd1 _15200_/B sky130_fd_sc_hd__xnor2_1
XFILLER_153_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16112__B1 _16106_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18652__A2 _11786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18958_ _18958_/A _18958_/B _19132_/B vssd1 vssd1 vccd1 vccd1 _19138_/C sky130_fd_sc_hd__nand3_1
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14674__B1 _14057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_591 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17909_ _17785_/X _17954_/B _17860_/B _17860_/A _17908_/Y vssd1 vssd1 vccd1 vccd1
+ _17959_/B sky130_fd_sc_hd__o221ai_4
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18889_ _19316_/B vssd1 vssd1 vccd1 vccd1 _18889_/X sky130_fd_sc_hd__buf_2
XANTENNA__21227__C _21638_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20747__B1 _20748_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20920_ _20920_/A _20920_/B _20920_/C vssd1 vssd1 vccd1 vccd1 _20923_/C sky130_fd_sc_hd__nand3_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12211__A _12211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14426__B1 _14351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1044 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17721__B _22900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20851_ _20849_/X _20797_/B _20850_/Y vssd1 vssd1 vccd1 vccd1 _20851_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19365__B1 _19350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20782_ _20782_/A _20782_/B vssd1 vssd1 vccd1 vccd1 _20782_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22521_ _13761_/B input57/X _22525_/S vssd1 vssd1 vccd1 vccd1 _22522_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22452_ _22452_/A vssd1 vssd1 vccd1 vccd1 _22723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21403_ _21403_/A vssd1 vssd1 vccd1 vccd1 _21403_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20278__A2 _15890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22383_ _12273_/B input62/X _22391_/S vssd1 vssd1 vccd1 vccd1 _22384_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21334_ _21351_/A vssd1 vssd1 vccd1 vccd1 _21725_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_191_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18891__A2 _18889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18628__C1 _18830_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21265_ _21243_/A _21243_/B _21243_/C vssd1 vssd1 vccd1 vccd1 _21265_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_190_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20216_ _20341_/A _20341_/B _22818_/Q vssd1 vssd1 vccd1 vccd1 _20217_/A sky130_fd_sc_hd__and3_1
X_21196_ _21185_/A _21187_/A _22841_/Q _21480_/A vssd1 vssd1 vccd1 vccd1 _21301_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__11647__D _11647_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20450__A2 _20449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17851__B1 _22902_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20147_ _20147_/A _20147_/B vssd1 vssd1 vccd1 vccd1 _20150_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19053__C1 _18795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ _20200_/A vssd1 vssd1 vccd1 vccd1 _20293_/B sky130_fd_sc_hd__buf_2
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13217__A _21480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20202__A2 _20115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18946__A3 _18953_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11920_ _12074_/A _12074_/B _11874_/A vssd1 vssd1 vccd1 vccd1 _11922_/A sky130_fd_sc_hd__a21o_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12121__A _18648_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _15978_/C _12003_/A _11846_/B _17313_/D _12050_/B vssd1 vssd1 vccd1 vccd1
+ _11851_/X sky130_fd_sc_hd__a32o_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18159__A1 _15888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _13973_/B _13907_/X _13970_/X _14593_/B _14775_/C vssd1 vssd1 vccd1 vccd1
+ _14573_/A sky130_fd_sc_hd__o311ai_1
X_11782_ _18116_/A _11430_/B _18507_/C _11846_/B vssd1 vssd1 vccd1 vccd1 _11782_/Y
+ sky130_fd_sc_hd__o211ai_2
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16709__A2 _11905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13521_ _13521_/A _13521_/B _13521_/C vssd1 vssd1 vccd1 vccd1 _13521_/Y sky130_fd_sc_hd__nand3_2
X_22719_ _22815_/CLK _22719_/D vssd1 vssd1 vccd1 vccd1 _22719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17382__A2 _17381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16240_ _15486_/A _15486_/B _15486_/C _14438_/A vssd1 vssd1 vccd1 vccd1 _16240_/X
+ sky130_fd_sc_hd__a31o_2
X_13452_ _13452_/A vssd1 vssd1 vccd1 vccd1 _13461_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16590__B1 _15918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12403_ _12403_/A _15631_/B _15631_/C _12403_/D vssd1 vssd1 vccd1 vccd1 _16294_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_90_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16171_ _16169_/X _16170_/X _16168_/A _16168_/B vssd1 vssd1 vccd1 vccd1 _16171_/Y
+ sky130_fd_sc_hd__o22ai_1
X_13383_ _13385_/B _13385_/C _13382_/Y vssd1 vssd1 vccd1 vccd1 _21251_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12600__C1 _16261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_831 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18331__A1 _16241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15122_ _15113_/X _15060_/X _15146_/A _15121_/X vssd1 vssd1 vccd1 vccd1 _15122_/X
+ sky130_fd_sc_hd__o211a_1
X_12334_ _12334_/A vssd1 vssd1 vccd1 vccd1 _12334_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18882__A2 _19313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19930_ _19970_/A _22923_/Q _19970_/C vssd1 vssd1 vccd1 vccd1 _19973_/A sky130_fd_sc_hd__and3_1
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15053_ _14996_/D _14934_/Y _15001_/C _15052_/X vssd1 vssd1 vccd1 vccd1 _15055_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__20216__C _22818_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12265_ _12396_/A vssd1 vssd1 vccd1 vccd1 _12824_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12941__D _13016_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater129_A _22871_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20426__C1 _20405_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14004_ _14001_/Y _14002_/X _14007_/A vssd1 vssd1 vccd1 vccd1 _14006_/B sky130_fd_sc_hd__o21ai_1
XFILLER_123_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19861_ _19788_/B _19837_/B _19788_/A _19796_/X vssd1 vssd1 vccd1 vccd1 _19861_/Y
+ sky130_fd_sc_hd__a31oi_1
X_12196_ _22961_/Q _22962_/Q vssd1 vssd1 vccd1 vccd1 _12208_/B sky130_fd_sc_hd__or2_2
XFILLER_96_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15448__A2 _19351_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18812_ _11502_/X _11503_/X _17646_/A vssd1 vssd1 vccd1 vccd1 _18812_/Y sky130_fd_sc_hd__o21ai_4
Xoutput82 _14324_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22685__CLK _22943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput93 _14326_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[1] sky130_fd_sc_hd__buf_2
X_19792_ _19792_/A vssd1 vssd1 vccd1 vccd1 _19901_/C sky130_fd_sc_hd__buf_2
XANTENNA__17525__C _17525_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18743_ _18743_/A _18743_/B vssd1 vssd1 vccd1 vccd1 _18748_/A sky130_fd_sc_hd__nand2_1
XFILLER_49_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15955_ _16400_/C _17816_/B _15703_/B _15870_/X vssd1 vssd1 vccd1 vccd1 _15955_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12131__A1 _18512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19595__B1 _19176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17822__A _17822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14906_ _14670_/A _14619_/X _14905_/X _14816_/Y vssd1 vssd1 vccd1 vccd1 _14906_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18674_ _18674_/A _18698_/A vssd1 vssd1 vccd1 vccd1 _18676_/B sky130_fd_sc_hd__nand2_1
X_15886_ _15886_/A _15886_/B vssd1 vssd1 vccd1 vccd1 _15886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12682__A2 _17401_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17625_ _17625_/A _17625_/B vssd1 vssd1 vccd1 vccd1 _17855_/A sky130_fd_sc_hd__nand2_2
XFILLER_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14837_ _14836_/A _14836_/B _14836_/C _14836_/D vssd1 vssd1 vccd1 vccd1 _14838_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15081__B1 _15082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17556_ _17404_/X _17402_/Y _17408_/Y vssd1 vssd1 vccd1 vccd1 _17556_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13631__A1 _21399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14768_ _14768_/A _14768_/B vssd1 vssd1 vccd1 vccd1 _14917_/B sky130_fd_sc_hd__xor2_1
XFILLER_147_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16507_ _16762_/A vssd1 vssd1 vccd1 vccd1 _16507_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13719_ _13725_/A vssd1 vssd1 vccd1 vccd1 _13810_/C sky130_fd_sc_hd__clkinv_2
XFILLER_189_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17487_ _17339_/X _17337_/A _17485_/Y _17486_/X vssd1 vssd1 vccd1 vccd1 _17491_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_32_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14699_ _22764_/Q _14699_/B vssd1 vssd1 vccd1 vccd1 _14791_/B sky130_fd_sc_hd__nand2_2
XFILLER_32_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19226_ _18131_/B _17525_/D _18131_/C _19218_/B _19195_/Y vssd1 vssd1 vccd1 vccd1
+ _19227_/A sky130_fd_sc_hd__a32o_1
XFILLER_177_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16438_ _16438_/A vssd1 vssd1 vccd1 vccd1 _17502_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16581__B1 _16580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22175__A _22229_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22103__C1 _22167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19114__A3 _19113_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19157_ _18996_/A _19007_/B _19002_/A _19002_/B vssd1 vssd1 vccd1 vccd1 _19185_/C
+ sky130_fd_sc_hd__o22ai_4
XFILLER_157_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16369_ _16369_/A _16627_/A _16369_/C vssd1 vssd1 vccd1 vccd1 _16377_/C sky130_fd_sc_hd__nand3_2
XANTENNA__18322__A1 _19322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_882 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_691 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18108_ _18108_/A _18108_/B vssd1 vssd1 vccd1 vccd1 _18109_/C sky130_fd_sc_hd__nand2_1
XFILLER_191_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19088_ _19088_/A _19088_/B _19088_/C vssd1 vssd1 vccd1 vccd1 _19089_/A sky130_fd_sc_hd__nand3_2
XFILLER_117_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16884__A1 _16879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18039_ _18039_/A _18065_/B vssd1 vssd1 vccd1 vccd1 _18040_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19484__A _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20680__A2 _17424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12206__A _15838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21050_ _21090_/A _21050_/B _21050_/C _21050_/D vssd1 vssd1 vccd1 vccd1 _21090_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18625__A2 _17391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20001_ _20001_/A vssd1 vssd1 vccd1 vccd1 _20001_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1054 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14111__A2 _14963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12122__A1 _15694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19586__B1 _18156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17732__A _17732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21952_ _21952_/A _21952_/B _21952_/C vssd1 vssd1 vccd1 vccd1 _21952_/X sky130_fd_sc_hd__and3_1
XFILLER_27_414 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20196__A1 _20195_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19050__A2 _16799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13870__A1 _13799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12673__A2 _12671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21254__A _21990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20903_ _20902_/A _20833_/Y _20776_/X vssd1 vssd1 vccd1 vccd1 _20903_/Y sky130_fd_sc_hd__a21oi_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21883_ _21760_/B _21846_/B _21886_/B vssd1 vssd1 vccd1 vccd1 _21892_/B sky130_fd_sc_hd__a21o_1
XFILLER_55_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12876__A _15746_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20834_ _20834_/A vssd1 vssd1 vccd1 vccd1 _20834_/X sky130_fd_sc_hd__buf_2
XFILLER_126_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16067__B _16067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20765_ _20762_/Y _20907_/A _20827_/D vssd1 vssd1 vccd1 vccd1 _20776_/A sky130_fd_sc_hd__a21o_1
XFILLER_126_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1036 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22504_ _22747_/Q input54/X _22508_/S vssd1 vssd1 vccd1 vccd1 _22505_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15375__B2 _15374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20696_ _20584_/A _20584_/B _13016_/C _16996_/A _20792_/C vssd1 vssd1 vccd1 vccd1
+ _20696_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_167_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22435_ _22717_/Q input56/X _22435_/S vssd1 vssd1 vccd1 vccd1 _22436_/A sky130_fd_sc_hd__mux2_1
XANTENNA__20105__D1 _16304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13925__A2 _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22366_ _22368_/A _22368_/B vssd1 vssd1 vccd1 vccd1 _22946_/D sky130_fd_sc_hd__nor2_1
XFILLER_163_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21317_ _21192_/A _21195_/Y _21203_/X _21201_/Y vssd1 vssd1 vccd1 vccd1 _21320_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_163_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_694 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12116__A _12116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22297_ _22297_/A _22297_/B _22295_/Y vssd1 vssd1 vccd1 vccd1 _22325_/B sky130_fd_sc_hd__or3b_1
XANTENNA__12346__D1 _20086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12050_ _19490_/B _12050_/B _19490_/A vssd1 vssd1 vccd1 vccd1 _12052_/A sky130_fd_sc_hd__and3_4
XFILLER_117_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21248_ _21248_/A _21248_/B _21248_/C vssd1 vssd1 vccd1 vccd1 _21261_/B sky130_fd_sc_hd__nand3_1
XFILLER_78_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21620__A1 _21383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15427__A _15797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21179_ _21179_/A _21179_/B _21179_/C vssd1 vssd1 vccd1 vccd1 _21181_/A sky130_fd_sc_hd__nand3_1
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20974__A3 _21017_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11674__B _11932_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17642__A _19687_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15740_ _15740_/A _15740_/B _15740_/C vssd1 vssd1 vccd1 vccd1 _15864_/A sky130_fd_sc_hd__nand3_4
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19041__A2 _17400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ _16772_/A vssd1 vssd1 vccd1 vccd1 _16100_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20187__A1 _12754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12664__A2 _20723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _11909_/C _11903_/B _11903_/C vssd1 vssd1 vccd1 vccd1 _12079_/C sky130_fd_sc_hd__nand3_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _15677_/A _15678_/C _15678_/D vssd1 vssd1 vccd1 vccd1 _15676_/C sky130_fd_sc_hd__nand3_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12883_ _12868_/X _20169_/A _12777_/X _12781_/X vssd1 vssd1 vccd1 vccd1 _12889_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17410_ _17410_/A vssd1 vssd1 vccd1 vccd1 _17410_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14635_/A vssd1 vssd1 vccd1 vccd1 _14622_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18390_ _18132_/Y _18136_/X _18172_/A vssd1 vssd1 vccd1 vccd1 _18390_/X sky130_fd_sc_hd__o21a_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _11837_/B _12084_/A _11831_/C vssd1 vssd1 vccd1 vccd1 _11834_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17341_/A _17341_/B _17341_/C _17341_/D vssd1 vssd1 vccd1 vccd1 _17341_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_42_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14553_ _14553_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14554_/A sky130_fd_sc_hd__nor2_1
X_11765_ _11995_/A vssd1 vssd1 vccd1 vccd1 _18319_/A sky130_fd_sc_hd__buf_2
XFILLER_92_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _13504_/A _13504_/B _13504_/C vssd1 vssd1 vccd1 vccd1 _13506_/A sky130_fd_sc_hd__or3_1
XFILLER_186_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17272_ _17272_/A _17272_/B _17272_/C vssd1 vssd1 vccd1 vccd1 _17273_/A sky130_fd_sc_hd__nand3_1
X_14484_ _13737_/X _13746_/X _13904_/Y vssd1 vssd1 vccd1 vccd1 _14484_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11696_ _11696_/A _11696_/B _11696_/C vssd1 vssd1 vccd1 vccd1 _12059_/B sky130_fd_sc_hd__nand3_2
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19011_ _19011_/A vssd1 vssd1 vccd1 vccd1 _19687_/D sky130_fd_sc_hd__clkbuf_2
X_16223_ _16940_/A _15450_/X _16247_/A vssd1 vssd1 vccd1 vccd1 _16532_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13435_ _21495_/B vssd1 vssd1 vccd1 vccd1 _21498_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_155_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18304__A1 _18305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11388__C1 _11727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16154_ _16151_/X _16130_/B _20284_/A _16153_/X vssd1 vssd1 vccd1 vccd1 _16154_/X
+ sky130_fd_sc_hd__a31o_1
X_13366_ _13521_/A _21448_/B _13521_/C vssd1 vssd1 vccd1 vccd1 _13366_/Y sky130_fd_sc_hd__nand3_2
XFILLER_10_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20111__A1 _16778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13129__B1 _13055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14326__C1 _14325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15105_ _15085_/A _15085_/B _15081_/X _14948_/C vssd1 vssd1 vccd1 vccd1 _15134_/A
+ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__17817__A _17817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20662__A2 _20551_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ _22818_/Q vssd1 vssd1 vccd1 vccd1 _12428_/B sky130_fd_sc_hd__inv_2
XFILLER_170_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16085_ _16093_/A _16093_/B _16134_/B vssd1 vssd1 vccd1 vccd1 _16085_/Y sky130_fd_sc_hd__nand3_1
X_13297_ _13297_/A _21329_/A vssd1 vssd1 vccd1 vccd1 _21495_/A sky130_fd_sc_hd__nand2_2
XFILLER_138_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19913_ _19913_/A _19913_/B _19913_/C vssd1 vssd1 vccd1 vccd1 _19914_/B sky130_fd_sc_hd__nor3_1
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ _18249_/A _12250_/D vssd1 vssd1 vccd1 vccd1 _12249_/B sky130_fd_sc_hd__nand2_1
X_15036_ _15036_/A vssd1 vssd1 vccd1 vccd1 _15098_/A sky130_fd_sc_hd__inv_2
XFILLER_174_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19454__D _19602_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11865__A _16712_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19844_ _19901_/C _19844_/B _19900_/A _19844_/D vssd1 vssd1 vccd1 vccd1 _19846_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15337__A _20611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20414__A2 _20429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ _12139_/A _12175_/A _12173_/Y _12174_/X vssd1 vssd1 vccd1 vccd1 _12181_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_96_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19775_ _19848_/A _19774_/C _17873_/A _19839_/D vssd1 vssd1 vccd1 vccd1 _19783_/B
+ sky130_fd_sc_hd__o2bb2ai_2
X_16987_ _16845_/A _16986_/Y _16908_/X vssd1 vssd1 vccd1 vccd1 _16989_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12104__A1 _11381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18726_ _18726_/A _18726_/B vssd1 vssd1 vccd1 vccd1 _18726_/Y sky130_fd_sc_hd__nand2_1
X_15938_ _15938_/A vssd1 vssd1 vccd1 vccd1 _15939_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18657_ _18657_/A vssd1 vssd1 vccd1 vccd1 _18865_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11863__B1 _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15869_ _17739_/A vssd1 vssd1 vccd1 vccd1 _17816_/A sky130_fd_sc_hd__buf_4
XANTENNA__12696__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17608_ _17910_/D _17726_/D _17726_/C _17607_/X _17502_/X vssd1 vssd1 vccd1 vccd1
+ _17608_/X sky130_fd_sc_hd__a311o_1
XFILLER_97_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18588_ _19443_/A _18960_/B _18960_/C vssd1 vssd1 vccd1 vccd1 _18595_/A sky130_fd_sc_hd__o21bai_1
XFILLER_178_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _17645_/D _18629_/B _19687_/C _17539_/D vssd1 vssd1 vccd1 vccd1 _17539_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13304__B _13304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20550_ _20442_/A _20442_/B _20549_/Y vssd1 vssd1 vccd1 vccd1 _20550_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_193_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20350__A1 _12734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19209_ _19201_/B _19201_/C _19201_/A vssd1 vssd1 vccd1 vccd1 _19209_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_22_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18533__D _19199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21240__C _21247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20481_ _20579_/A _20579_/B _20481_/C vssd1 vssd1 vccd1 vccd1 _20481_/Y sky130_fd_sc_hd__nand3_1
Xclkbuf_4_8_0_bq_clk_i clkbuf_4_9_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _22968_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22220_ _22220_/A vssd1 vssd1 vccd1 vccd1 _22304_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__22850__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20638__C1 _20178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18700__D1 _15991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12591__A1 _15631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22151_ _22094_/A _22096_/X _22290_/C _22290_/D vssd1 vssd1 vccd1 vccd1 _22151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21102_ _21122_/A _21122_/B _22942_/Q vssd1 vssd1 vccd1 vccd1 _21102_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22082_ _22084_/A _22026_/Y _22160_/A vssd1 vssd1 vccd1 vccd1 _22090_/A sky130_fd_sc_hd__o21bai_1
XFILLER_161_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16609__A1 _15918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16609__B2 _16351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21033_ _21008_/A _21008_/B _21031_/X _21062_/A vssd1 vssd1 vccd1 vccd1 _21067_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_99_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input1_A wb_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16490__C1 _17251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17462__A _17462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13990__A _14013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21935_ _21886_/A _21886_/B _21891_/A _21891_/B vssd1 vssd1 vccd1 vccd1 _21935_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_43_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16078__A _16129_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21866_ _21876_/A _21877_/A _21866_/C vssd1 vssd1 vccd1 vccd1 _21871_/A sky130_fd_sc_hd__nand3_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11606__B1 _15377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _20818_/A _20818_/B _20812_/Y _20816_/Y vssd1 vssd1 vccd1 vccd1 _20822_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_168_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21797_ _21782_/Y _21792_/X _21794_/Y _21796_/X vssd1 vssd1 vccd1 vccd1 _21797_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_179_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18534__B2 _17422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_444 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15710__A _16712_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ _11401_/Y _11895_/A _11895_/B vssd1 vssd1 vccd1 vccd1 _11554_/A sky130_fd_sc_hd__o21ai_1
X_20748_ _20748_/A _20748_/B _20748_/C vssd1 vssd1 vccd1 vccd1 _20751_/C sky130_fd_sc_hd__and3_1
XFILLER_168_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11481_ _22790_/Q vssd1 vssd1 vccd1 vccd1 _18115_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_20679_ _20678_/Y _20676_/Y _20685_/A _15919_/A vssd1 vssd1 vccd1 vccd1 _20682_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_7_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13220_ _13120_/A _13120_/B _21757_/A _13105_/Y _21638_/C vssd1 vssd1 vccd1 vccd1
+ _13221_/C sky130_fd_sc_hd__o2111ai_1
XANTENNA__18298__B1 _18305_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22418_ _22709_/Q input48/X _22424_/S vssd1 vssd1 vccd1 vccd1 _22419_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19836__B _20012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16899__A_N _22894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13151_ _21362_/A _13513_/B _21609_/B _21494_/B vssd1 vssd1 vccd1 vccd1 _13164_/A
+ sky130_fd_sc_hd__nand4_1
X_22349_ _22335_/B _22335_/A _22333_/B _22329_/Y vssd1 vssd1 vccd1 vccd1 _22352_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ _12102_/A _12102_/B _12102_/C vssd1 vssd1 vccd1 vccd1 _18208_/A sky130_fd_sc_hd__nand3_4
XFILLER_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13082_ _22841_/Q vssd1 vssd1 vccd1 vccd1 _21312_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input57_A wb_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16910_ _16792_/B _16787_/Y _16781_/Y _16782_/X vssd1 vssd1 vccd1 vccd1 _16919_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__11685__A _18203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12033_ _11693_/X _11736_/Y _11932_/A _11932_/B vssd1 vssd1 vccd1 vccd1 _12034_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_151_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17890_ _17890_/A _17890_/B vssd1 vssd1 vccd1 vccd1 _17891_/B sky130_fd_sc_hd__and2_1
XFILLER_132_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16841_ _16842_/A _16842_/B _16842_/C vssd1 vssd1 vccd1 vccd1 _16843_/A sky130_fd_sc_hd__a21o_1
XFILLER_120_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19560_ _19556_/Y _19557_/X _19558_/X _19559_/Y vssd1 vssd1 vccd1 vccd1 _19577_/B
+ sky130_fd_sc_hd__o22ai_1
X_16772_ _16772_/A _17405_/A _17406_/A vssd1 vssd1 vccd1 vccd1 _16773_/B sky130_fd_sc_hd__and3_1
XFILLER_59_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13984_ _13984_/A _14564_/C _13984_/C _14684_/B vssd1 vssd1 vccd1 vccd1 _13984_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18511_ _19614_/B _18999_/A _18507_/C _15774_/B _19351_/A vssd1 vssd1 vccd1 vccd1
+ _18511_/Y sky130_fd_sc_hd__a32oi_4
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15723_ _15723_/A vssd1 vssd1 vccd1 vccd1 _15723_/X sky130_fd_sc_hd__clkbuf_4
X_19491_ _19687_/D _17632_/A _19352_/A _19490_/Y vssd1 vssd1 vccd1 vccd1 _19491_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _15804_/C _20593_/C _16937_/B _12711_/X vssd1 vssd1 vccd1 vccd1 _12935_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18442_ _18571_/D _18442_/B _18442_/C vssd1 vssd1 vccd1 vccd1 _18443_/B sky130_fd_sc_hd__nand3_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _15648_/X _15650_/X _15652_/X _15653_/Y vssd1 vssd1 vccd1 vccd1 _15654_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15323__C _17532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12866_ _12510_/B _12564_/B _12865_/Y vssd1 vssd1 vccd1 vccd1 _12867_/C sky130_fd_sc_hd__a21oi_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14605_ _14605_/A _14953_/A _15026_/C _14605_/D vssd1 vssd1 vccd1 vccd1 _14605_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_159_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18373_ _18387_/A _18387_/B _18370_/X _18372_/X vssd1 vssd1 vccd1 vccd1 _18396_/A
+ sky130_fd_sc_hd__o2bb2ai_2
X_11817_ _11932_/A _11932_/B _11685_/X vssd1 vssd1 vccd1 vccd1 _11817_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _12046_/X _15495_/X _14439_/D vssd1 vssd1 vccd1 vccd1 _16771_/A sky130_fd_sc_hd__o21ai_4
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12540_/X _12783_/X _12792_/Y _12796_/Y vssd1 vssd1 vccd1 vccd1 _12863_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16716__A _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17341_/B _17324_/B _17324_/C vssd1 vssd1 vccd1 vccd1 _17333_/C sky130_fd_sc_hd__nand3_1
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22873__CLK _22915_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13745__A_N _13736_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _14541_/B _14541_/C vssd1 vssd1 vccd1 vccd1 _14536_/Y sky130_fd_sc_hd__nand2_1
X_11748_ _11762_/A vssd1 vssd1 vccd1 vccd1 _11932_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_926 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16435__B _16435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17255_ _17255_/A _17255_/B _17255_/C vssd1 vssd1 vccd1 vccd1 _17298_/B sky130_fd_sc_hd__nand3_2
XFILLER_128_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14467_ _14854_/A vssd1 vssd1 vccd1 vccd1 _14467_/X sky130_fd_sc_hd__clkbuf_2
X_11679_ _19316_/A vssd1 vssd1 vccd1 vccd1 _15580_/A sky130_fd_sc_hd__buf_4
XFILLER_174_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16206_ _16206_/A vssd1 vssd1 vccd1 vccd1 _16206_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12022__B1 _12006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13418_ _13494_/A _13495_/C vssd1 vssd1 vccd1 vccd1 _13491_/A sky130_fd_sc_hd__nand2_1
X_17186_ _17200_/A _17200_/B _17200_/C vssd1 vssd1 vccd1 vccd1 _17186_/X sky130_fd_sc_hd__and3_1
XFILLER_128_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14398_ _22442_/B vssd1 vssd1 vccd1 vccd1 _14398_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11376__A2 _11395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _16137_/A _16137_/B _16137_/C vssd1 vssd1 vccd1 vccd1 _16137_/Y sky130_fd_sc_hd__nand3_1
XFILLER_6_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13349_ _21383_/A _13343_/X _13346_/X _21216_/A _13329_/X vssd1 vssd1 vccd1 vccd1
+ _13349_/X sky130_fd_sc_hd__o221a_1
XFILLER_52_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19465__C _19614_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17500__A2 _18044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16068_ _16005_/A _16067_/Y _16098_/A _16155_/A vssd1 vssd1 vccd1 vccd1 _16068_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_97_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15019_ _15018_/A _15018_/B _15018_/C vssd1 vssd1 vccd1 vccd1 _15019_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19827_ _19827_/A _19827_/B vssd1 vssd1 vccd1 vccd1 _19827_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14078__A1 _14722_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14617__A3 _14765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19005__A2 _18893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19758_ _22919_/Q _19674_/A _19674_/B _19757_/Y vssd1 vssd1 vccd1 vccd1 _19759_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17016__A1 _16732_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18709_ _18709_/A _18709_/B _18709_/C vssd1 vssd1 vccd1 vccd1 _18722_/D sky130_fd_sc_hd__nand3_2
X_19689_ _19689_/A _19689_/B _19689_/C _19689_/D vssd1 vssd1 vccd1 vccd1 _19705_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_25_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_564 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21720_ _21219_/C _21522_/D _21654_/C _21654_/A _21717_/Y vssd1 vssd1 vccd1 vccd1
+ _21721_/B sky130_fd_sc_hd__a221oi_2
XFILLER_92_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20571__A1 _15325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21651_ _21463_/A _21651_/B vssd1 vssd1 vccd1 vccd1 _21651_/X sky130_fd_sc_hd__and2b_1
XFILLER_80_876 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18516__A1 _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_28 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15530__A _15530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18516__B2 _18514_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20602_ _20629_/C _20702_/B _20603_/B vssd1 vssd1 vccd1 vccd1 _20602_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_71_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20793__D _20793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21582_ _21582_/A _21582_/B _21582_/C vssd1 vssd1 vccd1 vccd1 _21936_/A sky130_fd_sc_hd__nand3_2
XFILLER_177_252 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_712 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20533_ _20568_/A _20534_/A _20568_/B vssd1 vssd1 vccd1 vccd1 _20535_/B sky130_fd_sc_hd__a21o_1
XFILLER_137_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_756 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20464_ _20464_/A _20464_/B vssd1 vssd1 vccd1 vccd1 _20581_/A sky130_fd_sc_hd__nand2_1
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22203_ _22258_/B vssd1 vssd1 vccd1 vccd1 _22212_/C sky130_fd_sc_hd__inv_2
XFILLER_165_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17457__A _17457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16361__A _16361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20395_ _20395_/A _20395_/B vssd1 vssd1 vccd1 vccd1 _20396_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22134_ _22134_/A _22134_/B vssd1 vssd1 vccd1 vccd1 _22137_/C sky130_fd_sc_hd__nand2_1
XFILLER_160_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20314__C _20314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22065_ _22064_/A _22064_/B _22064_/C _22064_/D vssd1 vssd1 vccd1 vccd1 _22135_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11524__C1 _18482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18610__A2_N _11879_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21016_ _21046_/A _21046_/B vssd1 vssd1 vccd1 vccd1 _21021_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21051__A2 _21017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20611__A _20611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18288__A _18288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15805__A2 _17427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22000__A1 _21841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22967_ _22968_/CLK _22967_/D vssd1 vssd1 vccd1 vccd1 _22967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_810 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22896__CLK _22952_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12720_ _20255_/B vssd1 vssd1 vccd1 vccd1 _12721_/A sky130_fd_sc_hd__buf_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21918_ _21917_/Y _21836_/Y _21915_/Y vssd1 vssd1 vccd1 vccd1 _21918_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22898_ _22951_/CLK _22898_/D vssd1 vssd1 vccd1 vccd1 _22898_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ _12651_/A _12651_/B _12651_/C vssd1 vssd1 vccd1 vccd1 _12898_/B sky130_fd_sc_hd__nand3_2
XFILLER_130_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21849_ _21610_/B _21740_/X _21848_/X _21742_/Y vssd1 vssd1 vccd1 vccd1 _21857_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_169_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11602_ _11459_/A _11459_/B _11778_/A _11778_/B vssd1 vssd1 vccd1 vccd1 _12003_/C
+ sky130_fd_sc_hd__a22oi_4
XFILLER_90_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15370_ _15370_/A _15370_/B _16322_/B vssd1 vssd1 vccd1 vccd1 _17424_/A sky130_fd_sc_hd__nand3_2
X_12582_ _15299_/C _15299_/D _12683_/A vssd1 vssd1 vccd1 vccd1 _12583_/C sky130_fd_sc_hd__and3_1
XFILLER_196_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14321_ _22586_/D input26/X _22586_/B vssd1 vssd1 vccd1 vccd1 _14413_/A sky130_fd_sc_hd__and3b_1
XFILLER_157_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11533_ _11533_/A _11533_/B vssd1 vssd1 vccd1 vccd1 _11536_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17040_ _17040_/A _17208_/A _17040_/C vssd1 vssd1 vccd1 vccd1 _17208_/B sky130_fd_sc_hd__nand3_4
XFILLER_156_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11464_ _11464_/A vssd1 vssd1 vccd1 vccd1 _15776_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11399__B _16308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14252_ _14153_/A _14285_/C _14248_/B _14248_/A vssd1 vssd1 vccd1 vccd1 _14253_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_171_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11358__A2 _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13203_ _21185_/A _13067_/A _13202_/Y vssd1 vssd1 vccd1 vccd1 _13517_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__12555__B2 _22824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14183_ _14117_/Y _14120_/Y _14118_/Y vssd1 vssd1 vccd1 vccd1 _14188_/C sky130_fd_sc_hd__a21o_1
X_11395_ _11395_/A _11450_/A vssd1 vssd1 vccd1 vccd1 _11395_/X sky130_fd_sc_hd__or2b_1
XFILLER_124_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16297__A2 _12378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13134_ _13449_/B vssd1 vssd1 vccd1 vccd1 _21367_/B sky130_fd_sc_hd__clkbuf_2
X_18991_ _11541_/X _19313_/A _18696_/X _19156_/D vssd1 vssd1 vccd1 vccd1 _18991_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_174_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ _18061_/B _17942_/B vssd1 vssd1 vccd1 vccd1 _17945_/A sky130_fd_sc_hd__or2_1
XANTENNA__19582__A _19687_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ _21448_/C _13330_/A vssd1 vssd1 vccd1 vccd1 _21341_/A sky130_fd_sc_hd__nand2_4
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11846__C _15776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ _12089_/A vssd1 vssd1 vccd1 vccd1 _12055_/A sky130_fd_sc_hd__clkbuf_1
X_17873_ _17873_/A vssd1 vssd1 vccd1 vccd1 _19987_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19612_ _19511_/A _19511_/B _19580_/Y vssd1 vssd1 vccd1 vccd1 _19612_/X sky130_fd_sc_hd__a21o_1
X_16824_ _19320_/A vssd1 vssd1 vccd1 vccd1 _18849_/D sky130_fd_sc_hd__buf_4
XFILLER_4_1110 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17533__C _18303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19543_ _19543_/A vssd1 vssd1 vccd1 vccd1 _19543_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16755_ _16753_/A _16753_/B _16733_/Y _16740_/Y _16853_/A vssd1 vssd1 vccd1 vccd1
+ _16866_/D sky130_fd_sc_hd__o221ai_4
XFILLER_111_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13967_ _14583_/C _14583_/D _14583_/B _14383_/A vssd1 vssd1 vccd1 vccd1 _14566_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15706_ _15706_/A _15707_/A vssd1 vssd1 vccd1 vccd1 _15740_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19474_ _19838_/A _17083_/X _19472_/Y _19473_/X vssd1 vssd1 vccd1 vccd1 _19636_/A
+ sky130_fd_sc_hd__o211ai_4
X_12918_ _12710_/Y _12724_/Y _12915_/Y _12917_/Y vssd1 vssd1 vccd1 vccd1 _13002_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_94_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16686_ _16686_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16686_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13898_ _13897_/Y _13849_/C _13963_/C vssd1 vssd1 vccd1 vccd1 _13899_/B sky130_fd_sc_hd__a21o_1
XANTENNA__16221__A2 _15489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18425_ _18773_/A _18774_/A vssd1 vssd1 vccd1 vccd1 _18425_/Y sky130_fd_sc_hd__nand2_1
X_15637_ _15637_/A vssd1 vssd1 vccd1 vccd1 _15938_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1028 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12849_ _12848_/Y _12488_/Y _12506_/Y vssd1 vssd1 vccd1 vccd1 _12851_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__15988__C _16781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14232__A1 _15050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18356_ _18520_/A _18356_/B vssd1 vssd1 vccd1 vccd1 _18356_/Y sky130_fd_sc_hd__nand2_1
X_15568_ _15568_/A _15568_/B vssd1 vssd1 vccd1 vccd1 _15571_/C sky130_fd_sc_hd__nand2_1
XANTENNA__15980__A1 _15797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17307_ _17307_/A _17307_/B _17307_/C vssd1 vssd1 vccd1 vccd1 _17475_/C sky130_fd_sc_hd__nand3_1
XFILLER_187_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14519_ _14498_/Y _14501_/X _14518_/Y vssd1 vssd1 vccd1 vccd1 _14540_/A sky130_fd_sc_hd__o21ai_2
X_18287_ _18194_/Y _18285_/X _18197_/Y _18286_/X vssd1 vssd1 vccd1 vccd1 _18291_/B
+ sky130_fd_sc_hd__a22oi_2
X_15499_ _15567_/A _15571_/A _15567_/B vssd1 vssd1 vccd1 vccd1 _15500_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_784 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17238_ _12379_/A _12379_/B _18203_/C vssd1 vssd1 vccd1 vccd1 _17238_/X sky130_fd_sc_hd__a21o_2
XANTENNA__15732__A1 _15427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17169_ _17169_/A _17169_/B vssd1 vssd1 vccd1 vccd1 _17180_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19474__A2 _17083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20180_ _20165_/A _20165_/B _20165_/C _20179_/X vssd1 vssd1 vccd1 vccd1 _20181_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_89_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19226__A2 _17525_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16460__A2 _15341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22821_ _22929_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _22821_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13045__A _13045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22752_ _22757_/CLK _22752_/D vssd1 vssd1 vccd1 vccd1 _22752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21703_ _21700_/X _21701_/X _21574_/A _21707_/B _21834_/B vssd1 vssd1 vccd1 vccd1
+ _21704_/C sky130_fd_sc_hd__o221ai_2
X_22683_ _22944_/CLK _22683_/D vssd1 vssd1 vccd1 vccd1 _22683_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13026__A2 _13016_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15420__B1 _15415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16356__A _20471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15260__A _15260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21634_ _21449_/B _21629_/Y _21963_/A _21633_/Y _21219_/C vssd1 vssd1 vccd1 vccd1
+ _21635_/D sky130_fd_sc_hd__o2111ai_1
XANTENNA__19162__A1 _15936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21565_ _21565_/A _21565_/B vssd1 vssd1 vccd1 vccd1 _21574_/A sky130_fd_sc_hd__nand2_2
XFILLER_165_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20516_ _20491_/Y _20501_/X _20513_/Y _20515_/X vssd1 vssd1 vccd1 vccd1 _20522_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_181_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21496_ _21496_/A _21607_/A vssd1 vssd1 vccd1 vccd1 _21716_/A sky130_fd_sc_hd__nand2_2
XFILLER_158_1008 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20447_ _20447_/A _20447_/B _20447_/C vssd1 vssd1 vccd1 vccd1 _20447_/Y sky130_fd_sc_hd__nor3_1
XFILLER_118_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15419__B _17131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20378_ _20403_/C _20378_/B vssd1 vssd1 vccd1 vccd1 _20378_/Y sky130_fd_sc_hd__nor2_2
XFILLER_161_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22117_ _22171_/B _22173_/D _22171_/A vssd1 vssd1 vccd1 vccd1 _22119_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22048_ _21939_/A _21939_/B _21946_/Y vssd1 vssd1 vccd1 vccd1 _22048_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_134_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15239__B1 _14990_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15435__A _22957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870_ _14775_/D _14571_/X _14791_/B _22766_/Q _14791_/A vssd1 vssd1 vccd1 vccd1
+ _14871_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13821_ _13821_/A _13821_/B vssd1 vssd1 vccd1 vccd1 _13821_/Y sky130_fd_sc_hd__nor2_2
XFILLER_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15154__B _15154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16540_ _16540_/A _16540_/B vssd1 vssd1 vccd1 vccd1 _16548_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13752_ _14808_/C vssd1 vssd1 vccd1 vccd1 _14892_/A sky130_fd_sc_hd__buf_2
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16739__B1 _16732_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12703_ _12790_/A vssd1 vssd1 vccd1 vccd1 _12716_/A sky130_fd_sc_hd__buf_4
X_16471_ _16471_/A vssd1 vssd1 vccd1 vccd1 _17631_/A sky130_fd_sc_hd__clkbuf_4
X_13683_ _13497_/X _21280_/B _13499_/X vssd1 vssd1 vccd1 vccd1 _13683_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18210_ _18277_/A _18276_/B _18212_/A vssd1 vssd1 vccd1 vccd1 _18232_/A sky130_fd_sc_hd__a21o_1
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15422_ _16477_/C vssd1 vssd1 vccd1 vccd1 _20129_/A sky130_fd_sc_hd__clkbuf_4
X_19190_ _19190_/A _19190_/B _19190_/C vssd1 vssd1 vccd1 vccd1 _19343_/C sky130_fd_sc_hd__nand3_2
X_12634_ _22823_/Q vssd1 vssd1 vccd1 vccd1 _20130_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_169_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19153__A1 _15888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11579__A2 _18663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18141_ _18141_/A _18337_/A vssd1 vssd1 vccd1 vccd1 _18141_/Y sky130_fd_sc_hd__nand2_2
XFILLER_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15353_ _12824_/A _16320_/A _15608_/C _15362_/D vssd1 vssd1 vccd1 vccd1 _15355_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_141_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12565_ _12565_/A vssd1 vssd1 vccd1 vccd1 _15299_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_157_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14304_ input20/X input19/X input22/X input21/X vssd1 vssd1 vccd1 vccd1 _14305_/D
+ sky130_fd_sc_hd__or4_1
X_18072_ _18071_/Y _18067_/A _18063_/X vssd1 vssd1 vccd1 vccd1 _18072_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11516_ _11583_/B vssd1 vssd1 vccd1 vccd1 _18445_/C sky130_fd_sc_hd__buf_2
XFILLER_156_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15284_ _22882_/Q _15284_/B vssd1 vssd1 vccd1 vccd1 _22870_/D sky130_fd_sc_hd__xnor2_1
XFILLER_89_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12496_ _15631_/A _12493_/Y _15306_/C vssd1 vssd1 vccd1 vccd1 _12497_/A sky130_fd_sc_hd__o21ai_1
XFILLER_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17023_ _16732_/A _16732_/B _16738_/X _16736_/Y vssd1 vssd1 vccd1 vccd1 _17023_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__22911__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17097__A _17341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14235_ _14198_/B _14198_/C _14198_/D _14234_/Y vssd1 vssd1 vccd1 vccd1 _14236_/C
+ sky130_fd_sc_hd__a31oi_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11447_ _11713_/B _15435_/B vssd1 vssd1 vccd1 vccd1 _11459_/B sky130_fd_sc_hd__and2_2
XFILLER_172_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11736__C1 _18093_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22460__A1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ _14165_/A _14165_/C _14054_/A vssd1 vssd1 vccd1 vccd1 _14166_/Y sky130_fd_sc_hd__a21oi_1
X_11378_ _11420_/A vssd1 vssd1 vccd1 vccd1 _11378_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_125_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11751__A2 _17422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13117_ _22841_/Q vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__inv_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _19132_/A _19132_/B _19132_/C _18973_/Y vssd1 vssd1 vccd1 vccd1 _19131_/A
+ sky130_fd_sc_hd__a31oi_4
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _14097_/A _14097_/B _14097_/C vssd1 vssd1 vccd1 vccd1 _14103_/C sky130_fd_sc_hd__nand3_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _19839_/B vssd1 vssd1 vccd1 vccd1 _19941_/A sky130_fd_sc_hd__clkbuf_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _22929_/Q _20314_/A vssd1 vssd1 vccd1 vccd1 _22909_/D sky130_fd_sc_hd__xor2_4
XFILLER_113_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20661__A2_N _20551_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17856_ _17779_/X _17787_/A _17858_/A _17778_/A vssd1 vssd1 vccd1 vccd1 _17857_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_22_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16807_ _12378_/B _15631_/X _15690_/X _18093_/C _16450_/B vssd1 vssd1 vccd1 vccd1
+ _16911_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17787_ _17787_/A _17787_/B vssd1 vssd1 vccd1 vccd1 _17799_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18719__A1 _11511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14999_ _14937_/X _14998_/X _14936_/X _14943_/X vssd1 vssd1 vccd1 vccd1 _15001_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA__15650__B1 _15649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17560__A _18659_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19526_ _19532_/A _19538_/B _19514_/X vssd1 vssd1 vccd1 vccd1 _19526_/Y sky130_fd_sc_hd__a21oi_1
X_16738_ _16710_/Y _16711_/Y _16098_/X _16737_/X vssd1 vssd1 vccd1 vccd1 _16738_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18375__B _18387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19457_ _19457_/A vssd1 vssd1 vccd1 vccd1 _19457_/Y sky130_fd_sc_hd__inv_2
X_16669_ _16669_/A vssd1 vssd1 vccd1 vccd1 _17226_/A sky130_fd_sc_hd__buf_2
XANTENNA__14205__A1 _14868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14205__B2 _14861_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18408_ _18559_/A _18408_/B _18408_/C vssd1 vssd1 vccd1 vccd1 _18408_/X sky130_fd_sc_hd__and3_1
X_19388_ _19338_/X _19344_/Y _19458_/B _19398_/C _19458_/A vssd1 vssd1 vccd1 vccd1
+ _19394_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19144__A1 _22914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18339_ _18339_/A _18339_/B _18339_/C vssd1 vssd1 vccd1 vccd1 _18340_/B sky130_fd_sc_hd__nand3_4
XANTENNA__13312__B _21480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12209__A _12209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21350_ _21460_/A _21344_/D _21349_/X vssd1 vssd1 vccd1 vccd1 _21509_/A sky130_fd_sc_hd__a21oi_1
XFILLER_147_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15705__A1 _15397_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20301_ _20292_/X _20296_/Y _20549_/A vssd1 vssd1 vccd1 vccd1 _20444_/A sky130_fd_sc_hd__o21ai_2
XFILLER_175_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21281_ _21281_/A _21419_/A _21281_/C vssd1 vssd1 vccd1 vccd1 _21419_/B sky130_fd_sc_hd__nand3_2
XFILLER_163_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20232_ _20232_/A _20236_/C vssd1 vssd1 vccd1 vccd1 _20232_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__22451__A1 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15469__B1 _12606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20163_ _12776_/X _12886_/X _12887_/X vssd1 vssd1 vccd1 vccd1 _20163_/X sky130_fd_sc_hd__o21a_1
XFILLER_130_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20094_ _20084_/Y _20085_/X _20088_/X _20093_/Y vssd1 vssd1 vccd1 vccd1 _20119_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_162_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14692__A1 _14270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16969__B1 _16976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15405__D _15799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22804_ _22804_/CLK _22804_/D vssd1 vssd1 vccd1 vccd1 _22804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20517__A1 _20514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20996_ _20990_/A _20954_/B _20906_/Y vssd1 vssd1 vccd1 vccd1 _21067_/A sky130_fd_sc_hd__a21oi_1
XFILLER_164_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_802 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22735_ _22735_/CLK _22735_/D vssd1 vssd1 vccd1 vccd1 _22735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_982 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21423__C _21560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22666_ _22959_/CLK _22666_/D vssd1 vssd1 vccd1 vccd1 _22666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22934__CLK _22937_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21617_ _21645_/C _21645_/D vssd1 vssd1 vccd1 vccd1 _21763_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19686__A2 _17647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22597_ _11349_/X input61/X _22597_/S vssd1 vssd1 vccd1 vccd1 _22598_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12350_ _20323_/A _15314_/A _20341_/C _20338_/C vssd1 vssd1 vccd1 vccd1 _12350_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_139_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21548_ _21548_/A _21548_/B vssd1 vssd1 vccd1 vccd1 _21553_/C sky130_fd_sc_hd__nand2_2
XFILLER_5_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11981__A2 _11979_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ _22799_/Q vssd1 vssd1 vccd1 vccd1 _11302_/A sky130_fd_sc_hd__inv_2
XFILLER_181_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12281_ _22690_/Q _22688_/Q _22689_/Q vssd1 vssd1 vccd1 vccd1 _12340_/A sky130_fd_sc_hd__nor3_2
X_21479_ _21466_/B _21482_/B _21486_/A _21478_/X vssd1 vssd1 vccd1 vccd1 _21490_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_135_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14020_ _14021_/A _14021_/B _13891_/A _14021_/D vssd1 vssd1 vccd1 vccd1 _14022_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17645__A _17652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15971_ _15971_/A _15971_/B vssd1 vssd1 vccd1 vccd1 _15971_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17710_ _17800_/D _17800_/A _17607_/X _17709_/Y vssd1 vssd1 vccd1 vccd1 _17721_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20502__C _20502_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14922_ _14923_/B _14923_/A vssd1 vssd1 vccd1 vccd1 _14924_/A sky130_fd_sc_hd__nor2_1
X_18690_ _18690_/A _18690_/B vssd1 vssd1 vccd1 vccd1 _18690_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17641_ _18629_/B vssd1 vssd1 vccd1 vccd1 _18830_/D sky130_fd_sc_hd__buf_2
XANTENNA__17082__C1 _17007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20221__D _20463_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14853_ _14885_/A _14885_/B _14805_/D vssd1 vssd1 vccd1 vccd1 _14883_/A sky130_fd_sc_hd__o21a_1
XFILLER_64_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13804_ _13808_/A _13881_/A vssd1 vssd1 vccd1 vccd1 _13807_/A sky130_fd_sc_hd__nand2_1
XFILLER_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17572_ _17626_/B _17626_/A _17571_/Y vssd1 vssd1 vccd1 vccd1 _17627_/A sky130_fd_sc_hd__o21ai_2
X_14784_ _15115_/A _15115_/B vssd1 vssd1 vccd1 vccd1 _15240_/C sky130_fd_sc_hd__nand2_2
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_10_0_bq_clk_i clkbuf_3_5_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _22959_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_17_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11996_ _11377_/A _18313_/A _18313_/B _12107_/A vssd1 vssd1 vccd1 vccd1 _18140_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_189_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19311_ _18514_/Y _19308_/X _19310_/X vssd1 vssd1 vccd1 vccd1 _19311_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_44_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16523_ _16476_/X _16515_/Y _16513_/X _16479_/X vssd1 vssd1 vccd1 vccd1 _16524_/B
+ sky130_fd_sc_hd__o211ai_1
X_13735_ _22759_/Q vssd1 vssd1 vccd1 vccd1 _13736_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19242_ _19085_/Y _19086_/Y _19240_/Y _19241_/Y vssd1 vssd1 vccd1 vccd1 _19242_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_143_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16454_ _16734_/A _16734_/B _16734_/C vssd1 vssd1 vccd1 vccd1 _16842_/A sky130_fd_sc_hd__nand3_2
XFILLER_43_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15331__C _20133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13666_ _13666_/A _13666_/B _13666_/C vssd1 vssd1 vccd1 vccd1 _13666_/X sky130_fd_sc_hd__and3_1
XFILLER_32_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15405_ _15893_/A _15776_/B _15799_/A _15799_/B vssd1 vssd1 vccd1 vccd1 _15406_/A
+ sky130_fd_sc_hd__nand4_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19173_ _19320_/A _19358_/C _19358_/D vssd1 vssd1 vccd1 vccd1 _19174_/B sky130_fd_sc_hd__and3_1
X_12617_ _12478_/Y _12479_/X _12621_/A vssd1 vssd1 vccd1 vccd1 _12618_/C sky130_fd_sc_hd__o21ai_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16385_ _16384_/X _15681_/C _15687_/Y vssd1 vssd1 vccd1 vccd1 _16386_/C sky130_fd_sc_hd__a21oi_1
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13597_ _13597_/A _13597_/B _13597_/C vssd1 vssd1 vccd1 vccd1 _13627_/B sky130_fd_sc_hd__nand3_2
XFILLER_157_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16724__A _19470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18124_ _12165_/A _18330_/A _18123_/Y vssd1 vssd1 vccd1 vccd1 _18363_/A sky130_fd_sc_hd__o21ai_1
X_15336_ _11415_/A _15718_/A _15329_/A vssd1 vssd1 vccd1 vccd1 _15336_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18885__B1 _18880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12548_ _12548_/A vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__buf_2
XANTENNA__17539__B _18629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18055_ _18055_/A _18055_/B vssd1 vssd1 vccd1 vccd1 _18055_/X sky130_fd_sc_hd__and2_1
XFILLER_129_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11868__A _18459_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16360__A1 _16586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15267_ _14990_/X _15253_/Y _15217_/B _15266_/Y _15260_/A vssd1 vssd1 vccd1 vccd1
+ _15268_/S sky130_fd_sc_hd__a311o_1
XFILLER_145_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12479_ _12479_/A _12479_/B _12543_/A vssd1 vssd1 vccd1 vccd1 _12479_/X sky130_fd_sc_hd__and3_1
XFILLER_172_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16360__B2 _16431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17006_ _17006_/A _17006_/B _17006_/C _17006_/D vssd1 vssd1 vccd1 vccd1 _17006_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_6_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14218_ _14779_/A vssd1 vssd1 vccd1 vccd1 _14276_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11587__B _11790_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15198_ _15210_/B _15197_/X vssd1 vssd1 vccd1 vccd1 _15199_/B sky130_fd_sc_hd__or2b_1
XFILLER_4_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16112__A1 _15901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14149_ _14161_/B _14149_/B _14161_/C vssd1 vssd1 vccd1 vccd1 _14149_/X sky130_fd_sc_hd__and3_1
XANTENNA__16112__B2 _16554_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18957_ _18957_/A _19132_/C _19132_/A vssd1 vssd1 vccd1 vccd1 _19138_/B sky130_fd_sc_hd__nand3_1
XFILLER_141_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17908_ _17919_/C _17908_/B vssd1 vssd1 vccd1 vccd1 _17908_/Y sky130_fd_sc_hd__xnor2_2
X_18888_ _18127_/B _12146_/Y _12148_/Y _18128_/C _18841_/B vssd1 vssd1 vccd1 vccd1
+ _19316_/B sky130_fd_sc_hd__o311a_1
XFILLER_39_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17839_ _19619_/D _17839_/B _17839_/C vssd1 vssd1 vccd1 vccd1 _17839_/X sky130_fd_sc_hd__and3_1
XANTENNA__22400__S _22402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20850_ _20695_/D _20797_/B _20848_/Y vssd1 vssd1 vccd1 vccd1 _20850_/Y sky130_fd_sc_hd__a21oi_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19365__A1 _16940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22957__CLK _22964_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19509_ _19652_/A _19506_/Y _19508_/X vssd1 vssd1 vccd1 vccd1 _19511_/A sky130_fd_sc_hd__o21a_1
XFILLER_35_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20781_ _20781_/A _20781_/B _20972_/D vssd1 vssd1 vccd1 vccd1 _20782_/B sky130_fd_sc_hd__nand3_2
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22520_ _22520_/A vssd1 vssd1 vccd1 vccd1 _22753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22451_ _13202_/A input60/X _22453_/S vssd1 vssd1 vccd1 vccd1 _22452_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21402_ _21390_/Y _21394_/Y _21401_/Y vssd1 vssd1 vccd1 vccd1 _21406_/B sky130_fd_sc_hd__a21o_1
X_22382_ _22439_/S vssd1 vssd1 vccd1 vccd1 _22391_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_191_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17449__B _17523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13952__A3 _13727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21333_ _21333_/A vssd1 vssd1 vccd1 vccd1 _21386_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18891__A3 _18890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18628__B1 _18629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21264_ _21257_/Y _21261_/Y _21263_/Y vssd1 vssd1 vccd1 vccd1 _21264_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22371__A _22439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13993__A _22866_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20215_ _20219_/B _20339_/A _20222_/A vssd1 vssd1 vccd1 vccd1 _20218_/A sky130_fd_sc_hd__o21ai_1
XFILLER_173_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17300__B1 _17304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21195_ _21851_/A _21195_/B _21195_/C _21851_/C vssd1 vssd1 vccd1 vccd1 _21195_/Y
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19840__A2 _17401_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20146_ _20149_/C _20149_/D vssd1 vssd1 vccd1 vccd1 _20147_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20077_ _20077_/A _20077_/B _20080_/A vssd1 vssd1 vccd1 vccd1 _20200_/A sky130_fd_sc_hd__nor3_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18800__B1 _11598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16809__A _19461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _18303_/C vssd1 vssd1 vccd1 vccd1 _12050_/B sky130_fd_sc_hd__buf_2
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18159__A2 _18156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15090__A1 _14990_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _12003_/B vssd1 vssd1 vccd1 vccd1 _11846_/B sky130_fd_sc_hd__clkbuf_4
X_20979_ _21044_/C _20979_/B vssd1 vssd1 vccd1 vccd1 _20980_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13520_ _13520_/A _13520_/B vssd1 vssd1 vccd1 vccd1 _13528_/A sky130_fd_sc_hd__nand2_1
XFILLER_14_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22718_ _22772_/CLK _22718_/D vssd1 vssd1 vccd1 vccd1 _22718_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__20910__A1 _20514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13451_ _13461_/A _13452_/A vssd1 vssd1 vccd1 vccd1 _13516_/D sky130_fd_sc_hd__nand2_1
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16590__A1 _16585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22649_ _22649_/A vssd1 vssd1 vccd1 vccd1 _22811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12402_ _12402_/A vssd1 vssd1 vccd1 vccd1 _15631_/B sky130_fd_sc_hd__buf_2
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16170_ _16174_/A _16111_/B _16111_/A _16118_/C vssd1 vssd1 vccd1 vccd1 _16170_/X
+ sky130_fd_sc_hd__o211a_1
X_13382_ _13384_/A _13381_/Y _13384_/B vssd1 vssd1 vccd1 vccd1 _13382_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12600__B1 _20471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18331__A2 _11988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20674__B1 _20853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15121_ _15120_/C _15120_/A _15120_/B vssd1 vssd1 vccd1 vccd1 _15121_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12333_ _12333_/A _12333_/B vssd1 vssd1 vccd1 vccd1 _12334_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15052_ _15118_/A _15215_/A _15118_/C _15051_/Y vssd1 vssd1 vccd1 vccd1 _15052_/X
+ sky130_fd_sc_hd__a31o_1
X_12264_ _12276_/A _12384_/A _12340_/D vssd1 vssd1 vccd1 vccd1 _12396_/A sky130_fd_sc_hd__nand3_2
XFILLER_181_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12364__C1 _12378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14003_ _14497_/A _14009_/B vssd1 vssd1 vccd1 vccd1 _14007_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18095__A1 _12116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19860_ _19860_/A _19913_/B _19860_/C vssd1 vssd1 vccd1 vccd1 _19860_/Y sky130_fd_sc_hd__nor3_4
X_12195_ _12195_/A vssd1 vssd1 vccd1 vccd1 _18228_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__21609__B _21609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18811_ _12064_/A _16758_/X _18626_/Y vssd1 vssd1 vccd1 vccd1 _18830_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__15448__A3 _12913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput83 _14357_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19791_ _19796_/A _19796_/B _19796_/C vssd1 vssd1 vccd1 vccd1 _19794_/B sky130_fd_sc_hd__nand3_2
Xoutput94 _14400_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17525__D _17525_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15954_ _17882_/C vssd1 vssd1 vccd1 vccd1 _17816_/B sky130_fd_sc_hd__buf_4
X_18742_ _18729_/Y _18730_/Y _18741_/Y _18731_/X vssd1 vssd1 vccd1 vccd1 _18743_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_23_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20729__A1 _20728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20729__B2 _20818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18398__A2 _18407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19595__B2 _17730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14905_ _15188_/B _14619_/X _14722_/Y _14726_/C vssd1 vssd1 vccd1 vccd1 _14905_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18673_ _19351_/A vssd1 vssd1 vccd1 vccd1 _19687_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15885_ _15812_/C _15812_/D _15824_/A _15824_/B vssd1 vssd1 vccd1 vccd1 _15886_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12682__A3 _12680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17624_ _17624_/A _17624_/B vssd1 vssd1 vccd1 vccd1 _17625_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12419__B1 _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14836_ _14836_/A _14836_/B _14836_/C _14836_/D vssd1 vssd1 vccd1 vccd1 _14982_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__21344__B _21848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _17663_/A _17663_/B _17541_/Y _17544_/Y vssd1 vssd1 vccd1 vccd1 _17559_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_17_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14767_ _14731_/A _14731_/C _14731_/B vssd1 vssd1 vccd1 vccd1 _14768_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__17358__B1 _22897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ _11980_/A _18674_/A _11980_/C vssd1 vssd1 vccd1 vccd1 _11979_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__13631__A2 _21489_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16506_ _16506_/A vssd1 vssd1 vccd1 vccd1 _16506_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16157__C _16157_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13718_ _22755_/Q vssd1 vssd1 vccd1 vccd1 _13725_/A sky130_fd_sc_hd__buf_4
XANTENNA__11642__A1 _11635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17486_ _17486_/A _17486_/B _17486_/C vssd1 vssd1 vccd1 vccd1 _17486_/X sky130_fd_sc_hd__and3_1
XANTENNA__15908__A1 _15903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14698_ _14889_/D vssd1 vssd1 vccd1 vccd1 _14951_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16437_ _16669_/A _16670_/A vssd1 vssd1 vccd1 vccd1 _16438_/A sky130_fd_sc_hd__nor2_1
X_19225_ _19037_/C _19224_/X _19037_/B vssd1 vssd1 vccd1 vccd1 _19229_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ _13664_/A _21250_/C _21250_/A _21195_/B _13650_/B vssd1 vssd1 vccd1 vccd1
+ _13649_/X sky130_fd_sc_hd__a32o_1
XFILLER_176_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16581__A1 _16435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19156_ _18984_/Y _19156_/B _19156_/C _19156_/D vssd1 vssd1 vccd1 vccd1 _19156_/Y
+ sky130_fd_sc_hd__nand4b_2
XFILLER_9_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16368_ _16369_/A _16627_/A _16367_/X _15653_/Y vssd1 vssd1 vccd1 vccd1 _16377_/B
+ sky130_fd_sc_hd__o2bb2ai_4
XANTENNA__22654__A1 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18107_ _18107_/A _18107_/B _18107_/C vssd1 vssd1 vccd1 vccd1 _18108_/B sky130_fd_sc_hd__and3_1
XANTENNA__18322__A2 _19322_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15319_ _15329_/A _15319_/B vssd1 vssd1 vccd1 vccd1 _15343_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11598__A _18156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19087_ _19028_/X _19032_/Y _19085_/Y _19086_/Y _19237_/A vssd1 vssd1 vccd1 vccd1
+ _19088_/C sky130_fd_sc_hd__o221ai_2
XANTENNA__16333__A1 _15792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16299_ _16299_/A _20678_/A _20870_/B _18130_/C vssd1 vssd1 vccd1 vccd1 _16299_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_145_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18038_ _18038_/A _18038_/B vssd1 vssd1 vccd1 vccd1 _18065_/B sky130_fd_sc_hd__nand2_1
XFILLER_145_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16884__A2 _17840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20968__A1 _20844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20000_ _19959_/A _19959_/B _19963_/A _19999_/Y vssd1 vssd1 vccd1 vccd1 _20026_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_114_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19989_ _19987_/X _19948_/A _19985_/X _19986_/X vssd1 vssd1 vccd1 vccd1 _20037_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12122__A2 _18848_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21951_ _21952_/C _21952_/A _21952_/B vssd1 vssd1 vccd1 vccd1 _21951_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20196__A2 _20065_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20902_ _20902_/A _20902_/B vssd1 vssd1 vccd1 vccd1 _20902_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21882_ _21882_/A _21882_/B vssd1 vssd1 vccd1 vccd1 _21886_/B sky130_fd_sc_hd__nand2_2
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19338__A1 _19340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20833_ _20907_/A _20906_/B _20994_/A _20832_/Y vssd1 vssd1 vccd1 vccd1 _20833_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_35_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16067__C _19470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18010__B2 _22903_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21696__A2 _21556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20764_ _20764_/A vssd1 vssd1 vccd1 vccd1 _20907_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22366__A _22368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_957 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22503_ _22503_/A vssd1 vssd1 vccd1 vccd1 _22746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16572__A1 _16435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20695_ _20695_/A _20695_/B _20695_/C _20695_/D vssd1 vssd1 vccd1 vccd1 _20796_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_195_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22434_ _22434_/A vssd1 vssd1 vccd1 vccd1 _22716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22365_ _22355_/A _22356_/A _22356_/B _22364_/A vssd1 vssd1 vccd1 vccd1 _22368_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17521__B1 _17523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11301__A _22799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21316_ _21316_/A _21467_/B vssd1 vssd1 vccd1 vccd1 _21320_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22296_ _22297_/A _22297_/B _22295_/Y vssd1 vssd1 vccd1 vccd1 _22298_/A sky130_fd_sc_hd__o21bai_1
XFILLER_11_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21247_ _21247_/A _21247_/B _21247_/C vssd1 vssd1 vccd1 vccd1 _21248_/C sky130_fd_sc_hd__nand3_1
XFILLER_132_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21178_ _13635_/A _21638_/B _21174_/Y _21177_/Y vssd1 vssd1 vccd1 vccd1 _21179_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17923__A _21082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20129_ _20129_/A _20129_/B _20675_/C _20323_/D vssd1 vssd1 vccd1 vccd1 _20129_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13228__A _22848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ _16947_/A vssd1 vssd1 vccd1 vccd1 _16772_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21384__A1 _21383_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20187__A2 _12894_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ _11576_/B _11902_/B _11902_/C vssd1 vssd1 vccd1 vccd1 _11903_/C sky130_fd_sc_hd__nand3b_1
X_15670_ _15666_/A _15668_/X _15673_/B _15673_/C vssd1 vssd1 vccd1 vccd1 _15678_/D
+ sky130_fd_sc_hd__o211ai_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12882_ _12882_/A vssd1 vssd1 vccd1 vccd1 _20182_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16260__B1 _17133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14626_/A _14621_/B _14621_/C _14626_/B vssd1 vssd1 vccd1 vccd1 _14635_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _11833_/A vssd1 vssd1 vccd1 vccd1 _12084_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14810__A1 _13820_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14059__A _22870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17340_ _17330_/Y _17337_/X _17339_/X vssd1 vssd1 vccd1 vccd1 _17340_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11624__A1 _18810_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _15176_/A vssd1 vssd1 vccd1 vccd1 _14552_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11764_/A _11764_/B _12146_/A _12146_/B vssd1 vssd1 vccd1 vccd1 _11995_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_187_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13503_ _13662_/B _13662_/C _13502_/Y vssd1 vssd1 vccd1 vccd1 _13506_/C sky130_fd_sc_hd__a21oi_4
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17271_ _17270_/Y _17180_/B _17168_/B vssd1 vssd1 vccd1 vccd1 _17272_/C sky130_fd_sc_hd__a21boi_1
XFILLER_42_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _14583_/B _13907_/X _13970_/X _14699_/B _14362_/X vssd1 vssd1 vccd1 vccd1
+ _14684_/C sky130_fd_sc_hd__o311ai_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16274__A _16274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11695_ _11689_/Y _11690_/Y _11687_/Y _11643_/Y vssd1 vssd1 vccd1 vccd1 _11696_/B
+ sky130_fd_sc_hd__o211ai_1
X_19010_ _19237_/A vssd1 vssd1 vccd1 vccd1 _19010_/X sky130_fd_sc_hd__clkbuf_2
X_16222_ _15589_/A _16236_/A _16221_/Y vssd1 vssd1 vccd1 vccd1 _16247_/A sky130_fd_sc_hd__o21ai_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13434_ _13434_/A vssd1 vssd1 vccd1 vccd1 _13434_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18304__A2 _18305_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11388__B1 _11404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16153_ _16153_/A _17006_/D _16157_/B vssd1 vssd1 vccd1 vccd1 _16153_/X sky130_fd_sc_hd__and3_1
X_13365_ _22849_/Q vssd1 vssd1 vccd1 vccd1 _21638_/B sky130_fd_sc_hd__buf_2
XFILLER_182_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12307__A _20130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20111__A2 _16779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13129__A1 _13112_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15104_ _15089_/B _15089_/A _15095_/B vssd1 vssd1 vccd1 vccd1 _15135_/A sky130_fd_sc_hd__o21ai_1
XFILLER_142_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_bq_clk_i clkbuf_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14326__B1 _14313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12316_ _12413_/A _12519_/B _12320_/A vssd1 vssd1 vccd1 vccd1 _16266_/A sky130_fd_sc_hd__a21oi_2
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16084_ _16073_/Y _16076_/Y _16056_/Y _16082_/Y _16083_/X vssd1 vssd1 vccd1 vccd1
+ _16084_/Y sky130_fd_sc_hd__a41oi_4
X_13296_ _13302_/A _13295_/X _13243_/A vssd1 vssd1 vccd1 vccd1 _21329_/A sky130_fd_sc_hd__o21ai_2
XFILLER_182_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19912_ _19913_/A _19913_/B _19913_/C vssd1 vssd1 vccd1 vccd1 _19914_/A sky130_fd_sc_hd__o21a_1
XFILLER_142_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15035_ _15035_/A _15035_/B _15035_/C vssd1 vssd1 vccd1 vccd1 _15036_/A sky130_fd_sc_hd__and3_1
XFILLER_142_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12247_ _18272_/A _12247_/B _12247_/C _12247_/D vssd1 vssd1 vccd1 vccd1 _12250_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_123_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19843_ _19909_/A _19909_/B vssd1 vssd1 vccd1 vccd1 _19852_/A sky130_fd_sc_hd__nor2_1
XFILLER_123_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12178_ _12006_/Y _11986_/X _12013_/Y vssd1 vssd1 vccd1 vccd1 _12181_/A sky130_fd_sc_hd__a21boi_1
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17833__A _17833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19774_ _19945_/C _19848_/A _19774_/C _19774_/D vssd1 vssd1 vccd1 vccd1 _19848_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_96_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16986_ _16986_/A _16986_/B vssd1 vssd1 vccd1 vccd1 _16986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18648__B _18648_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18725_ _18725_/A _18741_/C _18741_/D vssd1 vssd1 vccd1 vccd1 _18725_/X sky130_fd_sc_hd__and3_1
XFILLER_67_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15937_ _15932_/X _15792_/C _15792_/A _15935_/X _15936_/X vssd1 vssd1 vccd1 vccd1
+ _15937_/X sky130_fd_sc_hd__o32a_1
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19470__D _19470_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11881__A _18445_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17043__A2 _16884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18367__C _18367_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15868_ _17385_/C vssd1 vssd1 vccd1 vccd1 _17739_/A sky130_fd_sc_hd__buf_2
X_18656_ _15358_/X _19176_/A _18514_/Y _18512_/X _18511_/Y vssd1 vssd1 vccd1 vccd1
+ _18661_/A sky130_fd_sc_hd__o32ai_2
XANTENNA__11863__A1 _11859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17607_ _17607_/A vssd1 vssd1 vccd1 vccd1 _17607_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_184_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14819_ _15188_/B _14619_/X _14722_/Y _14726_/C _14816_/Y vssd1 vssd1 vccd1 vccd1
+ _14821_/B sky130_fd_sc_hd__o311a_1
X_18587_ _18587_/A _18587_/B vssd1 vssd1 vccd1 vccd1 _18960_/C sky130_fd_sc_hd__nand2_2
X_15799_ _15799_/A _15799_/B _16313_/C vssd1 vssd1 vccd1 vccd1 _15975_/B sky130_fd_sc_hd__and3_1
XFILLER_17_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18664__A _19346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17538_ _19507_/C vssd1 vssd1 vccd1 vccd1 _19687_/C sky130_fd_sc_hd__buf_2
XFILLER_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17469_ _17469_/A _17469_/B vssd1 vssd1 vccd1 vccd1 _17470_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20350__A2 _16611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19208_ _19208_/A _19223_/B vssd1 vssd1 vccd1 vccd1 _19208_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20480_ _15938_/A _12928_/A _20476_/Y _20479_/Y vssd1 vssd1 vccd1 vccd1 _20499_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_177_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19139_ _19293_/A _19294_/A _19134_/A _19134_/B _19138_/Y vssd1 vssd1 vccd1 vccd1
+ _19141_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_146_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20102__A2 _20110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16912__A _16912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22150_ _22150_/A _22150_/B _22681_/Q vssd1 vssd1 vccd1 vccd1 _22290_/D sky130_fd_sc_hd__nand3_2
XANTENNA__12591__A2 _12493_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16857__A2 _16594_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21101_ _21138_/B _21115_/B _21066_/X _21079_/Y vssd1 vssd1 vccd1 vccd1 _21122_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15528__A _15528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22081_ _22081_/A _22142_/A vssd1 vssd1 vccd1 vccd1 _22160_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14432__A _14432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16609__A2 _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21032_ _21008_/X _21006_/B _21031_/X vssd1 vssd1 vccd1 vccd1 _21032_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18839__A _19194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16490__B1 _16225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13990__B _14013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16359__A _20854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21934_ _21760_/B _21846_/B _21886_/B vssd1 vssd1 vccd1 vccd1 _21934_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_41_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16078__B _16078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21865_ _21865_/A _21986_/B _21865_/C vssd1 vssd1 vccd1 vccd1 _21891_/B sky130_fd_sc_hd__nand3_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11606__A1 _11285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20816_ _20816_/A _20816_/B vssd1 vssd1 vccd1 vccd1 _20816_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__20326__C1 _17532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21796_ _21899_/A _21802_/C _21799_/B vssd1 vssd1 vccd1 vccd1 _21796_/X sky130_fd_sc_hd__a21o_1
XFILLER_169_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20747_ _20748_/A _20748_/B _20748_/C vssd1 vssd1 vccd1 vccd1 _20751_/A sky130_fd_sc_hd__a21oi_1
XFILLER_169_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14607__A _14611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22675__CLK _22948_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15753__C1 _15727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11480_ _12094_/D vssd1 vssd1 vccd1 vccd1 _18130_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20678_ _20678_/A _20678_/B _20917_/A vssd1 vssd1 vccd1 vccd1 _20678_/Y sky130_fd_sc_hd__nand3_1
XFILLER_11_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18298__A1 _17822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22417_ _22417_/A vssd1 vssd1 vccd1 vccd1 _22708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13150_ _13502_/D vssd1 vssd1 vccd1 vccd1 _21494_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22348_ _22346_/B _22346_/A _22347_/Y vssd1 vssd1 vccd1 vccd1 _22356_/A sky130_fd_sc_hd__a21bo_1
XFILLER_100_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12101_ _12117_/A _12096_/Y _12098_/Y _17280_/A _18453_/C vssd1 vssd1 vccd1 vccd1
+ _12102_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_3_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13081_ _13301_/A _13073_/A _13234_/C _13304_/B vssd1 vssd1 vccd1 vccd1 _21351_/B
+ sky130_fd_sc_hd__o211ai_4
X_22279_ _22259_/X _22202_/A _22278_/Y vssd1 vssd1 vccd1 vccd1 _22317_/B sky130_fd_sc_hd__o21a_1
XFILLER_88_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12032_ _11762_/A _11762_/B _11685_/X vssd1 vssd1 vccd1 vccd1 _12034_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11685__B _18203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14061__B _14491_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16840_ _16840_/A _17189_/A vssd1 vssd1 vccd1 vccd1 _16846_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18470__B2 _18407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19571__C _22918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16771_ _16771_/A vssd1 vssd1 vccd1 vccd1 _17406_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13983_ _22867_/Q vssd1 vssd1 vccd1 vccd1 _14684_/B sky130_fd_sc_hd__buf_2
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15722_ _15649_/X _17108_/B _15959_/A _15721_/Y vssd1 vssd1 vccd1 vccd1 _15727_/A
+ sky130_fd_sc_hd__a22oi_4
X_18510_ _18510_/A vssd1 vssd1 vccd1 vccd1 _19351_/A sky130_fd_sc_hd__buf_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ _15988_/B _16078_/B _15696_/D _20355_/D vssd1 vssd1 vccd1 vccd1 _12934_/X
+ sky130_fd_sc_hd__and4_1
X_19490_ _19490_/A _19490_/B _19490_/C _19490_/D vssd1 vssd1 vccd1 vccd1 _19490_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16233__B1 _16486_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ _18402_/B _18402_/A _18307_/A _18309_/B vssd1 vssd1 vccd1 vccd1 _18443_/A
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ _15636_/Y _15640_/Y _15642_/X vssd1 vssd1 vccd1 vccd1 _15653_/Y sky130_fd_sc_hd__a21oi_4
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12865_ _12455_/Y _12480_/X _12508_/C _12508_/A vssd1 vssd1 vccd1 vccd1 _12865_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__21109__A1 _16585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16784__A1 _16778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _15050_/B _15026_/C _14729_/A _14605_/D vssd1 vssd1 vccd1 vccd1 _14604_/Y
+ sky130_fd_sc_hd__a22oi_1
X_18372_ _11345_/X _11351_/X _16276_/X _11821_/X _18371_/X vssd1 vssd1 vccd1 vccd1
+ _18372_/X sky130_fd_sc_hd__o32a_1
XANTENNA__15901__A _15901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11816_ _11761_/Y _11762_/X _11811_/Y _11815_/Y vssd1 vssd1 vccd1 vccd1 _11816_/Y
+ sky130_fd_sc_hd__o211ai_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15584_ _16241_/C _14430_/A _16241_/D _15536_/A vssd1 vssd1 vccd1 vccd1 _16770_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12792_/A _12792_/B _12794_/X _12795_/Y vssd1 vssd1 vccd1 vccd1 _12796_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17323_/A _17323_/B _17323_/C vssd1 vssd1 vccd1 vccd1 _17324_/C sky130_fd_sc_hd__nand3_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14540_/A _14540_/B _14540_/C vssd1 vssd1 vccd1 vccd1 _14535_/X sky130_fd_sc_hd__and3_1
X_11747_ _11703_/X _11724_/Y _11741_/Y _11746_/Y vssd1 vssd1 vccd1 vccd1 _11762_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17254_ _16040_/A _17391_/A _17257_/A vssd1 vssd1 vccd1 vccd1 _17255_/C sky130_fd_sc_hd__o21ai_1
XFILLER_175_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14466_ _14565_/A _14566_/A vssd1 vssd1 vccd1 vccd1 _14854_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11678_ _11819_/A vssd1 vssd1 vccd1 vccd1 _19316_/A sky130_fd_sc_hd__buf_2
XANTENNA__20883__A3 _15935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16205_ _16209_/A _16403_/A _16402_/B vssd1 vssd1 vccd1 vccd1 _16206_/A sky130_fd_sc_hd__and3_1
XANTENNA__18289__A1 _12116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13417_ _13419_/A _13419_/B vssd1 vssd1 vccd1 vccd1 _13495_/C sky130_fd_sc_hd__xnor2_1
X_17185_ _17331_/A vssd1 vssd1 vccd1 vccd1 _17200_/C sky130_fd_sc_hd__clkbuf_1
X_14397_ _14411_/A vssd1 vssd1 vccd1 vccd1 _14397_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16732__A _16732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16136_ _16126_/A _16126_/B _16126_/C _16122_/Y _15812_/D vssd1 vssd1 vccd1 vccd1
+ _16137_/C sky130_fd_sc_hd__a32oi_4
XANTENNA__13770__A1 _14181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13348_ _21448_/A _21494_/B _21990_/C vssd1 vssd1 vccd1 vccd1 _21216_/A sky130_fd_sc_hd__nand3_2
XFILLER_183_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16451__B _16451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16067_ _19470_/D _16067_/B _19470_/B _16067_/D vssd1 vssd1 vccd1 vccd1 _16067_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_170_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13279_ _13272_/A _13272_/B _13265_/A _13650_/B _13268_/X vssd1 vssd1 vccd1 vccd1
+ _13281_/A sky130_fd_sc_hd__o2111ai_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15018_ _15018_/A _15018_/B _15018_/C vssd1 vssd1 vccd1 vccd1 _15018_/X sky130_fd_sc_hd__and3_1
XFILLER_69_602 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20253__D1 _15991_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19826_ _22921_/Q _19892_/A _19892_/B vssd1 vssd1 vccd1 vccd1 _19890_/B sky130_fd_sc_hd__nand3b_1
XFILLER_64_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14078__A2 _14722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16472__B1 _16772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19757_ _19757_/A _19757_/B vssd1 vssd1 vccd1 vccd1 _19757_/Y sky130_fd_sc_hd__nor2_1
X_16969_ _16040_/A _16799_/X _16941_/X _16976_/B _16934_/X vssd1 vssd1 vccd1 vccd1
+ _16969_/X sky130_fd_sc_hd__o311a_1
XANTENNA__22545__A0 _22765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16179__A _16179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14483__C1 _14362_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17016__A2 _16742_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18708_ _12009_/X _19160_/A _18695_/X _18696_/X _18692_/Y vssd1 vssd1 vccd1 vccd1
+ _18709_/C sky130_fd_sc_hd__o221ai_4
X_19688_ _19585_/D _19689_/A _19689_/B _19689_/D vssd1 vssd1 vccd1 vccd1 _19705_/A
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__12500__A _12500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18639_ _18543_/A _18543_/B _18543_/C _18553_/A _18546_/C vssd1 vssd1 vccd1 vccd1
+ _18933_/C sky130_fd_sc_hd__a32oi_4
XFILLER_25_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20571__A2 _15326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21650_ _21650_/A _21650_/B _21650_/C vssd1 vssd1 vccd1 vccd1 _21650_/X sky130_fd_sc_hd__and3_1
XFILLER_40_719 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20429__A _20843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_888 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18516__A2 _11786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20601_ _20598_/X _20599_/Y _20600_/Y _20484_/Y vssd1 vssd1 vccd1 vccd1 _20603_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_71_1026 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16527__A1 _15545_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21581_ _22734_/Q vssd1 vssd1 vccd1 vccd1 _21582_/C sky130_fd_sc_hd__inv_2
XFILLER_33_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20532_ _20532_/A _20532_/B vssd1 vssd1 vccd1 vccd1 _20568_/B sky130_fd_sc_hd__nand2_1
XFILLER_193_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17738__A _19689_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20463_ _20463_/A _20463_/B _20463_/C vssd1 vssd1 vccd1 vccd1 _20464_/B sky130_fd_sc_hd__nand3_2
XFILLER_146_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16642__A _17806_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22202_ _22202_/A _22201_/Y vssd1 vssd1 vccd1 vccd1 _22258_/B sky130_fd_sc_hd__or2b_2
XFILLER_192_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17457__B _17523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20394_ _20393_/A _20393_/B _20393_/C vssd1 vssd1 vccd1 vccd1 _20395_/B sky130_fd_sc_hd__a21oi_2
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22133_ _22135_/A _22135_/D vssd1 vssd1 vccd1 vccd1 _22134_/B sky130_fd_sc_hd__nand2_1
XFILLER_134_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12316__A2 _12519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22064_ _22064_/A _22064_/B _22064_/C _22064_/D vssd1 vssd1 vccd1 vccd1 _22132_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA__20314__D _20442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11936__D _18093_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11524__B1 _18482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18452__A1 _12018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21015_ _20975_/D _20977_/B _21013_/X vssd1 vssd1 vccd1 vccd1 _21046_/B sky130_fd_sc_hd__a21oi_2
XFILLER_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21051__A3 _21017_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18288__B _19199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_1_0_bq_clk_i_A clkbuf_2_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22536__A0 _22761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21339__B2 _21739_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22000__A2 _21341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22966_ _22968_/CLK _22966_/D vssd1 vssd1 vccd1 vccd1 _22966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21917_ _21917_/A _21917_/B vssd1 vssd1 vccd1 vccd1 _21917_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22897_ _22952_/CLK _22897_/D vssd1 vssd1 vccd1 vccd1 _22897_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_167_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15721__A _16058_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12650_ _12544_/Y _12560_/Y _12562_/X _12510_/A _12510_/B vssd1 vssd1 vccd1 vccd1
+ _12651_/C sky130_fd_sc_hd__o2111ai_2
X_21848_ _21851_/A _21848_/B _21851_/C vssd1 vssd1 vccd1 vccd1 _21848_/X sky130_fd_sc_hd__and3_1
XFILLER_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11601_ _11936_/C vssd1 vssd1 vccd1 vccd1 _18810_/D sky130_fd_sc_hd__buf_4
XFILLER_168_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12581_ _20486_/C _12681_/A _12681_/B _12583_/A _12630_/A vssd1 vssd1 vccd1 vccd1
+ _12584_/A sky130_fd_sc_hd__a32o_1
XANTENNA__14337__A _14351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21779_ _21636_/X _21654_/C _21642_/Y vssd1 vssd1 vccd1 vccd1 _21779_/X sky130_fd_sc_hd__a21o_1
XFILLER_157_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ _14355_/A vssd1 vssd1 vccd1 vccd1 _14320_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13241__A _22847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11532_ _18706_/A _18093_/A _18093_/B vssd1 vssd1 vccd1 vccd1 _11533_/B sky130_fd_sc_hd__and3_1
XFILLER_157_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15726__C1 _15649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14251_ _14248_/A _14248_/B _14248_/C vssd1 vssd1 vccd1 vccd1 _14253_/C sky130_fd_sc_hd__a21bo_1
XFILLER_172_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11463_ _15888_/A vssd1 vssd1 vccd1 vccd1 _17083_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202_ _13202_/A vssd1 vssd1 vccd1 vccd1 _13202_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14182_ _14085_/B _14181_/Y _14143_/X _13924_/A _14120_/Y vssd1 vssd1 vccd1 vccd1
+ _14188_/B sky130_fd_sc_hd__o221ai_4
XFILLER_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11394_ _11394_/A vssd1 vssd1 vccd1 vccd1 _18259_/A sky130_fd_sc_hd__buf_4
XFILLER_192_790 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13133_ _13131_/X _13110_/Y _21580_/A _13055_/A vssd1 vssd1 vccd1 vccd1 _13449_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__20483__D1 _20678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18990_ _18990_/A vssd1 vssd1 vccd1 vccd1 _19185_/A sky130_fd_sc_hd__buf_2
XFILLER_174_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _19987_/D _19987_/A _17981_/D _21081_/B _17940_/B vssd1 vssd1 vccd1 vccd1
+ _17942_/B sky130_fd_sc_hd__o41a_1
XFILLER_155_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _13096_/A _13243_/A _13095_/A vssd1 vssd1 vccd1 vccd1 _13330_/A sky130_fd_sc_hd__a21o_2
XFILLER_155_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11846__D _15776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12015_ _11964_/X _11967_/Y _12007_/Y _12014_/X vssd1 vssd1 vccd1 vccd1 _12089_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_79_966 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17872_ _21083_/A _21083_/B _17872_/C vssd1 vssd1 vccd1 vccd1 _17872_/X sky130_fd_sc_hd__and3_1
XFILLER_94_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19611_ _19580_/Y _19581_/Y _19605_/Y _19610_/Y vssd1 vssd1 vccd1 vccd1 _19611_/X
+ sky130_fd_sc_hd__o211a_1
X_16823_ _16831_/B vssd1 vssd1 vccd1 vccd1 _16828_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13268__B1 _21629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17533__D _18303_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19542_ _19389_/C _19389_/B _19457_/Y vssd1 vssd1 vccd1 vccd1 _19543_/A sky130_fd_sc_hd__a21oi_1
XFILLER_19_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16754_ _16754_/A _16851_/A vssd1 vssd1 vccd1 vccd1 _16866_/C sky130_fd_sc_hd__nand2_1
X_13966_ _22762_/Q vssd1 vssd1 vccd1 vccd1 _14583_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12320__A _12320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15009__A1 _14503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15705_ _15397_/Y _15513_/Y _15700_/C vssd1 vssd1 vccd1 vccd1 _15707_/A sky130_fd_sc_hd__o21ai_1
X_12917_ _12917_/A _12917_/B vssd1 vssd1 vccd1 vccd1 _12917_/Y sky130_fd_sc_hd__nand2_1
X_16685_ _16685_/A _16685_/B _16685_/C vssd1 vssd1 vccd1 vccd1 _16698_/A sky130_fd_sc_hd__nand3_1
X_19473_ _19317_/Y _19330_/B _19479_/B _19479_/C vssd1 vssd1 vccd1 vccd1 _19473_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13897_ _13897_/A _13963_/B _14581_/D _13963_/D vssd1 vssd1 vccd1 vccd1 _13897_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18424_ _18773_/B vssd1 vssd1 vccd1 vccd1 _18774_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15631__A _15631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15636_ _15319_/B _15632_/Y _16720_/C _15634_/Y _20678_/A vssd1 vssd1 vccd1 vccd1
+ _15636_/Y sky130_fd_sc_hd__o2111ai_4
X_12848_ _12848_/A _12848_/B vssd1 vssd1 vccd1 vccd1 _12848_/Y sky130_fd_sc_hd__nand2_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__C1 _13022_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15567_ _15567_/A _15567_/B vssd1 vssd1 vccd1 vccd1 _15571_/B sky130_fd_sc_hd__nand2_1
X_18355_ _18355_/A _18355_/B vssd1 vssd1 vccd1 vccd1 _18356_/B sky130_fd_sc_hd__nand2_1
XANTENNA__15350__B _20605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _12769_/A _12560_/Y _20415_/A _13022_/D vssd1 vssd1 vccd1 vccd1 _12781_/B
+ sky130_fd_sc_hd__a211o_2
XANTENNA__15980__A2 _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19171__A2 _19167_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17306_ _17275_/Y _17285_/Y _17291_/Y _17591_/A vssd1 vssd1 vccd1 vccd1 _17307_/A
+ sky130_fd_sc_hd__o22a_1
X_14518_ _14522_/C _14522_/D vssd1 vssd1 vccd1 vccd1 _14518_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18286_ _15522_/X _15521_/X _18203_/A _15523_/X vssd1 vssd1 vccd1 vccd1 _18286_/X
+ sky130_fd_sc_hd__a211o_1
X_15498_ _15498_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _15571_/A sky130_fd_sc_hd__or2_1
XFILLER_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14449_ _14443_/X _16879_/B _14448_/X vssd1 vssd1 vccd1 vccd1 _22664_/D sky130_fd_sc_hd__a21o_1
XFILLER_175_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17237_ _20608_/A _17631_/A vssd1 vssd1 vccd1 vccd1 _17237_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15732__A2 _16039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19476__C _19476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17168_ _17168_/A _17168_/B vssd1 vssd1 vccd1 vccd1 _17170_/A sky130_fd_sc_hd__nand2_1
XFILLER_162_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16119_ _16047_/A _16047_/B _16047_/C _16047_/D vssd1 vssd1 vccd1 vccd1 _16119_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_142_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17099_ _16920_/Y _16922_/X _16923_/Y _16926_/Y vssd1 vssd1 vccd1 vccd1 _17099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15496__A1 _11721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19226__A3 _18131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15248__A1 _15230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19809_ _19809_/A _19809_/B vssd1 vssd1 vccd1 vccd1 _19811_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13326__A _22844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22820_ _22850_/CLK hold15/X vssd1 vssd1 vccd1 vccd1 _22820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18242__A1_N _12250_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22751_ _22751_/CLK _22751_/D vssd1 vssd1 vccd1 vccd1 _22751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13045__B _13045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21702_ _21815_/B _21702_/B vssd1 vssd1 vccd1 vccd1 _21834_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19013__A _19504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22682_ _22944_/CLK _22682_/D vssd1 vssd1 vccd1 vccd1 _22682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15260__B _15260_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21633_ _21633_/A _21633_/B vssd1 vssd1 vccd1 vccd1 _21633_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_551 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19162__A2 _19517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15708__C1 _15706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21564_ _21424_/A _21285_/C _21288_/Y _21289_/Y vssd1 vssd1 vccd1 vccd1 _21565_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_178_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18571__B _18571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18370__B1 _17427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20515_ _20514_/X _15935_/A _20244_/X _20328_/D _20512_/Y vssd1 vssd1 vccd1 vccd1
+ _20515_/X sky130_fd_sc_hd__o311a_1
XFILLER_154_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16920__A1 _16014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21495_ _21495_/A _21495_/B _21495_/C vssd1 vssd1 vccd1 vccd1 _21607_/A sky130_fd_sc_hd__nand3_1
XFILLER_165_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13195__C1 _21473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20446_ _20446_/A _20446_/B vssd1 vssd1 vccd1 vccd1 _20447_/C sky130_fd_sc_hd__nand2_1
XFILLER_180_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19870__B1 _19836_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20377_ _20362_/Y _20367_/Y _20403_/B vssd1 vssd1 vccd1 vccd1 _20378_/B sky130_fd_sc_hd__o21ai_1
XFILLER_192_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15487__A1 _15539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20480__A1 _15938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22116_ _21964_/X _21970_/X _22105_/X _22044_/A vssd1 vssd1 vccd1 vccd1 _22171_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_161_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22047_ _22039_/Y _22044_/X _22046_/X vssd1 vssd1 vccd1 vccd1 _22047_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22863__CLK _22944_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15435__B _15435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13820_ _13820_/A vssd1 vssd1 vccd1 vccd1 _13820_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13751_ _13984_/C vssd1 vssd1 vccd1 vccd1 _14808_/C sky130_fd_sc_hd__clkbuf_2
X_22949_ _22949_/CLK _22949_/D vssd1 vssd1 vccd1 vccd1 _22949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12702_ _12702_/A vssd1 vssd1 vccd1 vccd1 _12968_/A sky130_fd_sc_hd__buf_2
X_16470_ _17234_/A vssd1 vssd1 vccd1 vccd1 _19351_/B sky130_fd_sc_hd__buf_4
XFILLER_188_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13682_ _21422_/A vssd1 vssd1 vccd1 vccd1 _21424_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__20069__A _20069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15421_ _15703_/B _15703_/A _15420_/Y vssd1 vssd1 vccd1 vccd1 _15707_/B sky130_fd_sc_hd__a21oi_4
X_12633_ _20128_/A vssd1 vssd1 vccd1 vccd1 _20853_/A sky130_fd_sc_hd__buf_2
XFILLER_54_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14067__A _14564_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18140_ _18140_/A _18691_/C _18140_/C vssd1 vssd1 vccd1 vccd1 _18337_/A sky130_fd_sc_hd__nand3_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15352_ _15352_/A vssd1 vssd1 vccd1 vccd1 _20355_/A sky130_fd_sc_hd__buf_4
X_12564_ _12564_/A _12564_/B vssd1 vssd1 vccd1 vccd1 _12755_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303_ input16/X input15/X input18/X input17/X vssd1 vssd1 vccd1 vccd1 _14305_/C
+ sky130_fd_sc_hd__or4_1
X_18071_ _18042_/A _18070_/X _18040_/Y vssd1 vssd1 vccd1 vccd1 _18071_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_157_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11515_ _12090_/A _12090_/B vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__nor2_2
X_15283_ _22881_/Q _15287_/D _15288_/C vssd1 vssd1 vccd1 vccd1 _15284_/B sky130_fd_sc_hd__o21ai_1
XFILLER_89_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16372__C1 _15654_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12495_ _12532_/A vssd1 vssd1 vccd1 vccd1 _15306_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_141_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17022_ _16847_/A _16866_/A _16906_/X vssd1 vssd1 vccd1 vccd1 _17028_/A sky130_fd_sc_hd__a21oi_1
XFILLER_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14234_ _14188_/B _14188_/C _14188_/A vssd1 vssd1 vccd1 vccd1 _14234_/Y sky130_fd_sc_hd__a21oi_1
X_11446_ _22958_/Q vssd1 vssd1 vccd1 vccd1 _15435_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__17097__B _17310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11736__B1 _18093_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14165_ _14165_/A _14165_/B _14165_/C vssd1 vssd1 vccd1 vccd1 _14165_/X sky130_fd_sc_hd__and3_1
XFILLER_166_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11377_ _11377_/A vssd1 vssd1 vccd1 vccd1 _11394_/A sky130_fd_sc_hd__buf_2
XFILLER_152_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15478__A1 _19316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116_ _13330_/A vssd1 vssd1 vccd1 vccd1 _21448_/A sky130_fd_sc_hd__clkbuf_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21628__A _21724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18973_ _18955_/B _18955_/C _18955_/A vssd1 vssd1 vccd1 vccd1 _18973_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_140_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _14099_/B _14099_/C _14096_/C vssd1 vssd1 vccd1 vccd1 _14097_/C sky130_fd_sc_hd__nand3_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _19987_/D _19987_/A _17981_/D _21081_/B vssd1 vssd1 vccd1 vccd1 _17940_/A
+ sky130_fd_sc_hd__or4_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _12754_/X _12894_/Y _13041_/Y _13046_/Y vssd1 vssd1 vccd1 vccd1 _20314_/A
+ sky130_fd_sc_hd__o31a_2
XANTENNA__15626__A _20471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20223__A1 _12450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17855_ _17855_/A _17855_/B vssd1 vssd1 vccd1 vccd1 _17858_/A sky130_fd_sc_hd__or2_1
XFILLER_61_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12688__C _20355_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16806_ _16476_/X _16515_/Y _16513_/X _16479_/X vssd1 vssd1 vccd1 vccd1 _16812_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12050__A _19490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17786_ _17855_/A _17855_/B _17778_/A _17784_/Y _17785_/X vssd1 vssd1 vccd1 vccd1
+ _17787_/B sky130_fd_sc_hd__o311a_1
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14453__A2 _11438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14998_ _14998_/A _15212_/A _14998_/C vssd1 vssd1 vccd1 vccd1 _14998_/X sky130_fd_sc_hd__or3_1
XFILLER_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18719__A2 _18718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19525_ _19525_/A vssd1 vssd1 vccd1 vccd1 _19538_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16737_ _16737_/A vssd1 vssd1 vccd1 vccd1 _16737_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12985__A _15799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ _13949_/A vssd1 vssd1 vccd1 vccd1 _13949_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21723__A1 _21767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18375__C _18387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19456_ _19401_/X _19408_/X _19407_/X vssd1 vssd1 vccd1 vccd1 _19545_/A sky130_fd_sc_hd__a21bo_1
X_16668_ _16665_/X _17065_/A _16660_/Y vssd1 vssd1 vccd1 vccd1 _16675_/A sky130_fd_sc_hd__a21o_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15402__B2 _18512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18407_ _18407_/A _18407_/B vssd1 vssd1 vccd1 vccd1 _18408_/B sky130_fd_sc_hd__nor2_1
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19768__A _19842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15619_ _16715_/A _20098_/D _18876_/C vssd1 vssd1 vccd1 vccd1 _16332_/A sky130_fd_sc_hd__nand3_1
X_19387_ _19530_/B _19530_/C _19385_/Y _19386_/Y vssd1 vssd1 vccd1 vccd1 _19458_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16599_ _16599_/A _16599_/B _16599_/C vssd1 vssd1 vccd1 vccd1 _16602_/C sky130_fd_sc_hd__nand3_2
XFILLER_194_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18338_ _18339_/A _18339_/B _18338_/C vssd1 vssd1 vccd1 vccd1 _18484_/A sky130_fd_sc_hd__nand3_1
XFILLER_175_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16902__A1 _22893_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18269_ _22911_/Q vssd1 vssd1 vccd1 vccd1 _18432_/A sky130_fd_sc_hd__clkinv_2
XFILLER_129_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16192__A _20734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17719__C _17719_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20300_ _20300_/A _20300_/B _20300_/C vssd1 vssd1 vccd1 vccd1 _20549_/A sky130_fd_sc_hd__nand3_1
XFILLER_128_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21280_ _21280_/A _21280_/B vssd1 vssd1 vccd1 vccd1 _21282_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20231_ _20206_/Y _20446_/B _20211_/Y vssd1 vssd1 vccd1 vccd1 _20236_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__16115__C1 _15972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22886__CLK _22952_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15469__A1 _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15469__B2 _12607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20162_ _20162_/A _20167_/C vssd1 vssd1 vccd1 vccd1 _20165_/B sky130_fd_sc_hd__nand2_2
XFILLER_170_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20442__A _20442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20093_ _20093_/A _20093_/B vssd1 vssd1 vccd1 vccd1 _20093_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14692__A2 _15056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16969__A1 _16040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17751__A _19772_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22369__A input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22803_ _22803_/CLK _22803_/D vssd1 vssd1 vccd1 vccd1 _22803_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13652__B1 _21195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20995_ _21006_/A _21006_/B _21007_/C _21007_/B _21066_/A vssd1 vssd1 vccd1 vccd1
+ _20999_/A sky130_fd_sc_hd__a221o_1
XANTENNA__20517__A2 _15934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22734_ _22735_/CLK _22734_/D vssd1 vssd1 vccd1 vccd1 _22734_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17394__A1 _16040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17933__A3 _21044_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22665_ _22959_/CLK _22665_/D vssd1 vssd1 vccd1 vccd1 _22665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21616_ _21607_/X _21742_/A _21944_/A _21730_/A _22031_/A vssd1 vssd1 vccd1 vccd1
+ _21645_/D sky130_fd_sc_hd__o2111ai_2
XFILLER_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22596_ _22596_/A vssd1 vssd1 vccd1 vccd1 _22787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21547_ _21547_/A _21547_/B vssd1 vssd1 vccd1 vccd1 _21548_/B sky130_fd_sc_hd__nor2_1
XANTENNA__18894__B2 _18893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11300_ _11385_/C _11273_/X _11783_/C _11299_/X vssd1 vssd1 vccd1 vccd1 _11308_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_154_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11981__A3 _11980_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12280_ _12606_/A _12607_/A vssd1 vssd1 vccd1 vccd1 _12457_/A sky130_fd_sc_hd__nand2_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21478_ _21478_/A vssd1 vssd1 vccd1 vccd1 _21478_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12915__C1 _12601_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20429_ _20843_/A _20429_/B _20429_/C vssd1 vssd1 vccd1 vccd1 _20429_/X sky130_fd_sc_hd__or3_1
XANTENNA__19844__C _19900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20453__A1 _20723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17645__B _18830_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1069 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15446__A _15528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15970_ _15970_/A _15970_/B vssd1 vssd1 vccd1 vccd1 _15971_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input32_A wb_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14921_ _14921_/A _14921_/B vssd1 vssd1 vccd1 vccd1 _14923_/A sky130_fd_sc_hd__nand2_1
XFILLER_88_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17082__B1 _16098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17640_ _15840_/X _17440_/A _17633_/Y _17637_/Y vssd1 vssd1 vccd1 vccd1 _17661_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14852_ _14884_/B _14884_/C _14884_/A vssd1 vssd1 vccd1 vccd1 _14885_/A sky130_fd_sc_hd__a21oi_1
XFILLER_29_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15632__A1 _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13803_ _13834_/A _13974_/A _14200_/A vssd1 vssd1 vccd1 vccd1 _13881_/A sky130_fd_sc_hd__nand3_2
X_17571_ _17626_/B _17626_/A _17575_/B vssd1 vssd1 vccd1 vccd1 _17571_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14783_ _14861_/A vssd1 vssd1 vccd1 vccd1 _15115_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11995_ _11995_/A _11995_/B vssd1 vssd1 vccd1 vccd1 _12107_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19310_ _16711_/C _19480_/A _19481_/A _19618_/A _19470_/B vssd1 vssd1 vccd1 vccd1
+ _19310_/X sky130_fd_sc_hd__a32o_1
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16522_ _16248_/X _16060_/A _16472_/Y _16474_/Y vssd1 vssd1 vccd1 vccd1 _16524_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_21_1097 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13734_ _13869_/C vssd1 vssd1 vccd1 vccd1 _13736_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_188_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_112 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19241_ _19530_/A _19343_/A _19343_/B _19343_/C vssd1 vssd1 vccd1 vccd1 _19241_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16453_ _11820_/A _15341_/X _16257_/Y _16816_/A _16452_/X vssd1 vssd1 vccd1 vccd1
+ _16734_/C sky130_fd_sc_hd__o221ai_2
X_13665_ _13665_/A _13665_/B _13665_/C _13665_/D vssd1 vssd1 vccd1 vccd1 _13665_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA_repeater171_A _22690_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15331__D _16781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _12606_/X _12607_/X _11462_/A vssd1 vssd1 vccd1 vccd1 _15404_/X sky130_fd_sc_hd__a21o_2
X_12616_ _12456_/Y _12463_/Y _12455_/A vssd1 vssd1 vccd1 vccd1 _12621_/A sky130_fd_sc_hd__o21ai_1
XFILLER_157_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16384_ _15514_/X _15512_/Y _15682_/Y vssd1 vssd1 vccd1 vccd1 _16384_/X sky130_fd_sc_hd__a21o_1
X_19172_ _19016_/Y _19167_/Y _19334_/A vssd1 vssd1 vccd1 vccd1 _19174_/A sky130_fd_sc_hd__o21ai_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13520_/B _13593_/X _13663_/A _13595_/Y vssd1 vssd1 vccd1 vccd1 _13597_/C
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18334__B1 _15358_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16724__B _19470_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11957__B1 _16912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18123_ _19165_/A _19168_/C _18682_/C vssd1 vssd1 vccd1 vccd1 _18123_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__20677__D1 _17131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15335_ _15335_/A vssd1 vssd1 vccd1 vccd1 _15718_/A sky130_fd_sc_hd__buf_2
XANTENNA__20141__B1 _12718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12547_ _12547_/A vssd1 vssd1 vccd1 vccd1 _20514_/A sky130_fd_sc_hd__buf_2
XANTENNA__16345__C1 _20793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17539__C _19687_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14525__A _22874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18054_ _18051_/Y _18077_/A _18053_/Y _18015_/C vssd1 vssd1 vccd1 vccd1 _18057_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11868__B _17085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15266_ _15266_/A _15266_/B vssd1 vssd1 vccd1 vccd1 _15266_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12478_ _12479_/B _12543_/A _12479_/A vssd1 vssd1 vccd1 vccd1 _12478_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16360__A2 _17833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17005_ _17005_/A _17005_/B _17005_/C vssd1 vssd1 vccd1 vccd1 _17006_/C sky130_fd_sc_hd__nand3_2
X_14217_ _14255_/A _14255_/C _14255_/B vssd1 vssd1 vccd1 vccd1 _14256_/A sky130_fd_sc_hd__a21o_1
X_11429_ _11429_/A _11995_/B vssd1 vssd1 vccd1 vccd1 _11608_/A sky130_fd_sc_hd__nand2_2
XANTENNA__12045__A _19197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15197_ _15197_/A _15197_/B _15223_/A vssd1 vssd1 vccd1 vccd1 _15197_/X sky130_fd_sc_hd__or3_2
XFILLER_125_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16648__B1 _16351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148_ _14161_/B _14161_/C _14149_/B vssd1 vssd1 vccd1 vccd1 _14148_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16112__A2 _15901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14123__A1 _13930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18956_ _18958_/B _19132_/B vssd1 vssd1 vccd1 vccd1 _18957_/A sky130_fd_sc_hd__nand2_1
XFILLER_113_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14079_ _14079_/A _14489_/B vssd1 vssd1 vccd1 vccd1 _14083_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15871__A1 _15415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17907_ _17907_/A _17907_/B vssd1 vssd1 vccd1 vccd1 _17959_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18887_ _18887_/A _18887_/B _18887_/C vssd1 vssd1 vccd1 vccd1 _18897_/A sky130_fd_sc_hd__nand3_1
XFILLER_121_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13882__B1 _13823_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17838_ _21011_/A vssd1 vssd1 vccd1 vccd1 _17839_/C sky130_fd_sc_hd__buf_2
XFILLER_67_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21805__B _21805_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14426__A2 _14418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17769_ _17769_/A _17769_/B vssd1 vssd1 vccd1 vccd1 _17769_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13634__B1 _13126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19365__A2 _18718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19508_ _19346_/A _18629_/B _19651_/B _19651_/C vssd1 vssd1 vccd1 vccd1 _19508_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20780_ _21019_/A _21019_/B _20853_/A vssd1 vssd1 vccd1 vccd1 _20780_/Y sky130_fd_sc_hd__nand3_2
XFILLER_23_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19439_ _19439_/A _19439_/B vssd1 vssd1 vccd1 vccd1 _19561_/B sky130_fd_sc_hd__nand2_1
XANTENNA__15387__B1 _15358_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20380__B1 _20398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22450_ _22450_/A vssd1 vssd1 vccd1 vccd1 _22722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21401_ _21547_/B _21401_/B vssd1 vssd1 vccd1 vccd1 _21401_/Y sky130_fd_sc_hd__nor2_2
XFILLER_136_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11412__A2 _16482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22381_ _22381_/A vssd1 vssd1 vccd1 vccd1 _22692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21332_ _21332_/A _21332_/B _21332_/C vssd1 vssd1 vccd1 vccd1 _21333_/A sky130_fd_sc_hd__nand3_1
XFILLER_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19945__B _19945_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18628__A1 _18625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21263_ _13399_/C _21262_/Y _13494_/B _13495_/A vssd1 vssd1 vccd1 vccd1 _21263_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20214_ _20214_/A _20343_/A vssd1 vssd1 vccd1 vccd1 _20222_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21194_ _21495_/C vssd1 vssd1 vccd1 vccd1 _21851_/C sky130_fd_sc_hd__buf_2
XANTENNA__19840__A3 _17401_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20145_ _20143_/Y _20144_/Y _20155_/B vssd1 vssd1 vccd1 vccd1 _20149_/D sky130_fd_sc_hd__o21ai_1
XFILLER_106_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ _12792_/Y _20073_/Y _20075_/X vssd1 vssd1 vccd1 vccd1 _20080_/A sky130_fd_sc_hd__a21oi_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18800__A1 _15530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1097 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3_0_bq_clk_i clkbuf_2_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__16809__B _16809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22901__CLK _22951_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19356__A2 _15840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11945_/A _11777_/Y _11779_/X vssd1 vssd1 vccd1 vccd1 _11809_/A sky130_fd_sc_hd__a21oi_4
XFILLER_26_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20978_ _20977_/A _20977_/B _20977_/C vssd1 vssd1 vccd1 vccd1 _20979_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22717_ _22812_/CLK _22717_/D vssd1 vssd1 vccd1 vccd1 _22717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16825__A _19614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20910__A2 _16746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13450_ _13450_/A _21476_/C _13450_/C vssd1 vssd1 vccd1 vccd1 _13452_/A sky130_fd_sc_hd__nand3_1
X_22648_ _22811_/Q input54/X _22652_/S vssd1 vssd1 vccd1 vccd1 _22649_/A sky130_fd_sc_hd__mux2_1
XANTENNA__22112__A1 _21853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16590__A2 _16585_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ _12401_/A vssd1 vssd1 vccd1 vccd1 _12403_/A sky130_fd_sc_hd__buf_2
XFILLER_16_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16327__C1 _16062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ _21498_/D _21362_/B _21638_/C _21741_/B vssd1 vssd1 vccd1 vccd1 _13381_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_51_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22579_ _22579_/A vssd1 vssd1 vccd1 vccd1 _22780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ _15120_/A _15120_/B _15120_/C vssd1 vssd1 vccd1 vccd1 _15146_/A sky130_fd_sc_hd__nand3_1
XFILLER_51_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12332_ _12577_/A _12576_/A _12802_/C _12418_/A vssd1 vssd1 vccd1 vccd1 _12333_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_154_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_855 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _15064_/C _15114_/B _15154_/D _15118_/A vssd1 vssd1 vccd1 vccd1 _15051_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_182_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17656__A _19768_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ _22691_/Q vssd1 vssd1 vccd1 vccd1 _12340_/D sky130_fd_sc_hd__inv_2
XFILLER_181_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14002_ _14002_/A _14002_/B _14002_/C vssd1 vssd1 vccd1 vccd1 _14002_/X sky130_fd_sc_hd__and3_1
XANTENNA__18095__A2 _12114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12194_ _18214_/A _18214_/B _18214_/C vssd1 vssd1 vccd1 vccd1 _12195_/A sky130_fd_sc_hd__nand3_1
XFILLER_107_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17806__D _17806_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18810_ _18810_/A _19507_/B _19507_/C _18810_/D vssd1 vssd1 vccd1 vccd1 _18828_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_150_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19790_ _19796_/A _19796_/B _19796_/C vssd1 vssd1 vccd1 vccd1 _19790_/Y sky130_fd_sc_hd__a21oi_1
Xoutput84 _14364_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput95 _14402_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_62_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18741_ _18741_/A _18741_/B _18741_/C _18741_/D vssd1 vssd1 vccd1 vccd1 _18741_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_110_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15953_ _17525_/C vssd1 vssd1 vccd1 vccd1 _17882_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_103_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20729__A2 _15903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17391__A _17391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15904__A _15904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14904_ _14904_/A _14904_/B _14930_/B vssd1 vssd1 vccd1 vccd1 _14914_/C sky130_fd_sc_hd__and3_1
X_18672_ _18735_/A _18735_/B vssd1 vssd1 vccd1 vccd1 _18725_/A sky130_fd_sc_hd__nand2_1
X_15884_ _15842_/A _15842_/B _15853_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15945_/B
+ sky130_fd_sc_hd__o22ai_4
X_17623_ _17781_/B vssd1 vssd1 vccd1 vccd1 _17623_/Y sky130_fd_sc_hd__inv_2
X_14835_ _14834_/X _14673_/Y _14828_/Y _14829_/X _14675_/Y vssd1 vssd1 vccd1 vccd1
+ _14836_/D sky130_fd_sc_hd__o2111ai_2
XANTENNA__21344__C _21733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _17541_/Y _17544_/Y _17529_/X _17531_/X vssd1 vssd1 vccd1 vccd1 _17559_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_11978_ _11969_/A _12126_/A _11977_/Y vssd1 vssd1 vccd1 vccd1 _12137_/B sky130_fd_sc_hd__o21ai_1
X_14766_ _14911_/A _15082_/A _14911_/C vssd1 vssd1 vccd1 vccd1 _14768_/A sky130_fd_sc_hd__and3_1
XFILLER_189_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22351__A1 _22338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16505_ _17137_/A vssd1 vssd1 vccd1 vccd1 _16758_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16157__D _16157_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13717_ _13963_/A vssd1 vssd1 vccd1 vccd1 _13897_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17485_ _17485_/A _17485_/B vssd1 vssd1 vccd1 vccd1 _17485_/Y sky130_fd_sc_hd__nand2_1
X_14697_ _14716_/A _14716_/B vssd1 vssd1 vccd1 vccd1 _14710_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11642__A2 _11641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19224_ _18158_/X _19023_/X _19024_/Y _19026_/Y vssd1 vssd1 vccd1 vccd1 _19224_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16436_ _18258_/B _20069_/A vssd1 vssd1 vccd1 vccd1 _16670_/A sky130_fd_sc_hd__nor2_4
XFILLER_158_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13648_ _13647_/B _13647_/C _13647_/A vssd1 vssd1 vccd1 vccd1 _13671_/A sky130_fd_sc_hd__o21ai_1
XFILLER_60_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22103__A1 _13305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16581__A2 _16579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19156_/B _19156_/C _19154_/X _18984_/Y vssd1 vssd1 vccd1 vccd1 _19155_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16367_ _15616_/X _15657_/Y _15658_/Y _15660_/C vssd1 vssd1 vccd1 vccd1 _16367_/X
+ sky130_fd_sc_hd__o211a_1
X_13579_ _13579_/A vssd1 vssd1 vccd1 vccd1 _21445_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18106_ _16921_/X _12116_/X _18096_/Y _18105_/Y vssd1 vssd1 vccd1 vccd1 _18109_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__18322__A3 _16078_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15318_ _15482_/A _11988_/X _11464_/A _12578_/A _17532_/B vssd1 vssd1 vccd1 vccd1
+ _15319_/B sky130_fd_sc_hd__o2111ai_4
XANTENNA__21862__B1 _21376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19086_ _19086_/A _19086_/B vssd1 vssd1 vccd1 vccd1 _19086_/Y sky130_fd_sc_hd__nand2_2
X_16298_ _16450_/C vssd1 vssd1 vccd1 vccd1 _20870_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_173_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16333__A2 _16745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18037_ _18038_/A _18038_/B vssd1 vssd1 vccd1 vccd1 _18039_/A sky130_fd_sc_hd__or2_1
XFILLER_172_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15249_ _15259_/C vssd1 vssd1 vccd1 vccd1 _15249_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16884__A3 _16879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16470__A _17234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20417__A1 _20844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20968__A2 _17928_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12370__A3 _12403_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19988_ _19985_/X _19986_/X _19987_/X _19948_/A vssd1 vssd1 vccd1 vccd1 _19988_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14647__A2 _14181_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18939_ _18933_/X _18646_/X _18937_/Y _18938_/Y _18932_/Y vssd1 vssd1 vccd1 vccd1
+ _18941_/B sky130_fd_sc_hd__o221ai_1
XFILLER_140_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12658__A1 _12742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19035__B2 _19012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22924__CLK _22948_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21950_ _22037_/B _22122_/C _22037_/A vssd1 vssd1 vccd1 vccd1 _21952_/B sky130_fd_sc_hd__and3_1
XFILLER_55_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20901_ _20901_/A _20901_/B vssd1 vssd1 vccd1 vccd1 _20905_/A sky130_fd_sc_hd__nor2_2
XFILLER_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21881_ _21878_/X _21748_/Y _21879_/Y _21880_/Y vssd1 vssd1 vccd1 vccd1 _21882_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__19338__A2 _19340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20832_ _22936_/Q vssd1 vssd1 vccd1 vccd1 _20832_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21551__A _21551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18010__A2 _22904_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20763_ _20834_/A _20835_/A _20827_/D _20762_/Y vssd1 vssd1 vccd1 vccd1 _20776_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_196_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22502_ _22746_/Q input53/X _22508_/S vssd1 vssd1 vccd1 vccd1 _22503_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21270__B _21841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20694_ _20694_/A _20793_/D _20792_/A _20792_/B vssd1 vssd1 vccd1 vccd1 _20695_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_195_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22433_ _22716_/Q input55/X _22435_/S vssd1 vssd1 vccd1 vccd1 _22434_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20105__B1 _20471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22364_ _22364_/A _22364_/B vssd1 vssd1 vccd1 vccd1 _22945_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__17521__A1 _17523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22382__A _22439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21315_ _21851_/A _21315_/B _21851_/C vssd1 vssd1 vccd1 vccd1 _21467_/B sky130_fd_sc_hd__and3_1
XANTENNA__14335__A1 _11349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15532__B1 _12571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14335__B2 _13826_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22295_ _22211_/A _22290_/Y _22253_/A _22294_/Y vssd1 vssd1 vccd1 vccd1 _22295_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_191_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21246_ _21247_/B _21247_/C _21247_/A vssd1 vssd1 vccd1 vccd1 _21248_/B sky130_fd_sc_hd__a21o_1
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21177_ _21177_/A _21713_/C _21713_/A _21177_/D vssd1 vssd1 vccd1 vccd1 _21177_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_89_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20128_ _20128_/A vssd1 vssd1 vccd1 vccd1 _20323_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_133_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12950_ _20390_/C _12950_/B _12950_/C _12981_/D vssd1 vssd1 vccd1 vccd1 _12954_/B
+ sky130_fd_sc_hd__nand4_1
X_20059_ _20059_/A _20059_/B vssd1 vssd1 vccd1 vccd1 _20059_/Y sky130_fd_sc_hd__nor2_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21445__B _22231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21384__A2 _21341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11901_ _11902_/B _11902_/C _11576_/B vssd1 vssd1 vccd1 vccd1 _11903_/B sky130_fd_sc_hd__a21bo_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _12755_/X _12764_/Y _12874_/Y _12880_/Y vssd1 vssd1 vccd1 vccd1 _12882_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20592__B1 _16708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _14942_/A _14619_/X _14494_/B vssd1 vssd1 vccd1 vccd1 _14626_/B sky130_fd_sc_hd__o21ai_1
X_11832_ _11696_/C _11692_/Y _12247_/C _11831_/Y vssd1 vssd1 vccd1 vccd1 _11832_/Y
+ sky130_fd_sc_hd__o211ai_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14271__B1 _14861_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18537__B1 _11561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14551_/A vssd1 vssd1 vccd1 vccd1 _15176_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _22791_/Q _22790_/Q vssd1 vssd1 vccd1 vccd1 _12146_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11624__A2 _18328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21973__A2_N _22176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13517_/A _21495_/B _13517_/C _13502_/D vssd1 vssd1 vccd1 vccd1 _13502_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_14_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _17270_/A _17270_/B vssd1 vssd1 vccd1 vccd1 _17270_/Y sky130_fd_sc_hd__nand2_1
X_14482_ _14571_/A _14775_/A _14775_/C vssd1 vssd1 vccd1 vccd1 _14684_/A sky130_fd_sc_hd__o21ai_4
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11643_/Y _11649_/Y _11687_/Y vssd1 vssd1 vccd1 vccd1 _11696_/A sky130_fd_sc_hd__a21o_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16221_ _12929_/A _15489_/A _16476_/A vssd1 vssd1 vccd1 vccd1 _16221_/Y sky130_fd_sc_hd__o21ai_4
X_13433_ _13438_/A _13438_/B _13433_/C _13433_/D vssd1 vssd1 vccd1 vccd1 _13440_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19156__A_N _18984_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16152_ _15904_/X _15905_/X _12772_/X _12774_/X vssd1 vssd1 vccd1 vccd1 _16157_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__20647__A1 _20452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13364_ _13581_/A _21177_/D vssd1 vssd1 vccd1 vccd1 _13364_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__21844__B1 _22167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14326__A1 _12528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15103_ _15103_/A _15103_/B vssd1 vssd1 vccd1 vccd1 _22680_/D sky130_fd_sc_hd__nor2_1
X_12315_ _22695_/Q vssd1 vssd1 vccd1 vccd1 _12320_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17386__A _19694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16083_ _11561_/X _11563_/X _12765_/X vssd1 vssd1 vccd1 vccd1 _16083_/X sky130_fd_sc_hd__a21o_1
XFILLER_177_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13295_ _21188_/A vssd1 vssd1 vccd1 vccd1 _13295_/X sky130_fd_sc_hd__buf_2
XFILLER_138_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater134_A _22690_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19911_ _19908_/X _19991_/A vssd1 vssd1 vccd1 vccd1 _19913_/C sky130_fd_sc_hd__and2b_1
X_15034_ _15034_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15035_/C sky130_fd_sc_hd__xor2_1
XANTENNA__19265__A1 _11345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12246_ _12246_/A _12246_/B vssd1 vssd1 vccd1 vccd1 _12247_/D sky130_fd_sc_hd__nand2_1
XANTENNA__19265__B2 _12064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22947__CLK _22948_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__D1 _16106_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19842_ _19842_/A _19842_/B _19842_/C _19842_/D vssd1 vssd1 vccd1 vccd1 _19909_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__12726__A1_N _12583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ _12177_/A _12177_/B _12177_/C vssd1 vssd1 vccd1 vccd1 _12182_/C sky130_fd_sc_hd__nand3_2
XFILLER_110_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19017__A1 _11702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19773_ _15840_/A _19517_/A _19624_/A _17636_/A vssd1 vssd1 vccd1 vccd1 _19774_/C
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__17833__B _17833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13138__B _21480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16985_ _16988_/A _16988_/B _17188_/A _16981_/A vssd1 vssd1 vccd1 vccd1 _16989_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12042__B _22658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18724_ _18724_/A vssd1 vssd1 vccd1 vccd1 _18741_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18648__C _19016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15936_ _15936_/A vssd1 vssd1 vccd1 vccd1 _15936_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18367__D _18659_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18655_ _18655_/A vssd1 vssd1 vccd1 vccd1 _19176_/A sky130_fd_sc_hd__buf_2
X_15867_ _20678_/A vssd1 vssd1 vccd1 vccd1 _17385_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__11863__A2 _11861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17606_ _17611_/A _17611_/B vssd1 vssd1 vccd1 vccd1 _17607_/A sky130_fd_sc_hd__nand2_1
XFILLER_91_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14818_ _14818_/A vssd1 vssd1 vccd1 vccd1 _15188_/B sky130_fd_sc_hd__clkbuf_2
X_18586_ _18774_/A _18586_/B _18586_/C vssd1 vssd1 vccd1 vccd1 _18587_/B sky130_fd_sc_hd__nand3_1
XFILLER_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ _12922_/X _15797_/X _15775_/C _15775_/B vssd1 vssd1 vccd1 vccd1 _15801_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_45_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17537_ _17646_/A vssd1 vssd1 vccd1 vccd1 _18629_/B sky130_fd_sc_hd__buf_2
XFILLER_33_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14749_ _14836_/A _14749_/B vssd1 vssd1 vccd1 vccd1 _14751_/A sky130_fd_sc_hd__nand2_1
XFILLER_178_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16465__A _16465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17468_ _17466_/B _17467_/X _17466_/A vssd1 vssd1 vccd1 vccd1 _17469_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14014__B1 _13748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19207_ _19203_/X _19418_/B _19206_/Y vssd1 vssd1 vccd1 vccd1 _19223_/B sky130_fd_sc_hd__a21oi_1
X_16419_ _16419_/A _16421_/C _16419_/C vssd1 vssd1 vccd1 vccd1 _16695_/D sky130_fd_sc_hd__nand3_1
XFILLER_73_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17399_ _17390_/Y _17399_/B _17399_/C vssd1 vssd1 vccd1 vccd1 _17399_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_164_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11402__A _11502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20638__A1 _12606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19138_ _18607_/Y _19138_/B _19138_/C _19138_/D vssd1 vssd1 vccd1 vccd1 _19138_/Y
+ sky130_fd_sc_hd__nand4b_1
XFILLER_145_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20638__B2 _20734_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18700__B1 _19329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19069_ _19149_/A _19149_/B _19149_/C vssd1 vssd1 vccd1 vccd1 _19104_/A sky130_fd_sc_hd__nand3_1
XANTENNA__18830__D _18830_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16857__A3 _16594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15514__B1 _15700_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21100_ _21066_/X _21079_/Y _21115_/B _21138_/B vssd1 vssd1 vccd1 vccd1 _21122_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_191_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22080_ _22080_/A _22080_/B _22080_/C vssd1 vssd1 vccd1 vccd1 _22142_/A sky130_fd_sc_hd__nand3_1
XFILLER_114_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12879__A1 _12876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21031_ _21095_/A _21031_/B vssd1 vssd1 vccd1 vccd1 _21031_/X sky130_fd_sc_hd__and2_1
XANTENNA__16609__A3 _17875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18839__B _18839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17743__B _18305_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16490__A1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15544__A _15838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16490__B2 _16227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19016__A _19016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13990__C _14786_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21933_ _21933_/A _21933_/B vssd1 vssd1 vccd1 vccd1 _21996_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20574__B1 _20728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16078__C _16078_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21864_ _21865_/A _21986_/B _21865_/C vssd1 vssd1 vccd1 vccd1 _21891_/A sky130_fd_sc_hd__a21o_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20815_ _20810_/A _20810_/B _20813_/X vssd1 vssd1 vccd1 vccd1 _20816_/B sky130_fd_sc_hd__a21o_1
XFILLER_179_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11606__A2 _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21795_ _21783_/X _21785_/Y _21789_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _21899_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20746_ _21050_/C _20734_/A _20734_/C _20745_/X vssd1 vssd1 vccd1 vccd1 _20748_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15753__B1 _15727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20677_ _20605_/Y _20782_/A _20913_/A _20676_/Y _17131_/B vssd1 vssd1 vccd1 vccd1
+ _20682_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_195_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11312__A _22968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22416_ _22708_/Q input47/X _22424_/S vssd1 vssd1 vccd1 vccd1 _22417_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18298__A2 _18778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16822__B _16822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19836__D _19836_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15505__B1 _15504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22347_ _22347_/A _22686_/Q vssd1 vssd1 vccd1 vccd1 _22347_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12100_ _11381_/X _11731_/A _12099_/Y vssd1 vssd1 vccd1 vccd1 _12102_/B sky130_fd_sc_hd__o21ai_1
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ _13145_/A vssd1 vssd1 vccd1 vccd1 _13234_/C sky130_fd_sc_hd__buf_2
XFILLER_88_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15438__B _16473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22278_ _22243_/A _22243_/B _22317_/A _22277_/X vssd1 vssd1 vccd1 vccd1 _22278_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_5_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17258__B1 _15538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ _12055_/A _12055_/B _12088_/B vssd1 vssd1 vccd1 vccd1 _12039_/A sky130_fd_sc_hd__a21o_1
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21229_ _13338_/Y _13354_/B _13315_/X vssd1 vssd1 vccd1 vccd1 _21230_/C sky130_fd_sc_hd__a21boi_1
XANTENNA__11685__C _15580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14061__C _14512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22003__B1 _21733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16770_ _16770_/A vssd1 vssd1 vccd1 vccd1 _17405_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12098__A2 _11819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13982_ _22868_/Q vssd1 vssd1 vccd1 vccd1 _14564_/C sky130_fd_sc_hd__buf_2
XFILLER_101_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ _16058_/C _16809_/B _15960_/A _19154_/C vssd1 vssd1 vccd1 vccd1 _15721_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12933_ _12933_/A _12933_/B _12933_/C _12933_/D vssd1 vssd1 vccd1 vccd1 _12957_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18765__A _18765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16233__A1 _16225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18440_ _18438_/Y _18772_/D _18774_/B vssd1 vssd1 vccd1 vccd1 _18440_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _15343_/X _15651_/Y _15636_/Y _15640_/Y vssd1 vssd1 vccd1 vccd1 _15652_/X
+ sky130_fd_sc_hd__o211a_2
XANTENNA__13047__A1 _12754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12864_/A _12864_/B vssd1 vssd1 vccd1 vccd1 _12867_/B sky130_fd_sc_hd__nand2_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16784__A2 _16779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21109__A2 _16585_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14603_ _14892_/A vssd1 vssd1 vccd1 vccd1 _15026_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18371_ _18371_/A vssd1 vssd1 vccd1 vccd1 _18371_/X sky130_fd_sc_hd__buf_2
XANTENNA__15901__B _15901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ _11930_/A _11930_/B _11930_/C vssd1 vssd1 vccd1 vccd1 _11815_/Y sky130_fd_sc_hd__nand3_2
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15583_ _15583_/A _15583_/B _15583_/C vssd1 vssd1 vccd1 vccd1 _15672_/A sky130_fd_sc_hd__nand3_2
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12788_/B _12788_/C _12793_/X vssd1 vssd1 vccd1 vccd1 _12795_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17122_/A _17122_/B _17122_/C _17125_/X vssd1 vssd1 vccd1 vccd1 _17323_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_144_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _11606_/X _11744_/X _11745_/Y vssd1 vssd1 vccd1 vccd1 _11746_/Y sky130_fd_sc_hd__o21ai_1
X_14534_ _14540_/A _14540_/C _14540_/B _14541_/B _14541_/C vssd1 vssd1 vccd1 vccd1
+ _14534_/X sky130_fd_sc_hd__a32o_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19596__A _19842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17253_ _17142_/X _17252_/Y _17247_/A _17145_/B vssd1 vssd1 vccd1 vccd1 _17257_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11677_ _11738_/A _11737_/A _11706_/A vssd1 vssd1 vccd1 vccd1 _11819_/A sky130_fd_sc_hd__o21ai_4
XFILLER_105_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14465_ _14465_/A _14465_/B _14564_/C vssd1 vssd1 vccd1 vccd1 _14568_/A sky130_fd_sc_hd__nand3_4
XFILLER_30_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16204_ _15964_/Y _16038_/B _16657_/C _16203_/Y vssd1 vssd1 vccd1 vccd1 _16204_/Y
+ sky130_fd_sc_hd__o211ai_2
X_13416_ _13416_/A _13416_/B vssd1 vssd1 vccd1 vccd1 _13419_/B sky130_fd_sc_hd__nor2_1
X_17184_ _17184_/A _17184_/B _17184_/C vssd1 vssd1 vccd1 vccd1 _17331_/A sky130_fd_sc_hd__nand3_1
XANTENNA__18289__A2 _16248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14396_ _14410_/A vssd1 vssd1 vccd1 vccd1 _14396_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16732__B _16732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21293__A1 _22672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16135_ _15824_/C _16017_/X _16093_/B _16093_/A vssd1 vssd1 vccd1 vccd1 _16137_/B
+ sky130_fd_sc_hd__o211ai_2
X_13347_ _21448_/C vssd1 vssd1 vccd1 vccd1 _21990_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_182_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16066_ _18328_/A vssd1 vssd1 vccd1 vccd1 _19470_/B sky130_fd_sc_hd__buf_4
X_13278_ _13282_/B vssd1 vssd1 vccd1 vccd1 _13413_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_143_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12229_ _12225_/A _12195_/A _12230_/C vssd1 vssd1 vccd1 vccd1 _12231_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13149__A _22845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15017_ _15017_/A _15017_/B vssd1 vssd1 vccd1 vccd1 _15018_/C sky130_fd_sc_hd__nor2_1
XFILLER_130_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12730__B1 _12601_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19825_ _19881_/B _19818_/B _19761_/Y _19750_/X vssd1 vssd1 vccd1 vccd1 _19892_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12988__A _12988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16472__A1 _19351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A _17313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16472__B2 _17631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19756_ _19891_/D _19827_/B vssd1 vssd1 vccd1 vccd1 _19759_/A sky130_fd_sc_hd__nand2_1
X_16968_ _16934_/X _16937_/Y _15840_/A _15934_/A vssd1 vssd1 vccd1 vccd1 _16968_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__22545__A1 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18707_ _18707_/A _18707_/B vssd1 vssd1 vccd1 vccd1 _18709_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15919_ _15919_/A vssd1 vssd1 vccd1 vccd1 _15919_/X sky130_fd_sc_hd__buf_6
X_19687_ _19687_/A _19687_/B _19687_/C _19687_/D vssd1 vssd1 vccd1 vccd1 _19689_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16899_ _22894_/Q _16899_/B _16899_/C vssd1 vssd1 vccd1 vccd1 _16899_/Y sky130_fd_sc_hd__nand3b_2
XANTENNA__18675__A _22798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18638_ _18635_/X _18637_/X _18619_/Y _18835_/A vssd1 vssd1 vccd1 vccd1 _18638_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18569_ _18569_/A _18569_/B _18569_/C vssd1 vssd1 vccd1 vccd1 _18570_/A sky130_fd_sc_hd__nand3_1
XANTENNA__15983__B1 _15810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20429__B _20429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20600_ _20599_/B _20475_/C _20599_/A vssd1 vssd1 vccd1 vccd1 _20600_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21580_ _21580_/A _21580_/B vssd1 vssd1 vccd1 vccd1 _21582_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16527__A2 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1038 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20531_ _20531_/A _20531_/B _20531_/C vssd1 vssd1 vccd1 vccd1 _20653_/A sky130_fd_sc_hd__nand3_2
XFILLER_165_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19477__A1 _15580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20462_ _20462_/A vssd1 vssd1 vccd1 vccd1 _20587_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22201_ _21932_/Y _22200_/Y _22166_/Y _22198_/Y vssd1 vssd1 vccd1 vccd1 _22201_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15539__A _15539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20393_ _20393_/A _20393_/B _20393_/C vssd1 vssd1 vccd1 vccd1 _20395_/A sky130_fd_sc_hd__and3_1
XFILLER_133_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22132_ _22132_/A _22132_/B vssd1 vssd1 vccd1 vccd1 _22135_/D sky130_fd_sc_hd__nand2_1
XFILLER_160_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22660__A _22662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22063_ _22113_/A _22059_/Y _22051_/Y _22054_/Y vssd1 vssd1 vccd1 vccd1 _22064_/D
+ sky130_fd_sc_hd__o211ai_2
XFILLER_102_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18988__B1 _18880_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21587__A2 _13521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21014_ _21082_/A _21010_/X _21044_/B _20975_/D _21013_/X vssd1 vssd1 vccd1 vccd1
+ _21046_/A sky130_fd_sc_hd__o311a_1
XANTENNA__18452__A2 _16248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18288__C _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22536__A1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21339__A2 _21725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22965_ _22968_/CLK _22965_/D vssd1 vssd1 vccd1 vccd1 _22965_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_114_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17412__B1 _15355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21916_ _21917_/A _21917_/B _21915_/Y vssd1 vssd1 vccd1 vccd1 _21916_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__13029__A1 _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22896_ _22952_/CLK _22896_/D vssd1 vssd1 vccd1 vccd1 _22896_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17963__A1 _17226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15721__B _16809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21847_ _21847_/A _21847_/B vssd1 vssd1 vccd1 vccd1 _21889_/A sky130_fd_sc_hd__nor2_1
XFILLER_167_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1099 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11600_ _11600_/A _11600_/B _11600_/C vssd1 vssd1 vccd1 vccd1 _11647_/B sky130_fd_sc_hd__nand3_2
XFILLER_24_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12580_ _12576_/X _12577_/X _17532_/A _20101_/C _12579_/X vssd1 vssd1 vccd1 vccd1
+ _12630_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21778_ _21790_/A _21790_/B _21789_/B _21778_/D vssd1 vssd1 vccd1 vccd1 _21781_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_169_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11531_ _11796_/A vssd1 vssd1 vccd1 vccd1 _18706_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11460__B1 _11506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20729_ _20728_/A _15903_/X _20255_/A _20728_/C _20818_/A vssd1 vssd1 vccd1 vccd1
+ _20730_/B sky130_fd_sc_hd__o32a_2
XFILLER_169_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _14250_/A _14250_/B _14250_/C vssd1 vssd1 vccd1 vccd1 _14250_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__19468__A1 _17427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11462_ _11462_/A vssd1 vssd1 vccd1 vccd1 _15888_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16765__A2_N _16496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20355__A _20355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _22723_/Q vssd1 vssd1 vccd1 vccd1 _13202_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1012 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14181_ _14181_/A _14684_/B _14181_/C vssd1 vssd1 vccd1 vccd1 _14181_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__12555__A3 _12567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11393_ _11911_/A _11381_/X _11392_/Y vssd1 vssd1 vccd1 vccd1 _11393_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_152_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13132_ _13145_/A vssd1 vssd1 vccd1 vccd1 _21580_/A sky130_fd_sc_hd__buf_2
XFILLER_48_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input62_A wb_dat_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17940_ _17940_/A _17940_/B vssd1 vssd1 vccd1 vccd1 _18061_/B sky130_fd_sc_hd__nor2_1
XFILLER_151_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _13145_/A vssd1 vssd1 vccd1 vccd1 _13243_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12014_ _12013_/Y _11986_/X _12006_/Y vssd1 vssd1 vccd1 vccd1 _12014_/X sky130_fd_sc_hd__a21o_1
X_17871_ _17871_/A _17897_/A _17871_/C vssd1 vssd1 vccd1 vccd1 _17897_/B sky130_fd_sc_hd__nand3_1
XFILLER_79_978 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19610_ _19610_/A _19610_/B _19610_/C vssd1 vssd1 vccd1 vccd1 _19610_/Y sky130_fd_sc_hd__nand3_1
X_16822_ _16822_/A _16822_/B _16822_/C vssd1 vssd1 vccd1 vccd1 _16831_/B sky130_fd_sc_hd__nand3_1
XFILLER_4_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19541_ _19457_/Y _19389_/X _19650_/A _19540_/Y vssd1 vssd1 vccd1 vccd1 _19545_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_4_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16753_ _16753_/A _16753_/B vssd1 vssd1 vccd1 vccd1 _16851_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13965_ _14581_/B _13973_/A vssd1 vssd1 vccd1 vccd1 _14565_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15704_ _15704_/A _15704_/B vssd1 vssd1 vccd1 vccd1 _15706_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19943__A2 _19461_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19472_ _19168_/Y _19323_/X _19330_/B _19479_/B _19479_/C vssd1 vssd1 vccd1 vccd1
+ _19472_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12916_ _12916_/A _12916_/B vssd1 vssd1 vccd1 vccd1 _12917_/B sky130_fd_sc_hd__nor2_1
XFILLER_185_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16684_ _16438_/A _16426_/X _16664_/B _16664_/C vssd1 vssd1 vccd1 vccd1 _16685_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_111_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13896_ _13896_/A _22759_/Q _22758_/Q vssd1 vssd1 vccd1 vccd1 _14581_/D sky130_fd_sc_hd__nor3_2
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18423_ _18423_/A _18423_/B _18423_/C vssd1 vssd1 vccd1 vccd1 _18773_/B sky130_fd_sc_hd__nand3_1
XFILLER_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15635_ _20355_/A vssd1 vssd1 vccd1 vccd1 _20678_/A sky130_fd_sc_hd__buf_2
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12847_ _12400_/X _20358_/A _20250_/C _20129_/B _12792_/A vssd1 vssd1 vccd1 vccd1
+ _12848_/B sky130_fd_sc_hd__o2111ai_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _18354_/A _18354_/B vssd1 vssd1 vccd1 vccd1 _18520_/A sky130_fd_sc_hd__nand2_2
X_15566_ _15566_/A vssd1 vssd1 vccd1 vccd1 _15566_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15350__C _18876_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12778_ _12968_/D vssd1 vssd1 vccd1 vccd1 _13022_/D sky130_fd_sc_hd__buf_2
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17178_/Y _17172_/A _17181_/Y _17180_/X vssd1 vssd1 vccd1 vccd1 _17475_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_30_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14517_ _14516_/C _14516_/B _14505_/X vssd1 vssd1 vccd1 vccd1 _14522_/D sky130_fd_sc_hd__a21bo_1
XANTENNA__17839__A _19619_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18285_ _11308_/A _11308_/B _15530_/X _15531_/X vssd1 vssd1 vccd1 vccd1 _18285_/X
+ sky130_fd_sc_hd__a22o_1
X_11729_ _16256_/A _16256_/B vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12794__A3 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15497_ _15521_/A _15522_/A _12672_/A _15523_/A vssd1 vssd1 vccd1 vccd1 _15498_/B
+ sky130_fd_sc_hd__a211o_2
XANTENNA__16914__C1 _11666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17236_ _15723_/X _17379_/A _17235_/Y vssd1 vssd1 vccd1 vccd1 _17236_/X sky130_fd_sc_hd__o21a_1
X_14448_ _14448_/A vssd1 vssd1 vccd1 vccd1 _14448_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11887__A _19202_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17167_ _17169_/A _17169_/B _17180_/B _17180_/C vssd1 vssd1 vccd1 vccd1 _17167_/Y
+ sky130_fd_sc_hd__nand4_1
X_14379_ _14410_/A vssd1 vssd1 vccd1 vccd1 _14379_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14263__A _14512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16118_ _16169_/D _16174_/A _16118_/C vssd1 vssd1 vccd1 vccd1 _16186_/A sky130_fd_sc_hd__or3_1
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_964 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17098_ _16919_/A _16919_/B _16919_/C _17095_/X vssd1 vssd1 vccd1 vccd1 _17098_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16049_ _16049_/A vssd1 vssd1 vccd1 vccd1 _16130_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13900__C1 _13815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16445__A1 _16397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22665__CLK _22959_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19808_ _19808_/A _19808_/B vssd1 vssd1 vccd1 vccd1 _19809_/B sky130_fd_sc_hd__and2_1
XANTENNA__14456__B1 _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19739_ _19650_/A _19650_/B _19650_/C _19650_/D _19652_/Y vssd1 vssd1 vccd1 vccd1
+ _19740_/B sky130_fd_sc_hd__a41o_1
XANTENNA__18198__A1 _12050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15822__A _19317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22750_ _22771_/CLK _22750_/D vssd1 vssd1 vccd1 vccd1 _22750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21701_ _21701_/A vssd1 vssd1 vccd1 vccd1 _21701_/X sky130_fd_sc_hd__buf_2
XFILLER_80_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15956__B1 _15955_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22681_ _22944_/CLK _22681_/D vssd1 vssd1 vccd1 vccd1 _22681_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19770__A1_N _19836_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_664 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21632_ _21632_/A vssd1 vssd1 vccd1 vccd1 _21963_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18852__B _18854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_563 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15708__B1 _15700_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21563_ _21566_/A _21566_/B _21930_/A _21562_/Y vssd1 vssd1 vccd1 vccd1 _21568_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_166_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19155__A1_N _19156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18370__A1 _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18370__B2 _12116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18571__C _18571_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20514_ _20514_/A vssd1 vssd1 vccd1 vccd1 _20514_/X sky130_fd_sc_hd__buf_2
XFILLER_165_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21494_ _21851_/A _21494_/B _21495_/C vssd1 vssd1 vccd1 vccd1 _21610_/A sky130_fd_sc_hd__nand3_2
XANTENNA__16920__A2 _17443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20445_ _20549_/B _20549_/D _20422_/Y vssd1 vssd1 vccd1 vccd1 _20445_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_146_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20376_ _20376_/A vssd1 vssd1 vccd1 vccd1 _20403_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15419__D _19154_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22115_ _22115_/A vssd1 vssd1 vccd1 vccd1 _22173_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20480__A2 _12928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15892__C1 _11506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22046_ _21952_/C _21952_/B _22045_/Y vssd1 vssd1 vccd1 vccd1 _22046_/X sky130_fd_sc_hd__a21o_1
XANTENNA__19622__A1 _18107_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20341__C _20341_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14447__B1 _18259_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15435__C _15435_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14462__A3 _14785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13750_ _13750_/A _13750_/B vssd1 vssd1 vccd1 vccd1 _13984_/C sky130_fd_sc_hd__nand2_1
X_22948_ _22948_/CLK _22948_/D vssd1 vssd1 vccd1 vccd1 _22948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17936__B2 _17840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ _12701_/A vssd1 vssd1 vccd1 vccd1 _12702_/A sky130_fd_sc_hd__buf_2
XANTENNA__11681__B1 _11667_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13681_ _21280_/B _13497_/X _13499_/X _13680_/Y vssd1 vssd1 vccd1 vccd1 _21422_/A
+ sky130_fd_sc_hd__o211ai_4
X_22879_ _22944_/CLK input73/X vssd1 vssd1 vccd1 vccd1 _22879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15420_ _15703_/B _15419_/Y _15415_/X vssd1 vssd1 vccd1 vccd1 _15420_/Y sky130_fd_sc_hd__a21oi_1
X_12632_ _15901_/C vssd1 vssd1 vccd1 vccd1 _16498_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_145_1150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15351_ _12009_/A _16300_/A _15350_/Y vssd1 vssd1 vccd1 vccd1 _15368_/A sky130_fd_sc_hd__o21ai_1
X_12563_ _12544_/Y _12560_/Y _12562_/X vssd1 vssd1 vccd1 vccd1 _12564_/B sky130_fd_sc_hd__o21a_1
XFILLER_156_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14302_ input14/X input13/X _14302_/C vssd1 vssd1 vccd1 vccd1 _14305_/B sky130_fd_sc_hd__or3_1
X_11514_ _11551_/B _11551_/C vssd1 vssd1 vccd1 vccd1 _11553_/B sky130_fd_sc_hd__nand2_1
XFILLER_196_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18070_ _17957_/A _17962_/Y _17999_/A vssd1 vssd1 vccd1 vccd1 _18070_/X sky130_fd_sc_hd__o21a_1
XFILLER_141_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12494_ _12288_/A _12401_/A _12385_/A vssd1 vssd1 vccd1 vccd1 _12532_/A sky130_fd_sc_hd__o21ai_2
X_15282_ _15282_/A _15282_/B vssd1 vssd1 vccd1 vccd1 _22869_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17021_ _16906_/X _16907_/Y _17017_/Y _17020_/Y vssd1 vssd1 vccd1 vccd1 _17036_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__22445__A0 _13659_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11445_ _11407_/B _11675_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _11459_/A sky130_fd_sc_hd__nand3b_4
X_14233_ _14238_/A _14238_/B _14233_/C _14233_/D vssd1 vssd1 vccd1 vccd1 _14236_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17097__C _17341_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18113__A1 _18279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11736__A1 _11502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11500__A _18131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ _14248_/A _14248_/C _14248_/B vssd1 vssd1 vccd1 vccd1 _14172_/A sky130_fd_sc_hd__a21boi_1
XFILLER_109_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11376_ _11450_/A _11395_/A _11980_/B _11306_/X vssd1 vssd1 vccd1 vccd1 _11380_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__19861__A1 _19788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15478__A2 _16059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13115_ _13513_/A vssd1 vssd1 vccd1 vccd1 _21362_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18972_ _18972_/A _18972_/B vssd1 vssd1 vccd1 vccd1 _22894_/D sky130_fd_sc_hd__xnor2_1
XFILLER_140_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15907__A _15988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22688__CLK _22690_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14095_ _14178_/B _14093_/Y _14178_/C vssd1 vssd1 vccd1 vccd1 _14097_/B sky130_fd_sc_hd__o21ai_1
XFILLER_140_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17923_ _21082_/C vssd1 vssd1 vccd1 vccd1 _21081_/B sky130_fd_sc_hd__buf_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _12754_/X _12894_/Y _13045_/Y vssd1 vssd1 vccd1 vccd1 _13046_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_79_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18002__B _18044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17854_ _17910_/D _17910_/C _17910_/A _17502_/X vssd1 vssd1 vccd1 vccd1 _17854_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_94_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16805_ _16908_/A _16908_/B _16908_/C vssd1 vssd1 vccd1 vccd1 _17189_/B sky130_fd_sc_hd__nand3_2
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17785_ _17785_/A _17785_/B _17776_/A vssd1 vssd1 vccd1 vccd1 _17785_/X sky130_fd_sc_hd__or3b_4
XFILLER_54_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12050__B _12050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15064__D _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14997_ _14997_/A vssd1 vssd1 vccd1 vccd1 _15212_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19524_ _19510_/Y _19513_/Y _19514_/X _19532_/A vssd1 vssd1 vccd1 vccd1 _19524_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15650__A2 _16397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16736_ _16724_/X _16725_/Y _16743_/C vssd1 vssd1 vccd1 vccd1 _16736_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__21363__B _21629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13948_ _13948_/A vssd1 vssd1 vccd1 vccd1 _13948_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19455_ _19455_/A _19945_/B _19455_/C vssd1 vssd1 vccd1 vccd1 _19455_/X sky130_fd_sc_hd__and3_1
X_16667_ _16667_/A vssd1 vssd1 vccd1 vccd1 _17065_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__21082__C _21082_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ _13881_/A _13986_/A _13873_/X _13877_/Y _14889_/D vssd1 vssd1 vccd1 vccd1
+ _13879_/X sky130_fd_sc_hd__o2111a_1
XANTENNA__18953__A _18953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18406_ _18404_/Y _18405_/X _18396_/Y _18398_/Y vssd1 vssd1 vccd1 vccd1 _18406_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13162__A _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15618_ _15904_/A _15905_/A _15617_/X _12827_/X _20675_/A vssd1 vssd1 vccd1 vccd1
+ _15646_/A sky130_fd_sc_hd__o221ai_4
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19386_ _19386_/A vssd1 vssd1 vccd1 vccd1 _19386_/Y sky130_fd_sc_hd__inv_2
X_16598_ _16598_/A _16598_/B vssd1 vssd1 vccd1 vccd1 _16599_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13287__A1_N _13340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18337_ _18337_/A vssd1 vssd1 vccd1 vccd1 _18337_/X sky130_fd_sc_hd__clkbuf_2
X_15549_ _16964_/A vssd1 vssd1 vccd1 vccd1 _19507_/B sky130_fd_sc_hd__buf_4
XFILLER_148_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18268_ _18268_/A _18268_/B vssd1 vssd1 vccd1 vccd1 _18435_/A sky130_fd_sc_hd__or2_1
XANTENNA__16192__B _16192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13177__B1 _13633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17219_ _17219_/A _17219_/B vssd1 vssd1 vccd1 vccd1 _17220_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_3_5_0_bq_clk_i clkbuf_3_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_bq_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18199_ _11502_/X _11503_/X _19047_/B vssd1 vssd1 vccd1 vccd1 _18199_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_144_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20230_ _20236_/A _20236_/B vssd1 vssd1 vccd1 vccd1 _20232_/A sky130_fd_sc_hd__nand2_1
XANTENNA__20723__A _20723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15469__A2 _11568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20161_ _20200_/A _20161_/B vssd1 vssd1 vccd1 vccd1 _20167_/C sky130_fd_sc_hd__nor2_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14721__A _14892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20092_ _20092_/A _20092_/B _20346_/C vssd1 vssd1 vccd1 vccd1 _20093_/B sky130_fd_sc_hd__and3_2
XFILLER_112_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16969__A2 _16799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21962__A2 _21853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22369__B input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22802_ _22802_/CLK _22802_/D vssd1 vssd1 vccd1 vccd1 _22802_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14492__A2_N _14611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994_ _20994_/A _20994_/B _20906_/C vssd1 vssd1 vccd1 vccd1 _21007_/C sky130_fd_sc_hd__nor3b_1
XFILLER_37_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22733_ _22733_/CLK _22733_/D vssd1 vssd1 vccd1 vccd1 _22733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15271__B _15271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17394__A2 _17393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22664_ _22959_/CLK _22664_/D vssd1 vssd1 vccd1 vccd1 _22664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21615_ _21615_/A vssd1 vssd1 vccd1 vccd1 _22031_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_187_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22595_ _11860_/C input60/X _22597_/S vssd1 vssd1 vccd1 vccd1 _22596_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17146__A2 _17400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15157__A1 _15188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21546_ _21546_/A _21546_/B vssd1 vssd1 vccd1 vccd1 _21548_/A sky130_fd_sc_hd__nand2_1
XFILLER_154_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19694__A _19694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21477_ _21596_/A vssd1 vssd1 vccd1 vccd1 _21486_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12416__A _20130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22830__CLK _22850_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11320__A _11790_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20428_ _20429_/C _20414_/X _20426_/X _20427_/Y _20545_/A vssd1 vssd1 vccd1 vccd1
+ _20431_/B sky130_fd_sc_hd__o221ai_1
XFILLER_175_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17854__B1 _17502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15727__A _15727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20453__A2 _20734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20359_ _20359_/A _20359_/B _20359_/C vssd1 vssd1 vccd1 vccd1 _20359_/X sky130_fd_sc_hd__or3_1
XFILLER_150_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18103__A _18896_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14132__A2 _14191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19056__C1 _19651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22029_ _22029_/A _22029_/B vssd1 vssd1 vccd1 vccd1 _22072_/B sky130_fd_sc_hd__nand2_2
X_14920_ _14919_/A _14919_/B _14919_/C vssd1 vssd1 vccd1 vccd1 _14921_/B sky130_fd_sc_hd__a21o_1
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input25_A wb_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851_ _14825_/C _14902_/B _14825_/A _14826_/A vssd1 vssd1 vccd1 vccd1 _14916_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_91_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15632__A2 _15631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _22867_/Q vssd1 vssd1 vccd1 vccd1 _14200_/A sky130_fd_sc_hd__buf_2
X_17570_ _17442_/X _17439_/X _17564_/A _17433_/B vssd1 vssd1 vccd1 vccd1 _17575_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_95_1100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14782_ _14805_/A _14895_/B vssd1 vssd1 vccd1 vccd1 _14885_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11994_ _12107_/C vssd1 vssd1 vccd1 vccd1 _18313_/B sky130_fd_sc_hd__clkinv_2
XFILLER_95_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16521_ _16535_/A _16535_/B _16534_/B vssd1 vssd1 vccd1 vccd1 _16521_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13733_ _22758_/Q _13733_/B vssd1 vssd1 vccd1 vccd1 _13869_/C sky130_fd_sc_hd__nand2_1
XFILLER_17_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19240_ _19240_/A _19240_/B _19240_/C _19240_/D vssd1 vssd1 vccd1 vccd1 _19240_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_182_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ _16452_/A vssd1 vssd1 vccd1 vccd1 _16452_/X sky130_fd_sc_hd__buf_2
XANTENNA__16593__B1 _16599_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13664_ _13664_/A _13664_/B _21878_/C _13664_/D vssd1 vssd1 vccd1 vccd1 _13665_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_32_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15403_ _15403_/A vssd1 vssd1 vccd1 vccd1 _15403_/X sky130_fd_sc_hd__buf_2
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19171_ _19016_/Y _19167_/Y _19334_/A _19170_/X vssd1 vssd1 vccd1 vccd1 _19171_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12615_ _12456_/Y _12463_/Y _12455_/A _12621_/B vssd1 vssd1 vccd1 vccd1 _12618_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16383_ _16391_/A _16391_/B _16636_/B vssd1 vssd1 vccd1 vccd1 _16386_/B sky130_fd_sc_hd__nand3_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13595_ _13319_/X _13213_/X _13521_/Y vssd1 vssd1 vccd1 vccd1 _13595_/Y sky130_fd_sc_hd__o21ai_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11957__A1 _11502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18122_ _18483_/B vssd1 vssd1 vccd1 vccd1 _19168_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__16724__C _17385_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15334_ _16313_/C vssd1 vssd1 vccd1 vccd1 _16720_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_12_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16345__B1 _15978_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20141__A1 _12721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ _12546_/A vssd1 vssd1 vccd1 vccd1 _12645_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20141__B2 _16708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17539__D _17539_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18053_ _18053_/A _18053_/B _18053_/C vssd1 vssd1 vccd1 vccd1 _18053_/Y sky130_fd_sc_hd__nand3_1
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16896__B2 _16650_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15265_ _14845_/B _15263_/A _15263_/B vssd1 vssd1 vccd1 vccd1 _15265_/X sky130_fd_sc_hd__o21ba_1
XFILLER_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11868__C _16106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ _12500_/A _12501_/A _22822_/Q vssd1 vssd1 vccd1 vccd1 _12479_/A sky130_fd_sc_hd__o21ai_1
XFILLER_138_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16360__A3 _17833_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ _16709_/Y _17081_/A _16554_/C _16994_/Y _17313_/A vssd1 vssd1 vccd1 vccd1
+ _17005_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14216_ _14267_/A _14265_/A _14265_/B _14215_/X vssd1 vssd1 vccd1 vccd1 _14255_/B
+ sky130_fd_sc_hd__a31o_1
X_11428_ _11430_/C _11428_/B _18674_/A vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__18637__A2 _17400_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15196_ _15161_/A _15160_/A _15160_/B _15163_/X vssd1 vssd1 vccd1 vccd1 _15197_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__16648__A1 _16613_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15637__A _15637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ _11593_/A _11594_/A vssd1 vssd1 vccd1 vccd1 _12008_/A sky130_fd_sc_hd__nor2_2
X_14147_ _14147_/A _14147_/B _14147_/C _14147_/D vssd1 vssd1 vccd1 vccd1 _14151_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_180_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16112__A3 _12913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__C1 _15988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14123__A2 _13930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18955_ _18955_/A _18955_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _19132_/B sky130_fd_sc_hd__nand3_2
X_14078_ _14722_/C _14722_/A _14210_/A _14079_/A vssd1 vssd1 vccd1 vccd1 _14082_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17906_ _17919_/C _17908_/B vssd1 vssd1 vccd1 vccd1 _17907_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13029_ _12579_/X _13016_/X _13018_/X vssd1 vssd1 vccd1 vccd1 _13029_/Y sky130_fd_sc_hd__a21oi_1
X_18886_ _18707_/B _18692_/Y _18696_/X _18695_/X vssd1 vssd1 vccd1 vccd1 _18887_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__13882__A1 _13820_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17837_ _21011_/C vssd1 vssd1 vccd1 vccd1 _17839_/B sky130_fd_sc_hd__buf_2
XANTENNA__21805__C _22231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17768_ _17768_/A _17768_/B _17768_/C vssd1 vssd1 vccd1 vccd1 _17769_/B sky130_fd_sc_hd__or3_1
XFILLER_82_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13634__B2 _13434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_642 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19507_ _19507_/A _19507_/B _19507_/C _19507_/D vssd1 vssd1 vccd1 vccd1 _19651_/C
+ sky130_fd_sc_hd__nand4_2
X_16719_ _16719_/A vssd1 vssd1 vccd1 vccd1 _16743_/C sky130_fd_sc_hd__buf_2
XFILLER_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17699_ _17699_/A _17699_/B _17699_/C vssd1 vssd1 vccd1 vccd1 _17701_/B sky130_fd_sc_hd__nand3_1
XFILLER_34_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19438_ _19437_/Y _19427_/C _19428_/A vssd1 vssd1 vccd1 vccd1 _19439_/B sky130_fd_sc_hd__a21boi_2
XANTENNA__15387__A1 _17423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_628 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19369_ _19364_/Y _19365_/X _19366_/Y _19368_/Y vssd1 vssd1 vccd1 vccd1 _19369_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_176_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11354__A_N _11334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1080 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22853__CLK _22937_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21400_ _21399_/B _21399_/C _21689_/A _13361_/X vssd1 vssd1 vccd1 vccd1 _21401_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__20437__B _20554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22380_ _12387_/B input61/X _22380_/S vssd1 vssd1 vccd1 vccd1 _22381_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14435__B _22967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21331_ _21466_/A _21466_/B _21591_/B _21467_/A _21850_/A vssd1 vssd1 vccd1 vccd1
+ _21332_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_175_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1007 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21262_ _13387_/X _13391_/A _13392_/A vssd1 vssd1 vccd1 vccd1 _21262_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_151_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18628__A2 _18627_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20213_ _20213_/A _20213_/B _20338_/C vssd1 vssd1 vccd1 vccd1 _20343_/A sky130_fd_sc_hd__nand3_2
XFILLER_116_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21193_ _21495_/A vssd1 vssd1 vccd1 vccd1 _21851_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20144_ _20132_/X _20142_/B _20137_/X vssd1 vssd1 vccd1 vccd1 _20144_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_77_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20075_ _12525_/A _12525_/B _20415_/A vssd1 vssd1 vccd1 vccd1 _20075_/X sky130_fd_sc_hd__a21o_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21284__A _21423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18800__A2 _15531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16811__A1 _19012_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16809__C _17133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19689__A _19689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ _20977_/A _20977_/B _20977_/C vssd1 vssd1 vccd1 vccd1 _21044_/C sky130_fd_sc_hd__nand3_1
XFILLER_122_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22360__A2 _22338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22716_ _22812_/CLK _22716_/D vssd1 vssd1 vccd1 vccd1 _22716_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19839__D _19839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16825__B _18849_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13389__B1 _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22647_ _22647_/A vssd1 vssd1 vccd1 vccd1 _22810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11939__A1 _12111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12400_ _12606_/A _12607_/A _12574_/A vssd1 vssd1 vccd1 vccd1 _12400_/X sky130_fd_sc_hd__a21o_1
X_13380_ _21609_/B vssd1 vssd1 vccd1 vccd1 _21741_/B sky130_fd_sc_hd__buf_2
XANTENNA__16327__B1 _16996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22578_ _22780_/Q input55/X _22580_/S vssd1 vssd1 vccd1 vccd1 _22579_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12600__A2 _15450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_672 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12331_ _12447_/A _16256_/D _12348_/A vssd1 vssd1 vccd1 vccd1 _12333_/A sky130_fd_sc_hd__nand3_1
X_21529_ _21529_/A _21529_/B _21529_/C vssd1 vssd1 vccd1 vccd1 _21530_/A sky130_fd_sc_hd__nand3_1
XFILLER_166_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15050_ _15050_/A _15050_/B _15050_/C vssd1 vssd1 vccd1 vccd1 _15118_/C sky130_fd_sc_hd__and3_1
X_12262_ _22690_/Q vssd1 vssd1 vccd1 vccd1 _12384_/A sky130_fd_sc_hd__clkinv_2
XFILLER_107_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14001_ _14002_/B _14002_/C _14002_/A vssd1 vssd1 vccd1 vccd1 _14001_/Y sky130_fd_sc_hd__a21oi_1
X_12193_ _12183_/Y _12184_/Y _12182_/C _12182_/D vssd1 vssd1 vccd1 vccd1 _18214_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_134_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15176__B _15180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput85 _14368_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput96 _14405_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[22] sky130_fd_sc_hd__buf_2
XANTENNA__17672__A _17672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18740_ _18666_/X _18664_/X _18827_/A _18826_/A vssd1 vssd1 vccd1 vccd1 _18741_/B
+ sky130_fd_sc_hd__o211ai_1
X_15952_ _15952_/A _15952_/B _15952_/C vssd1 vssd1 vccd1 vccd1 _16034_/A sky130_fd_sc_hd__nand3_1
XFILLER_89_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20729__A3 _20255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14903_ _14904_/B _14930_/B _14904_/A vssd1 vssd1 vccd1 vccd1 _14972_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__18252__B1 _19443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18671_ _18668_/X _18669_/X _18662_/A _18826_/A vssd1 vssd1 vccd1 vccd1 _18735_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_23_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15883_ _15883_/A _15883_/B vssd1 vssd1 vccd1 vccd1 _15883_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17622_ _17622_/A _17622_/B vssd1 vssd1 vccd1 vccd1 _17800_/A sky130_fd_sc_hd__nand2_2
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15605__A2 _16318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14834_ _14834_/A _15186_/D _14834_/C vssd1 vssd1 vccd1 vccd1 _14834_/X sky130_fd_sc_hd__and3_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17553_ _17553_/A vssd1 vssd1 vccd1 vccd1 _17628_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14765_ _14765_/A _14963_/C _14765_/C vssd1 vssd1 vccd1 vccd1 _14769_/A sky130_fd_sc_hd__and3_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ _15904_/A _15905_/A _12127_/A _18325_/A vssd1 vssd1 vccd1 vccd1 _11977_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ _16504_/A vssd1 vssd1 vccd1 vccd1 _16519_/B sky130_fd_sc_hd__inv_2
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22876__CLK _22916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13716_ _22754_/Q _22753_/Q _22752_/Q vssd1 vssd1 vccd1 vccd1 _13963_/A sky130_fd_sc_hd__nor3_4
X_17484_ _17490_/A _17490_/B _17490_/C vssd1 vssd1 vccd1 vccd1 _17484_/X sky130_fd_sc_hd__and3_1
XFILLER_177_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14696_ _14696_/A vssd1 vssd1 vccd1 vccd1 _14716_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19223_ _19223_/A _19223_/B vssd1 vssd1 vccd1 vccd1 _19229_/A sky130_fd_sc_hd__nand2_1
XFILLER_177_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16435_ _18259_/B _16435_/B vssd1 vssd1 vccd1 vccd1 _16669_/A sky130_fd_sc_hd__nor2_4
X_13647_ _13647_/A _13647_/B _13647_/C vssd1 vssd1 vccd1 vccd1 _13647_/Y sky130_fd_sc_hd__nor3_1
XFILLER_108_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22103__A2 _13305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19154_ _19614_/B _19614_/C _19154_/C vssd1 vssd1 vccd1 vccd1 _19154_/X sky130_fd_sc_hd__and3_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16377_/A _16370_/B _16364_/Y _16365_/X vssd1 vssd1 vccd1 vccd1 _16366_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13578_ _13319_/X _13213_/X _13521_/Y _13662_/A _13361_/X vssd1 vssd1 vccd1 vccd1
+ _13578_/X sky130_fd_sc_hd__o32a_1
XANTENNA__21311__B1 _13519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18105_ _19061_/A _18848_/C _19317_/D _18367_/C vssd1 vssd1 vccd1 vccd1 _18105_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_118_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15317_ _12292_/A _15369_/B _12577_/X vssd1 vssd1 vccd1 vccd1 _17532_/B sky130_fd_sc_hd__a21o_4
X_19085_ _19085_/A _19085_/B vssd1 vssd1 vccd1 vccd1 _19085_/Y sky130_fd_sc_hd__nand2_2
XFILLER_118_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21862__A1 _13305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12529_ _12550_/C _12549_/A vssd1 vssd1 vccd1 vccd1 _12773_/A sky130_fd_sc_hd__and2_1
X_16297_ _12403_/D _12378_/A _15981_/X vssd1 vssd1 vccd1 vccd1 _16299_/A sky130_fd_sc_hd__a21oi_1
XFILLER_173_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16751__A _16751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18036_ _18036_/A _18036_/B vssd1 vssd1 vccd1 vccd1 _18038_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15248_ _15230_/A _15247_/A _15246_/X vssd1 vssd1 vccd1 vccd1 _15259_/C sky130_fd_sc_hd__o21ba_2
XFILLER_173_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20417__A2 _15890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__A _11895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _15179_/A vssd1 vssd1 vccd1 vccd1 _22682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19987_ _19987_/A _19987_/B _19987_/C _19987_/D vssd1 vssd1 vccd1 vccd1 _19987_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14647__A3 _14181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18938_ _18938_/A _18938_/B vssd1 vssd1 vccd1 vccd1 _18938_/Y sky130_fd_sc_hd__nand2_1
.ends

