VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bqmain
  CLASS BLOCK ;
  FOREIGN bqmain ;
  ORIGIN 0.000 0.000 ;
  SIZE 554.570 BY 565.290 ;
  PIN bq_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END bq_clk_i
  PIN nreset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 561.290 23.370 565.290 ;
    END
  END nreset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 552.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 552.400 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END wb_adr_i[24]
  PIN wb_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END wb_adr_i[25]
  PIN wb_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END wb_adr_i[26]
  PIN wb_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END wb_adr_i[27]
  PIN wb_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END wb_adr_i[28]
  PIN wb_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END wb_adr_i[29]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END wb_adr_i[30]
  PIN wb_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 4.000 ;
    END
  END wb_adr_i[31]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 4.000 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 0.000 510.050 4.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 4.000 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 0.000 484.750 4.000 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END wb_dat_o[9]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END wb_rst_i
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END wb_we_i
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 23.840 554.570 24.440 ;
    END
  END x[0]
  PIN x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 493.040 554.570 493.640 ;
    END
  END x[10]
  PIN x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 539.960 554.570 540.560 ;
    END
  END x[11]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 70.760 554.570 71.360 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 117.680 554.570 118.280 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 164.600 554.570 165.200 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 211.520 554.570 212.120 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 258.440 554.570 259.040 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 305.360 554.570 305.960 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 352.280 554.570 352.880 ;
    END
  END x[7]
  PIN x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 399.200 554.570 399.800 ;
    END
  END x[8]
  PIN x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.570 446.120 554.570 446.720 ;
    END
  END x[9]
  PIN y[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 561.290 65.690 565.290 ;
    END
  END y[0]
  PIN y[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 561.290 488.890 565.290 ;
    END
  END y[10]
  PIN y[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 561.290 531.210 565.290 ;
    END
  END y[11]
  PIN y[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 561.290 108.010 565.290 ;
    END
  END y[1]
  PIN y[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 561.290 150.330 565.290 ;
    END
  END y[2]
  PIN y[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 561.290 192.650 565.290 ;
    END
  END y[3]
  PIN y[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 561.290 234.970 565.290 ;
    END
  END y[4]
  PIN y[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 561.290 277.290 565.290 ;
    END
  END y[5]
  PIN y[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 561.290 319.610 565.290 ;
    END
  END y[6]
  PIN y[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 561.290 361.930 565.290 ;
    END
  END y[7]
  PIN y[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 561.290 404.250 565.290 ;
    END
  END y[8]
  PIN y[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 561.290 446.570 565.290 ;
    END
  END y[9]
  OBS
      LAYER nwell ;
        RECT 5.330 550.745 548.970 552.350 ;
        RECT 5.330 545.305 548.970 548.135 ;
        RECT 5.330 539.865 548.970 542.695 ;
        RECT 5.330 534.425 548.970 537.255 ;
        RECT 5.330 528.985 548.970 531.815 ;
        RECT 5.330 523.545 548.970 526.375 ;
        RECT 5.330 518.105 548.970 520.935 ;
        RECT 5.330 512.665 548.970 515.495 ;
        RECT 5.330 507.225 548.970 510.055 ;
        RECT 5.330 501.785 548.970 504.615 ;
        RECT 5.330 496.345 548.970 499.175 ;
        RECT 5.330 490.905 548.970 493.735 ;
        RECT 5.330 485.465 548.970 488.295 ;
        RECT 5.330 480.025 548.970 482.855 ;
        RECT 5.330 474.585 548.970 477.415 ;
        RECT 5.330 469.145 548.970 471.975 ;
        RECT 5.330 463.705 548.970 466.535 ;
        RECT 5.330 458.265 548.970 461.095 ;
        RECT 5.330 452.825 548.970 455.655 ;
        RECT 5.330 447.385 548.970 450.215 ;
        RECT 5.330 441.945 548.970 444.775 ;
        RECT 5.330 436.505 548.970 439.335 ;
        RECT 5.330 431.065 548.970 433.895 ;
        RECT 5.330 425.625 548.970 428.455 ;
        RECT 5.330 420.185 548.970 423.015 ;
        RECT 5.330 414.745 548.970 417.575 ;
        RECT 5.330 409.305 548.970 412.135 ;
        RECT 5.330 403.865 548.970 406.695 ;
        RECT 5.330 398.425 548.970 401.255 ;
        RECT 5.330 392.985 548.970 395.815 ;
        RECT 5.330 387.545 548.970 390.375 ;
        RECT 5.330 382.105 548.970 384.935 ;
        RECT 5.330 376.665 548.970 379.495 ;
        RECT 5.330 371.225 548.970 374.055 ;
        RECT 5.330 365.785 548.970 368.615 ;
        RECT 5.330 360.345 548.970 363.175 ;
        RECT 5.330 354.905 548.970 357.735 ;
        RECT 5.330 349.465 548.970 352.295 ;
        RECT 5.330 344.025 548.970 346.855 ;
        RECT 5.330 338.585 548.970 341.415 ;
        RECT 5.330 333.145 548.970 335.975 ;
        RECT 5.330 327.705 548.970 330.535 ;
        RECT 5.330 322.265 548.970 325.095 ;
        RECT 5.330 316.825 548.970 319.655 ;
        RECT 5.330 311.385 548.970 314.215 ;
        RECT 5.330 305.945 548.970 308.775 ;
        RECT 5.330 300.505 548.970 303.335 ;
        RECT 5.330 295.065 548.970 297.895 ;
        RECT 5.330 289.625 548.970 292.455 ;
        RECT 5.330 284.185 548.970 287.015 ;
        RECT 5.330 278.745 548.970 281.575 ;
        RECT 5.330 273.305 548.970 276.135 ;
        RECT 5.330 267.865 548.970 270.695 ;
        RECT 5.330 262.425 548.970 265.255 ;
        RECT 5.330 256.985 548.970 259.815 ;
        RECT 5.330 251.545 548.970 254.375 ;
        RECT 5.330 246.105 548.970 248.935 ;
        RECT 5.330 240.665 548.970 243.495 ;
        RECT 5.330 235.225 548.970 238.055 ;
        RECT 5.330 229.785 548.970 232.615 ;
        RECT 5.330 224.345 548.970 227.175 ;
        RECT 5.330 218.905 548.970 221.735 ;
        RECT 5.330 213.465 548.970 216.295 ;
        RECT 5.330 208.025 548.970 210.855 ;
        RECT 5.330 202.585 548.970 205.415 ;
        RECT 5.330 197.145 548.970 199.975 ;
        RECT 5.330 191.705 548.970 194.535 ;
        RECT 5.330 186.265 548.970 189.095 ;
        RECT 5.330 180.825 548.970 183.655 ;
        RECT 5.330 175.385 548.970 178.215 ;
        RECT 5.330 169.945 548.970 172.775 ;
        RECT 5.330 164.505 548.970 167.335 ;
        RECT 5.330 159.065 548.970 161.895 ;
        RECT 5.330 153.625 548.970 156.455 ;
        RECT 5.330 148.185 548.970 151.015 ;
        RECT 5.330 142.745 548.970 145.575 ;
        RECT 5.330 137.305 548.970 140.135 ;
        RECT 5.330 131.865 548.970 134.695 ;
        RECT 5.330 126.425 548.970 129.255 ;
        RECT 5.330 120.985 548.970 123.815 ;
        RECT 5.330 115.545 548.970 118.375 ;
        RECT 5.330 110.105 548.970 112.935 ;
        RECT 5.330 104.665 548.970 107.495 ;
        RECT 5.330 99.225 548.970 102.055 ;
        RECT 5.330 93.785 548.970 96.615 ;
        RECT 5.330 88.345 548.970 91.175 ;
        RECT 5.330 82.905 548.970 85.735 ;
        RECT 5.330 77.465 548.970 80.295 ;
        RECT 5.330 72.025 548.970 74.855 ;
        RECT 5.330 66.585 548.970 69.415 ;
        RECT 5.330 61.145 548.970 63.975 ;
        RECT 5.330 55.705 548.970 58.535 ;
        RECT 5.330 50.265 548.970 53.095 ;
        RECT 5.330 44.825 548.970 47.655 ;
        RECT 5.330 39.385 548.970 42.215 ;
        RECT 5.330 33.945 548.970 36.775 ;
        RECT 5.330 28.505 548.970 31.335 ;
        RECT 5.330 23.065 548.970 25.895 ;
        RECT 5.330 17.625 548.970 20.455 ;
        RECT 5.330 12.185 548.970 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 548.780 552.245 ;
      LAYER met1 ;
        RECT 5.520 0.040 548.780 552.400 ;
      LAYER met2 ;
        RECT 7.000 561.010 22.810 562.090 ;
        RECT 23.650 561.010 65.130 562.090 ;
        RECT 65.970 561.010 107.450 562.090 ;
        RECT 108.290 561.010 149.770 562.090 ;
        RECT 150.610 561.010 192.090 562.090 ;
        RECT 192.930 561.010 234.410 562.090 ;
        RECT 235.250 561.010 276.730 562.090 ;
        RECT 277.570 561.010 319.050 562.090 ;
        RECT 319.890 561.010 361.370 562.090 ;
        RECT 362.210 561.010 403.690 562.090 ;
        RECT 404.530 561.010 446.010 562.090 ;
        RECT 446.850 561.010 488.330 562.090 ;
        RECT 489.170 561.010 530.650 562.090 ;
        RECT 531.490 561.010 547.300 562.090 ;
        RECT 7.000 4.280 547.300 561.010 ;
        RECT 7.000 0.010 18.670 4.280 ;
        RECT 19.510 0.010 23.730 4.280 ;
        RECT 24.570 0.010 28.790 4.280 ;
        RECT 29.630 0.010 33.850 4.280 ;
        RECT 34.690 0.010 38.910 4.280 ;
        RECT 39.750 0.010 43.970 4.280 ;
        RECT 44.810 0.010 49.030 4.280 ;
        RECT 49.870 0.010 54.090 4.280 ;
        RECT 54.930 0.010 59.150 4.280 ;
        RECT 59.990 0.010 64.210 4.280 ;
        RECT 65.050 0.010 69.270 4.280 ;
        RECT 70.110 0.010 74.330 4.280 ;
        RECT 75.170 0.010 79.390 4.280 ;
        RECT 80.230 0.010 84.450 4.280 ;
        RECT 85.290 0.010 89.510 4.280 ;
        RECT 90.350 0.010 94.570 4.280 ;
        RECT 95.410 0.010 99.630 4.280 ;
        RECT 100.470 0.010 104.690 4.280 ;
        RECT 105.530 0.010 109.750 4.280 ;
        RECT 110.590 0.010 114.810 4.280 ;
        RECT 115.650 0.010 119.870 4.280 ;
        RECT 120.710 0.010 124.930 4.280 ;
        RECT 125.770 0.010 129.990 4.280 ;
        RECT 130.830 0.010 135.050 4.280 ;
        RECT 135.890 0.010 140.110 4.280 ;
        RECT 140.950 0.010 145.170 4.280 ;
        RECT 146.010 0.010 150.230 4.280 ;
        RECT 151.070 0.010 155.290 4.280 ;
        RECT 156.130 0.010 160.350 4.280 ;
        RECT 161.190 0.010 165.410 4.280 ;
        RECT 166.250 0.010 170.470 4.280 ;
        RECT 171.310 0.010 175.530 4.280 ;
        RECT 176.370 0.010 180.590 4.280 ;
        RECT 181.430 0.010 185.650 4.280 ;
        RECT 186.490 0.010 190.710 4.280 ;
        RECT 191.550 0.010 195.770 4.280 ;
        RECT 196.610 0.010 200.830 4.280 ;
        RECT 201.670 0.010 205.890 4.280 ;
        RECT 206.730 0.010 210.950 4.280 ;
        RECT 211.790 0.010 216.010 4.280 ;
        RECT 216.850 0.010 221.070 4.280 ;
        RECT 221.910 0.010 226.130 4.280 ;
        RECT 226.970 0.010 231.190 4.280 ;
        RECT 232.030 0.010 236.250 4.280 ;
        RECT 237.090 0.010 241.310 4.280 ;
        RECT 242.150 0.010 246.370 4.280 ;
        RECT 247.210 0.010 251.430 4.280 ;
        RECT 252.270 0.010 256.490 4.280 ;
        RECT 257.330 0.010 261.550 4.280 ;
        RECT 262.390 0.010 266.610 4.280 ;
        RECT 267.450 0.010 271.670 4.280 ;
        RECT 272.510 0.010 276.730 4.280 ;
        RECT 277.570 0.010 281.790 4.280 ;
        RECT 282.630 0.010 286.850 4.280 ;
        RECT 287.690 0.010 291.910 4.280 ;
        RECT 292.750 0.010 296.970 4.280 ;
        RECT 297.810 0.010 302.030 4.280 ;
        RECT 302.870 0.010 307.090 4.280 ;
        RECT 307.930 0.010 312.150 4.280 ;
        RECT 312.990 0.010 317.210 4.280 ;
        RECT 318.050 0.010 322.270 4.280 ;
        RECT 323.110 0.010 327.330 4.280 ;
        RECT 328.170 0.010 332.390 4.280 ;
        RECT 333.230 0.010 337.450 4.280 ;
        RECT 338.290 0.010 342.510 4.280 ;
        RECT 343.350 0.010 347.570 4.280 ;
        RECT 348.410 0.010 352.630 4.280 ;
        RECT 353.470 0.010 357.690 4.280 ;
        RECT 358.530 0.010 362.750 4.280 ;
        RECT 363.590 0.010 367.810 4.280 ;
        RECT 368.650 0.010 372.870 4.280 ;
        RECT 373.710 0.010 377.930 4.280 ;
        RECT 378.770 0.010 382.990 4.280 ;
        RECT 383.830 0.010 388.050 4.280 ;
        RECT 388.890 0.010 393.110 4.280 ;
        RECT 393.950 0.010 398.170 4.280 ;
        RECT 399.010 0.010 403.230 4.280 ;
        RECT 404.070 0.010 408.290 4.280 ;
        RECT 409.130 0.010 413.350 4.280 ;
        RECT 414.190 0.010 418.410 4.280 ;
        RECT 419.250 0.010 423.470 4.280 ;
        RECT 424.310 0.010 428.530 4.280 ;
        RECT 429.370 0.010 433.590 4.280 ;
        RECT 434.430 0.010 438.650 4.280 ;
        RECT 439.490 0.010 443.710 4.280 ;
        RECT 444.550 0.010 448.770 4.280 ;
        RECT 449.610 0.010 453.830 4.280 ;
        RECT 454.670 0.010 458.890 4.280 ;
        RECT 459.730 0.010 463.950 4.280 ;
        RECT 464.790 0.010 469.010 4.280 ;
        RECT 469.850 0.010 474.070 4.280 ;
        RECT 474.910 0.010 479.130 4.280 ;
        RECT 479.970 0.010 484.190 4.280 ;
        RECT 485.030 0.010 489.250 4.280 ;
        RECT 490.090 0.010 494.310 4.280 ;
        RECT 495.150 0.010 499.370 4.280 ;
        RECT 500.210 0.010 504.430 4.280 ;
        RECT 505.270 0.010 509.490 4.280 ;
        RECT 510.330 0.010 514.550 4.280 ;
        RECT 515.390 0.010 519.610 4.280 ;
        RECT 520.450 0.010 524.670 4.280 ;
        RECT 525.510 0.010 529.730 4.280 ;
        RECT 530.570 0.010 534.790 4.280 ;
        RECT 535.630 0.010 547.300 4.280 ;
      LAYER met3 ;
        RECT 10.185 540.960 550.570 552.325 ;
        RECT 10.185 539.560 550.170 540.960 ;
        RECT 10.185 494.040 550.570 539.560 ;
        RECT 10.185 492.640 550.170 494.040 ;
        RECT 10.185 447.120 550.570 492.640 ;
        RECT 10.185 445.720 550.170 447.120 ;
        RECT 10.185 400.200 550.570 445.720 ;
        RECT 10.185 398.800 550.170 400.200 ;
        RECT 10.185 353.280 550.570 398.800 ;
        RECT 10.185 351.880 550.170 353.280 ;
        RECT 10.185 306.360 550.570 351.880 ;
        RECT 10.185 304.960 550.170 306.360 ;
        RECT 10.185 259.440 550.570 304.960 ;
        RECT 10.185 258.040 550.170 259.440 ;
        RECT 10.185 212.520 550.570 258.040 ;
        RECT 10.185 211.120 550.170 212.520 ;
        RECT 10.185 165.600 550.570 211.120 ;
        RECT 10.185 164.200 550.170 165.600 ;
        RECT 10.185 118.680 550.570 164.200 ;
        RECT 10.185 117.280 550.170 118.680 ;
        RECT 10.185 71.760 550.570 117.280 ;
        RECT 10.185 70.360 550.170 71.760 ;
        RECT 10.185 24.840 550.570 70.360 ;
        RECT 10.185 23.440 550.170 24.840 ;
        RECT 10.185 8.335 550.570 23.440 ;
      LAYER met4 ;
        RECT 15.935 10.240 20.640 551.305 ;
        RECT 23.040 10.240 97.440 551.305 ;
        RECT 99.840 10.240 174.240 551.305 ;
        RECT 176.640 10.240 251.040 551.305 ;
        RECT 253.440 10.240 327.840 551.305 ;
        RECT 330.240 10.240 404.640 551.305 ;
        RECT 407.040 10.240 481.440 551.305 ;
        RECT 483.840 10.240 544.345 551.305 ;
        RECT 15.935 9.695 544.345 10.240 ;
  END
END bqmain
END LIBRARY

