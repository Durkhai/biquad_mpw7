* NGSPICE file created from bqmain.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt bqmain bq_clk_i nreset vccd1 vssd1 wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11]
+ wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18]
+ wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24]
+ wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30]
+ wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8]
+ wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12]
+ wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19]
+ wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25]
+ wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31]
+ wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9]
+ wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15]
+ wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21]
+ wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28]
+ wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5]
+ wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rst_i wb_stb_i wb_we_i x[0] x[10]
+ x[11] x[1] x[2] x[3] x[4] x[5] x[6] x[7] x[8] x[9] y[0] y[10] y[11] y[1] y[2] y[3]
+ y[4] y[5] y[6] y[7] y[8] y[9]
XANTENNA__11866__B1 _19363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18869_ _18670_/Y _18627_/Y _18465_/X vssd1 vssd1 vccd1 vccd1 _18869_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23119__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18794__A1 _12130_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16198__A _17631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20900_ _12674_/X _20471_/Y _20899_/Y vssd1 vssd1 vccd1 vccd1 _20900_/Y sky130_fd_sc_hd__o21ai_1
X_21880_ _21880_/A vssd1 vssd1 vccd1 vccd1 _22121_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11881__A3 _18952_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19338__A3 _19951_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20831_ _21121_/B _20887_/A _20887_/B vssd1 vssd1 vccd1 vccd1 _20841_/A sky130_fd_sc_hd__nand3_1
XANTENNA__21832__A _21832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19507__A1_N _19656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23550_ _23578_/CLK _23550_/D vssd1 vssd1 vccd1 vccd1 _23550_/Q sky130_fd_sc_hd__dfxtp_1
X_20762_ _20761_/B _20761_/C _23561_/Q vssd1 vssd1 vccd1 vccd1 _21030_/A sky130_fd_sc_hd__a21bo_1
XFILLER_39_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22501_ _22501_/A _22501_/B _22501_/C _22501_/D vssd1 vssd1 vccd1 vccd1 _22541_/D
+ sky130_fd_sc_hd__nand4_1
XANTENNA__16021__A2 _16073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23481_ _23518_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 _23481_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20693_ _20624_/X _20631_/X _20636_/X _20667_/B vssd1 vssd1 vccd1 vccd1 _20695_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16364__C _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13350__A _23472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22432_ _22434_/A _22434_/D vssd1 vssd1 vccd1 vccd1 _22457_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22363_ _22363_/A vssd1 vssd1 vccd1 vccd1 _22636_/C sky130_fd_sc_hd__buf_2
XANTENNA__19675__C _19675_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21314_ _21314_/A vssd1 vssd1 vccd1 vccd1 _21502_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22294_ _22476_/A _22476_/B _22569_/B vssd1 vssd1 vccd1 vccd1 _22362_/A sky130_fd_sc_hd__nand3_2
XFILLER_151_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21245_ _21414_/A _21415_/A _21240_/Y _21255_/A vssd1 vssd1 vccd1 vccd1 _21245_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14181__A _14181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21176_ _21369_/A _21370_/A _21176_/C _21182_/D vssd1 vssd1 vccd1 vccd1 _21179_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20127_ _20039_/B _20039_/A _20310_/C _20201_/C _20201_/A vssd1 vssd1 vccd1 vccd1
+ _20128_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_132_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15835__A2 _16027_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20058_ _20058_/A _20058_/B vssd1 vssd1 vccd1 vccd1 _20060_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13525__A _13547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11900_ _18849_/C vssd1 vssd1 vccd1 vccd1 _19548_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16539__C _16539_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16574__A_N _16294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12880_ _12606_/Y _12668_/X _12608_/X vssd1 vssd1 vccd1 vccd1 _12880_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_172_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _16027_/A vssd1 vssd1 vccd1 vccd1 _19180_/C sky130_fd_sc_hd__clkbuf_4
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18537__A1 _12378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18537__B2 _17591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18419__B1_N _23537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14550_ _14550_/A vssd1 vssd1 vccd1 vccd1 _14550_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16548__B1 _16549_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ _12183_/A vssd1 vssd1 vccd1 vccd1 _12343_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _22064_/C vssd1 vssd1 vccd1 vccd1 _22381_/C sky130_fd_sc_hd__buf_2
XFILLER_53_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _14492_/C _14380_/B _14410_/Y _14405_/Y vssd1 vssd1 vccd1 vccd1 _14486_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _23584_/Q vssd1 vssd1 vccd1 vccd1 _11720_/A sky130_fd_sc_hd__buf_2
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16220_ _16233_/B _16710_/A vssd1 vssd1 vccd1 vccd1 _16222_/A sky130_fd_sc_hd__nand2_1
XFILLER_186_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13432_ _13732_/A _13431_/X _13407_/Y _13410_/X _13433_/A vssd1 vssd1 vccd1 vccd1
+ _13432_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_155_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _17592_/A _17590_/A _16447_/A _15766_/X _18756_/A vssd1 vssd1 vccd1 vccd1
+ _16152_/A sky130_fd_sc_hd__o221ai_4
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ _13620_/C _13351_/X _13357_/Y _13362_/Y vssd1 vssd1 vccd1 vccd1 _13364_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_158_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23524__CLK _23538_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15102_ _15102_/A _15102_/B vssd1 vssd1 vccd1 vccd1 _15446_/B sky130_fd_sc_hd__nand2_2
XFILLER_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20805__B _21065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12314_ _12508_/A _16529_/C _16500_/D _12327_/A vssd1 vssd1 vccd1 vccd1 _12314_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16082_ _16022_/A _15895_/C _16021_/Y vssd1 vssd1 vccd1 vccd1 _16084_/B sky130_fd_sc_hd__a21o_1
X_13294_ _22361_/C vssd1 vssd1 vccd1 vccd1 _21891_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19910_ _19928_/C _19928_/D vssd1 vssd1 vccd1 vccd1 _19911_/A sky130_fd_sc_hd__nand2_1
X_15033_ _15036_/A _15033_/B _15033_/C vssd1 vssd1 vccd1 vccd1 _15050_/A sky130_fd_sc_hd__nand3b_2
XFILLER_181_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12245_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12245_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__19265__A2 _20366_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19841_ _19848_/A _19868_/A _19949_/D vssd1 vssd1 vccd1 vccd1 _19841_/Y sky130_fd_sc_hd__nand3_1
X_12176_ _12173_/X _12174_/X _18600_/C _12175_/X vssd1 vssd1 vccd1 vccd1 _12177_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19772_ _19772_/A vssd1 vssd1 vccd1 vccd1 _19772_/Y sky130_fd_sc_hd__inv_2
X_16984_ _17010_/C _16761_/Y _16983_/Y vssd1 vssd1 vccd1 vccd1 _16984_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18723_ _12473_/C _12473_/A _12473_/B _12480_/B vssd1 vssd1 vccd1 vccd1 _18723_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_7_1154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output56_A _14619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15935_ _15640_/Y _15917_/Y _17885_/A _16372_/A _15925_/Y vssd1 vssd1 vccd1 vccd1
+ _16281_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17579__A2 _17565_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18654_ _18973_/B vssd1 vssd1 vccd1 vccd1 _18972_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _15985_/C _15866_/B vssd1 vssd1 vccd1 vccd1 _15867_/C sky130_fd_sc_hd__nor2_1
XANTENNA__15353__C _15353_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17605_ _17605_/A _17605_/B _20055_/C _20055_/D vssd1 vssd1 vccd1 vccd1 _17605_/Y
+ sky130_fd_sc_hd__nand4_4
X_14817_ _14835_/C _23505_/Q vssd1 vssd1 vccd1 vccd1 _14855_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18585_ _18568_/A _18584_/Y _18576_/A vssd1 vssd1 vccd1 vccd1 _18586_/C sky130_fd_sc_hd__o21ai_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15797_ _15797_/A vssd1 vssd1 vccd1 vccd1 _17465_/A sky130_fd_sc_hd__buf_4
XANTENNA__16746__A _17898_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17536_ _17536_/A vssd1 vssd1 vccd1 vccd1 _18208_/A sky130_fd_sc_hd__buf_2
XANTENNA__15650__A _17098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14748_ _14961_/A vssd1 vssd1 vccd1 vccd1 _15439_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22186__C _22186_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17467_ _17597_/A vssd1 vssd1 vccd1 vccd1 _17467_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14679_ _23338_/Q _14668_/X _14673_/X _23306_/Q _14678_/X vssd1 vssd1 vccd1 vccd1
+ _14679_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15800__D _19308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19206_ _19013_/X _19192_/Y _19197_/Y _19201_/Y _19205_/X vssd1 vssd1 vccd1 vccd1
+ _19206_/X sky130_fd_sc_hd__a41o_1
X_16418_ _16418_/A vssd1 vssd1 vccd1 vccd1 _16474_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17398_ _17395_/Y _17806_/A _17397_/Y _17239_/X vssd1 vssd1 vccd1 vccd1 _17493_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_192_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19137_ _19354_/A _19354_/B _19391_/A vssd1 vssd1 vccd1 vccd1 _19140_/B sky130_fd_sc_hd__nand3_1
XFILLER_118_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_439 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16349_ _16581_/A _16581_/B _16276_/A vssd1 vssd1 vccd1 vccd1 _16771_/B sky130_fd_sc_hd__a21o_1
XFILLER_157_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19068_ _18889_/Y _18867_/Y _18885_/Y vssd1 vssd1 vccd1 vccd1 _19069_/C sky130_fd_sc_hd__a21oi_4
XFILLER_145_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18019_ _18022_/A _18022_/B _18015_/X _18018_/X vssd1 vssd1 vccd1 vccd1 _18028_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_172_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19792__A _19792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21030_ _21030_/A _21030_/B _21030_/C vssd1 vssd1 vccd1 vccd1 _21031_/C sky130_fd_sc_hd__nand3_1
XANTENNA__21063__A2 _21061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19661__C1 _19659_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23464__D _23476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11839__B1 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19016__B _19148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22981_ _23038_/S vssd1 vssd1 vccd1 vccd1 _22990_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_41_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22563__A2 _22059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21932_ _21783_/X _21755_/X _21760_/X vssd1 vssd1 vccd1 vccd1 _21936_/B sky130_fd_sc_hd__a21bo_4
XFILLER_94_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21863_ _22107_/D _22455_/A _21859_/A _21859_/B vssd1 vssd1 vccd1 vccd1 _21864_/C
+ sky130_fd_sc_hd__o211ai_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20814_ _20814_/A vssd1 vssd1 vccd1 vccd1 _21278_/A sky130_fd_sc_hd__clkbuf_2
X_21794_ _13561_/A _22564_/C _21792_/Y _21793_/Y vssd1 vssd1 vccd1 vccd1 _21794_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_179_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19192__A1 _16437_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19192__B2 _19649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23533_ _23558_/CLK _23533_/D vssd1 vssd1 vccd1 vccd1 _23533_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20745_ _20868_/A _20738_/A _20747_/C vssd1 vssd1 vccd1 vccd1 _20748_/A sky130_fd_sc_hd__a21o_1
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22079__A1 _21936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23464_ _23559_/CLK _23476_/Q vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
X_20676_ _20676_/A _20676_/B vssd1 vssd1 vccd1 vccd1 _20676_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22415_ _22288_/B _22288_/A _22289_/B vssd1 vssd1 vccd1 vccd1 _22415_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_164_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23395_ _23395_/CLK _23395_/D vssd1 vssd1 vccd1 vccd1 _23395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_878 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22346_ _22346_/A _22346_/B _22445_/C _22445_/D vssd1 vssd1 vccd1 vccd1 _22351_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_128_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22277_ _22364_/B vssd1 vssd1 vccd1 vccd1 _22479_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12030_ _12130_/A vssd1 vssd1 vccd1 vccd1 _12051_/A sky130_fd_sc_hd__buf_4
X_21228_ _21228_/A _21228_/B _21228_/C _21228_/D vssd1 vssd1 vccd1 vccd1 _21333_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_105_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21159_ _21159_/A _21159_/B vssd1 vssd1 vccd1 vccd1 _21228_/B sky130_fd_sc_hd__nand2_1
XANTENNA__22003__A1 _13642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23200__A0 _15664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16481__A2 _16451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13981_ _13972_/X _14795_/C _13985_/D _14246_/A _14791_/B vssd1 vssd1 vccd1 vccd1
+ _14150_/D sky130_fd_sc_hd__a32o_1
XFILLER_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18758__A1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13255__A _13660_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15720_ _15798_/A _15799_/A vssd1 vssd1 vccd1 vccd1 _16200_/A sky130_fd_sc_hd__nand2_1
XFILLER_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12932_ _12932_/A vssd1 vssd1 vccd1 vccd1 _13177_/A sky130_fd_sc_hd__buf_2
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15651_ _16921_/C _16113_/A _15641_/Y _15650_/Y vssd1 vssd1 vccd1 vccd1 _15651_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _12709_/A _12862_/X _12858_/A vssd1 vssd1 vccd1 vccd1 _12867_/B sky130_fd_sc_hd__o21ai_4
XFILLER_73_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17981__A2 _20210_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _13603_/X _14550_/X _14526_/X _12875_/B _14601_/X vssd1 vssd1 vccd1 vccd1
+ _14602_/X sky130_fd_sc_hd__a221o_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _18405_/A _18370_/B _18370_/C vssd1 vssd1 vccd1 vccd1 _18371_/B sky130_fd_sc_hd__nor3_1
X_11814_ _11814_/A vssd1 vssd1 vccd1 vccd1 _12238_/A sky130_fd_sc_hd__buf_2
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _23512_/Q _15582_/B vssd1 vssd1 vccd1 vccd1 _23500_/D sky130_fd_sc_hd__xnor2_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12794_/A _12794_/B vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17326_/B _17326_/C _17134_/A vssd1 vssd1 vccd1 vccd1 _17322_/C sky130_fd_sc_hd__a21bo_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14533_ _14535_/A _14538_/A _14538_/B _14538_/C vssd1 vssd1 vccd1 vccd1 _23184_/D
+ sky130_fd_sc_hd__nor4_2
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19877__A _20003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11745_/A _12100_/C vssd1 vssd1 vccd1 vccd1 _11746_/C sky130_fd_sc_hd__nand2_1
XFILLER_187_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17252_/A _17433_/A vssd1 vssd1 vccd1 vccd1 _17252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14464_ _14465_/A _14465_/B _14465_/C _14465_/D vssd1 vssd1 vccd1 vccd1 _14464_/Y
+ sky130_fd_sc_hd__a22oi_1
X_11676_ _11980_/A vssd1 vssd1 vccd1 vccd1 _11676_/X sky130_fd_sc_hd__buf_2
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _15761_/X _15920_/B _15631_/B _15637_/D _15932_/A vssd1 vssd1 vccd1 vccd1
+ _16203_/Y sky130_fd_sc_hd__a41oi_4
X_13415_ _13486_/A vssd1 vssd1 vccd1 vccd1 _13415_/X sky130_fd_sc_hd__buf_2
XFILLER_179_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17183_ _16954_/Y _17173_/B _16944_/X vssd1 vssd1 vccd1 vccd1 _17183_/Y sky130_fd_sc_hd__o21ai_1
X_14395_ _14395_/A _14395_/B vssd1 vssd1 vccd1 vccd1 _14396_/C sky130_fd_sc_hd__nand2_1
XANTENNA__17828__C _23528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_856 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_630 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16134_ _12208_/A _16377_/A _15975_/B _16128_/X _16610_/A vssd1 vssd1 vccd1 vccd1
+ _16135_/C sky130_fd_sc_hd__o221ai_2
XFILLER_155_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21293__A2 _20471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13346_ _23325_/Q vssd1 vssd1 vccd1 vccd1 _13394_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16065_ _19196_/A vssd1 vssd1 vccd1 vccd1 _19670_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_185_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13277_ _13642_/A vssd1 vssd1 vccd1 vccd1 _13469_/A sky130_fd_sc_hd__buf_2
XFILLER_142_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15016_ _14058_/X _15366_/A _14903_/B _14872_/Y vssd1 vssd1 vccd1 vccd1 _15022_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_12228_ _12203_/Y _12220_/Y _12540_/B _12532_/B vssd1 vssd1 vccd1 vccd1 _12542_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_64_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12191__C1 _12308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22793__A2 _22560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19824_ _19802_/A _19802_/B _19823_/Y vssd1 vssd1 vccd1 vccd1 _19836_/A sky130_fd_sc_hd__o21ai_1
XFILLER_123_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12159_ _12159_/A _12159_/B _12159_/C vssd1 vssd1 vccd1 vccd1 _12159_/X sky130_fd_sc_hd__and3_1
XFILLER_116_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19755_ _19755_/A _19755_/B vssd1 vssd1 vccd1 vccd1 _19755_/Y sky130_fd_sc_hd__nand2_1
X_16967_ _18161_/C vssd1 vssd1 vccd1 vccd1 _18277_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_111_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15680__B1 _14569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19946__B1 _23396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17860__A _17860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18706_ _18706_/A _18706_/B vssd1 vssd1 vccd1 vccd1 _18708_/A sky130_fd_sc_hd__nand2_1
X_15918_ _15921_/C _15918_/B _15918_/C vssd1 vssd1 vccd1 vccd1 _15937_/A sky130_fd_sc_hd__nand3b_4
XANTENNA__18213__A3 _17324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19686_ _19686_/A _19688_/A _19688_/B vssd1 vssd1 vccd1 vccd1 _19740_/A sky130_fd_sc_hd__nand3_2
XFILLER_64_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16898_ _16904_/A _16908_/A _16913_/B vssd1 vssd1 vccd1 vccd1 _16898_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17421__A1 _12237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_707 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_567 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15849_ _15753_/B _15975_/A _15844_/A vssd1 vssd1 vccd1 vccd1 _15858_/A sky130_fd_sc_hd__o21ai_1
XFILLER_52_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18637_ _18443_/A _18453_/A _18804_/A vssd1 vssd1 vccd1 vccd1 _18639_/A sky130_fd_sc_hd__o21ai_2
XFILLER_91_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18394__C _18417_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18568_ _18568_/A _18568_/B _18568_/C vssd1 vssd1 vccd1 vccd1 _18569_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19174__A1 _16437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12797__A1 _20957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19174__B2 _12323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17519_ _17699_/A _17519_/B vssd1 vssd1 vccd1 vccd1 _17523_/B sky130_fd_sc_hd__nand2_1
X_18499_ _18499_/A _18499_/B _18499_/C vssd1 vssd1 vccd1 vccd1 _18529_/A sky130_fd_sc_hd__nand3_1
XFILLER_71_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12509__A _12509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20530_ _13056_/X _12766_/X _13053_/X _20676_/A _20670_/A vssd1 vssd1 vccd1 vccd1
+ _20530_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20461_ _20902_/B _23458_/Q vssd1 vssd1 vccd1 vccd1 _20612_/A sky130_fd_sc_hd__nor2_1
XANTENNA__14724__A _23597_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19331__D1 _19543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22200_ _22200_/A _22200_/B _22200_/C vssd1 vssd1 vccd1 vccd1 _22200_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__23459__D _23471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23180_ _23412_/Q input30/X _23182_/S vssd1 vssd1 vccd1 vccd1 _23181_/A sky130_fd_sc_hd__mux2_1
X_20392_ _20392_/A _20392_/B vssd1 vssd1 vccd1 vccd1 _20393_/B sky130_fd_sc_hd__nand2_1
XFILLER_134_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13985__D _13985_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20164__C _20164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22131_ _21922_/B _22012_/Y _22062_/X vssd1 vssd1 vccd1 vccd1 _22136_/B sky130_fd_sc_hd__a21o_1
XFILLER_145_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22062_ _13803_/A _13803_/B _13469_/A vssd1 vssd1 vccd1 vccd1 _22062_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20461__A _20902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21013_ _20999_/X _21003_/X _21006_/Y _21012_/X vssd1 vssd1 vccd1 vccd1 _21243_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_59_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22964_ _23316_/Q input30/X _22966_/S vssd1 vssd1 vccd1 vccd1 _22965_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15018__A3 _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21915_ _22045_/A _22045_/B _22269_/C _22043_/A _22364_/B vssd1 vssd1 vccd1 vccd1
+ _21918_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_167_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22895_ _22895_/A _22895_/B vssd1 vssd1 vccd1 vccd1 _23578_/D sky130_fd_sc_hd__nor2_1
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21846_ _21836_/Y _21837_/Y _21834_/Y _21826_/X vssd1 vssd1 vccd1 vccd1 _21847_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_71_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16536__D _17326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21777_ _21777_/A _21777_/B vssd1 vssd1 vccd1 vccd1 _22364_/B sky130_fd_sc_hd__nand2_4
XFILLER_90_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23516_ _23518_/CLK input52/X vssd1 vssd1 vccd1 vccd1 _23516_/Q sky130_fd_sc_hd__dfxtp_1
X_20728_ _20728_/A vssd1 vssd1 vccd1 vccd1 _20728_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23447_ _23559_/CLK hold25/X vssd1 vssd1 vccd1 vccd1 _23447_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_165_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14634__A _14688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20659_ _20479_/X _20639_/Y _20894_/A _20641_/A vssd1 vssd1 vccd1 vccd1 _20662_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11748__C1 _11743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13200_ _13147_/A _13147_/B _13147_/C vssd1 vssd1 vccd1 vccd1 _13201_/C sky130_fd_sc_hd__a21o_1
XFILLER_183_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14180_ _14180_/A _14180_/B _14180_/C vssd1 vssd1 vccd1 vccd1 _14220_/A sky130_fd_sc_hd__nand3_4
XFILLER_178_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23378_ _23378_/CLK _23378_/D vssd1 vssd1 vccd1 vccd1 _23378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _13131_/A vssd1 vssd1 vccd1 vccd1 _21435_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22329_ _22332_/A _22332_/B _22332_/C vssd1 vssd1 vccd1 vccd1 _22333_/A sky130_fd_sc_hd__a21o_1
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16151__B2 _15766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22224__A1 _21988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13062_ _13055_/X _13060_/X _13061_/Y vssd1 vssd1 vccd1 vccd1 _13062_/X sky130_fd_sc_hd__o21a_1
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12013_ _18859_/B _18859_/C _12306_/A _12262_/B vssd1 vssd1 vccd1 vccd1 _12013_/Y
+ sky130_fd_sc_hd__nand4_2
X_17870_ _17988_/A _17982_/A _17982_/B vssd1 vssd1 vccd1 vccd1 _17874_/A sky130_fd_sc_hd__a21oi_1
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16821_ _16821_/A _17449_/A _17040_/A _17041_/C vssd1 vssd1 vccd1 vccd1 _16821_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_120_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12601__B _12601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_bq_clk_i clkbuf_4_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _23571_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_87_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19540_ _19540_/A _19540_/B vssd1 vssd1 vccd1 vccd1 _19542_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16752_ _16266_/A _16266_/B _16266_/C _16281_/D _16275_/A vssd1 vssd1 vccd1 vccd1
+ _16752_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_150_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13964_ _14331_/C _14331_/A vssd1 vssd1 vccd1 vccd1 _13964_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20538__A1 _20957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15703_ _23419_/Q _15727_/B _15656_/X vssd1 vssd1 vccd1 vccd1 _15815_/A sky130_fd_sc_hd__o21a_2
X_12915_ _12915_/A vssd1 vssd1 vccd1 vccd1 _13158_/A sky130_fd_sc_hd__clkbuf_2
X_19471_ _19471_/A _19471_/B vssd1 vssd1 vccd1 vccd1 _19471_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16683_ _16683_/A vssd1 vssd1 vccd1 vccd1 _16683_/X sky130_fd_sc_hd__buf_4
XFILLER_80_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13895_ _23504_/Q vssd1 vssd1 vccd1 vccd1 _14936_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18422_ _18407_/C _18408_/B _18430_/A _18420_/X vssd1 vssd1 vccd1 vccd1 _18423_/B
+ sky130_fd_sc_hd__a211oi_1
X_15634_ _15634_/A _15634_/B _15634_/C vssd1 vssd1 vccd1 vccd1 _15927_/A sky130_fd_sc_hd__nand3_1
XFILLER_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15965__A1 _16523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12846_ _12846_/A _12901_/B vssd1 vssd1 vccd1 vccd1 _12896_/A sky130_fd_sc_hd__nand2_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _18296_/X _18295_/X _18267_/Y vssd1 vssd1 vccd1 vccd1 _18353_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15565_ _15468_/X _15538_/A _15538_/D _15564_/Y _15559_/A vssd1 vssd1 vccd1 vccd1
+ _15566_/S sky130_fd_sc_hd__a311o_4
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12777_/A _12901_/A _12845_/A vssd1 vssd1 vccd1 vccd1 _12779_/B sky130_fd_sc_hd__nand3_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17506_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14633_/A _14519_/D _14633_/B _14633_/C vssd1 vssd1 vccd1 vccd1 _14516_/X
+ sky130_fd_sc_hd__or4_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18284_ _18284_/A _18284_/B vssd1 vssd1 vccd1 vccd1 _18285_/B sky130_fd_sc_hd__nor2_1
X_11728_ _16661_/C vssd1 vssd1 vccd1 vccd1 _19161_/A sky130_fd_sc_hd__buf_2
X_15496_ _15496_/A vssd1 vssd1 vccd1 vccd1 _15516_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17235_ _17235_/A vssd1 vssd1 vccd1 vccd1 _19949_/D sky130_fd_sc_hd__buf_2
XFILLER_119_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447_ _14806_/A vssd1 vssd1 vccd1 vccd1 _15208_/A sky130_fd_sc_hd__clkbuf_2
X_11659_ _23387_/Q _23386_/Q vssd1 vssd1 vccd1 vccd1 _11983_/A sky130_fd_sc_hd__nor2_2
XFILLER_174_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14544__A _14693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_962 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17166_ _17166_/A _17166_/B _17350_/A _17170_/B vssd1 vssd1 vccd1 vccd1 _17167_/D
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18667__B1 _18665_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14378_ _15017_/D vssd1 vssd1 vccd1 vccd1 _15358_/A sky130_fd_sc_hd__buf_2
XFILLER_128_675 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16117_ _17326_/D _17035_/C _18172_/A _18219_/D _15926_/X vssd1 vssd1 vccd1 vccd1
+ _16275_/A sky130_fd_sc_hd__a41o_2
XFILLER_31_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12951__A1 _12640_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16257__A2_N _16254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13329_ _13660_/C vssd1 vssd1 vccd1 vccd1 _13701_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17097_ _16856_/Y _17093_/Y _15991_/A _17096_/X _15807_/A vssd1 vssd1 vccd1 vccd1
+ _17097_/Y sky130_fd_sc_hd__o2111ai_2
XFILLER_6_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17890__A1 _17643_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16048_ _11792_/A _11792_/B _15821_/A _16451_/C vssd1 vssd1 vccd1 vccd1 _16490_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19807_ _19807_/A vssd1 vssd1 vccd1 vccd1 _19807_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17999_ _17999_/A _17999_/B _18085_/B _17999_/D vssd1 vssd1 vccd1 vccd1 _18022_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22518__A2 _22521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15653__B1 _16661_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19738_ _19719_/Y _19893_/A _19726_/X vssd1 vssd1 vccd1 vccd1 _19880_/B sky130_fd_sc_hd__a21o_1
XFILLER_42_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19669_ _19670_/A _18455_/A _18461_/C _20209_/A _16066_/C vssd1 vssd1 vccd1 vccd1
+ _19669_/X sky130_fd_sc_hd__o32a_1
X_21700_ _21717_/B _21717_/A vssd1 vssd1 vccd1 vccd1 _21700_/Y sky130_fd_sc_hd__nand2_1
X_22680_ _22677_/Y _22549_/B _22675_/Y _22676_/Y vssd1 vssd1 vccd1 vccd1 _22680_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21631_ _21631_/A _21631_/B _21631_/C vssd1 vssd1 vccd1 vccd1 _21631_/Y sky130_fd_sc_hd__nand3_1
X_21562_ _21428_/X _21552_/A _21561_/Y _21559_/B vssd1 vssd1 vccd1 vccd1 _21564_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23301_ _23397_/CLK _23301_/D vssd1 vssd1 vccd1 vccd1 _23301_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20513_ _20556_/A _20556_/B _13032_/X vssd1 vssd1 vccd1 vccd1 _20515_/B sky130_fd_sc_hd__a21o_1
XFILLER_166_759 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21493_ _21493_/A _21493_/B _21493_/C vssd1 vssd1 vccd1 vccd1 _21495_/B sky130_fd_sc_hd__and3_1
XFILLER_176_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20444_ _20444_/A _20444_/B vssd1 vssd1 vccd1 vccd1 _23537_/D sky130_fd_sc_hd__nor2_1
X_23232_ _23232_/A vssd1 vssd1 vccd1 vccd1 _23434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20375_ _20428_/B _20428_/C vssd1 vssd1 vccd1 vccd1 _20401_/B sky130_fd_sc_hd__xor2_1
X_23163_ _23404_/Q input21/X _23167_/S vssd1 vssd1 vccd1 vccd1 _23164_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22114_ _21979_/B _21977_/B _21975_/Y vssd1 vssd1 vccd1 vccd1 _22115_/B sky130_fd_sc_hd__a21oi_2
XFILLER_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23094_ _23094_/A vssd1 vssd1 vccd1 vccd1 _23373_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__22047__A_N _14614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22045_ _22045_/A _22045_/B vssd1 vssd1 vccd1 vccd1 _22045_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__19083__B1 _19082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12702__A _23447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16436__A2 _11883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17094__C1 _16591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_798 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22947_ _23308_/Q input21/X _22951_/S vssd1 vssd1 vccd1 vccd1 _22948_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17936__A2 _18208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_846 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12700_ _20670_/C _21271_/B _20663_/D _21054_/C vssd1 vssd1 vccd1 vccd1 _12700_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13407__C1 _22145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ _13680_/A _13680_/B _13680_/C _13680_/D vssd1 vssd1 vccd1 vccd1 _13680_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_141_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22878_ _22878_/A _22878_/B _22887_/C vssd1 vssd1 vccd1 vccd1 _22881_/B sky130_fd_sc_hd__nand3_1
XFILLER_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12631_ _23448_/Q vssd1 vssd1 vccd1 vccd1 _12632_/A sky130_fd_sc_hd__inv_2
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21829_ _21829_/A vssd1 vssd1 vccd1 vccd1 _22754_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15350_ _15350_/A _15353_/C _15350_/C vssd1 vssd1 vccd1 vccd1 _15350_/X sky130_fd_sc_hd__and3_1
XFILLER_34_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12562_ _12396_/A _12396_/B _12396_/C vssd1 vssd1 vccd1 vccd1 _12563_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__16357__D1 _16046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14301_ _14307_/A _14310_/C vssd1 vssd1 vccd1 vccd1 _14303_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15281_ _15292_/B _15292_/A vssd1 vssd1 vccd1 vccd1 _15392_/B sky130_fd_sc_hd__and2_1
XFILLER_184_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12493_ _12492_/Y _12161_/Y _12158_/A _12198_/B vssd1 vssd1 vccd1 vccd1 _12494_/C
+ sky130_fd_sc_hd__a22oi_1
X_17020_ _17381_/A _17019_/A _17019_/B _17019_/C vssd1 vssd1 vccd1 vccd1 _17020_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14232_ _14215_/Y _14218_/Y _14816_/A _14228_/B vssd1 vssd1 vccd1 vccd1 _14826_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_184_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23265__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19310__A1 _19304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12933__A1 _12571_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16124__A1 _11971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ _15253_/C _14163_/B _15253_/A _14252_/D vssd1 vssd1 vccd1 vccd1 _14164_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__21909__B _22064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_0_0_bq_clk_i_A clkbuf_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13114_ _21050_/C _13119_/A _13119_/B _13116_/C _21050_/D vssd1 vssd1 vccd1 vccd1
+ _13114_/X sky130_fd_sc_hd__a32o_1
XFILLER_124_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14094_ _14094_/A vssd1 vssd1 vccd1 vccd1 _14094_/X sky130_fd_sc_hd__clkbuf_2
X_18971_ _18971_/A vssd1 vssd1 vccd1 vccd1 _18971_/X sky130_fd_sc_hd__buf_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15195__A _15195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20532__C _23455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17922_ _17922_/A vssd1 vssd1 vccd1 vccd1 _17922_/X sky130_fd_sc_hd__buf_2
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13708__A _22145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13045_ _12867_/A _12867_/B _12867_/C _13044_/Y _12900_/A vssd1 vssd1 vccd1 vccd1
+ _13048_/B sky130_fd_sc_hd__a32oi_4
XFILLER_79_732 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17853_ _17853_/A vssd1 vssd1 vccd1 vccd1 _17982_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16804_ _16804_/A _16804_/B vssd1 vssd1 vccd1 vccd1 _17040_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17784_ _17768_/Y _17773_/Y _17771_/Y vssd1 vssd1 vccd1 vccd1 _17784_/Y sky130_fd_sc_hd__a21oi_1
X_14996_ _14887_/B _15099_/A _14992_/Y _15104_/A _14469_/C vssd1 vssd1 vccd1 vccd1
+ _15004_/C sky130_fd_sc_hd__o2111ai_2
XANTENNA__23562__D _23562_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19523_ _19523_/A _19577_/C vssd1 vssd1 vccd1 vccd1 _19526_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13947_ _13977_/B _14001_/A _13945_/X _14094_/A _13908_/C vssd1 vssd1 vccd1 vccd1
+ _13951_/A sky130_fd_sc_hd__o311ai_2
X_16735_ _16735_/A _16735_/B _16735_/C vssd1 vssd1 vccd1 vccd1 _16739_/B sky130_fd_sc_hd__nand3_1
XFILLER_75_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16457__C _17845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19454_ _19449_/Y _19450_/X _19461_/A vssd1 vssd1 vccd1 vccd1 _19456_/A sky130_fd_sc_hd__o21a_1
X_16666_ _16781_/B _16665_/X _14631_/X vssd1 vssd1 vccd1 vccd1 _16669_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__15938__A1 _16921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ _14863_/C vssd1 vssd1 vccd1 vccd1 _14001_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18405_ _18405_/A vssd1 vssd1 vccd1 vccd1 _18407_/A sky130_fd_sc_hd__inv_2
XFILLER_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15617_ _15622_/A _15712_/C _15631_/B _15624_/A vssd1 vssd1 vccd1 vccd1 _15618_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12829_ _20961_/A _12796_/A _12828_/Y vssd1 vssd1 vccd1 vccd1 _12835_/C sky130_fd_sc_hd__o21ai_2
X_19385_ _19385_/A _19385_/B _19385_/C vssd1 vssd1 vccd1 vccd1 _19468_/A sky130_fd_sc_hd__nand3_2
X_16597_ _16597_/A _16597_/B _16597_/C vssd1 vssd1 vccd1 vccd1 _16647_/A sky130_fd_sc_hd__nand3_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18336_ _18335_/B _17323_/X _17324_/X _18378_/C _18335_/D vssd1 vssd1 vccd1 vccd1
+ _18337_/B sky130_fd_sc_hd__a32o_1
X_15548_ _15548_/A vssd1 vssd1 vccd1 vccd1 _15548_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11975__A2 _11902_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11898__A _18461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_562 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18267_ _18267_/A vssd1 vssd1 vccd1 vccd1 _18267_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15479_ _15479_/A _15479_/B vssd1 vssd1 vccd1 vccd1 _23280_/D sky130_fd_sc_hd__nand2_1
XFILLER_175_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ _17218_/A vssd1 vssd1 vccd1 vccd1 _17536_/A sky130_fd_sc_hd__clkbuf_2
X_18198_ _18252_/A _18252_/B _18198_/C vssd1 vssd1 vccd1 vccd1 _18302_/C sky130_fd_sc_hd__nor3_2
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12506__B _12506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17149_ _17149_/A _17631_/A _17712_/D vssd1 vssd1 vccd1 vccd1 _17150_/B sky130_fd_sc_hd__and3_1
XFILLER_190_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17312__B1 _16908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14126__B1 _14070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20160_ _20160_/A _20160_/B vssd1 vssd1 vccd1 vccd1 _20167_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16666__A2 _16665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20091_ _19996_/A _19996_/B _19996_/C _19963_/B vssd1 vssd1 vccd1 vccd1 _20091_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_97_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12152__A2 _12324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_884 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15626__B1 _15664_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22801_ _22756_/D _22756_/B _22861_/C _22800_/X vssd1 vssd1 vccd1 vccd1 _22801_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19024__B _19029_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20993_ _20846_/A _20847_/A _20847_/B vssd1 vssd1 vccd1 vccd1 _20995_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__14449__A _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13353__A _23325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22732_ _22537_/X _22729_/C _22697_/X vssd1 vssd1 vccd1 vccd1 _22732_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15929__A1 _16281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16051__B1 _17226_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22663_ _22716_/A _22663_/B _22663_/C _22663_/D vssd1 vssd1 vccd1 vccd1 _22725_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__14062__C1 _14760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14601__A1 _23580_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14601__B2 _14188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21614_ _21529_/X _21614_/B _21614_/C _21614_/D vssd1 vssd1 vccd1 vccd1 _21614_/Y
+ sky130_fd_sc_hd__nand4b_2
XANTENNA__19040__A _19040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22594_ _22594_/A _22594_/B _22594_/C vssd1 vssd1 vccd1 vccd1 _22605_/A sky130_fd_sc_hd__nand3_1
XFILLER_187_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21545_ _21545_/A _21635_/A _21592_/A _21635_/B vssd1 vssd1 vccd1 vccd1 _21545_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14184__A _14184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11601__A _23397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13707__A3 _21987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19694__B _19799_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21476_ _21476_/A _21476_/B vssd1 vssd1 vccd1 vccd1 _21477_/B sky130_fd_sc_hd__xor2_1
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11718__A2 _11670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23215_ _14631_/X input11/X _23217_/S vssd1 vssd1 vccd1 vccd1 _23216_/A sky130_fd_sc_hd__mux2_1
X_20427_ _20314_/X _20368_/C _20269_/B _20371_/B vssd1 vssd1 vccd1 vccd1 _20427_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17321__B1_N _17134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23146_ _23146_/A vssd1 vssd1 vccd1 vccd1 _23396_/D sky130_fd_sc_hd__clkbuf_1
X_20358_ _20359_/B _20355_/Y _20356_/Y _20357_/Y vssd1 vssd1 vccd1 vccd1 _20358_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_122_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15865__B1 _12518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20289_ _20284_/X _20287_/X _20288_/X vssd1 vssd1 vccd1 vccd1 _20295_/B sky130_fd_sc_hd__a21bo_2
XFILLER_121_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23077_ _23077_/A vssd1 vssd1 vccd1 vccd1 _23365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15446__C _15446_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12143__A2 _12110_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17606__A1 _14599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22028_ _22028_/A _22028_/B vssd1 vssd1 vccd1 vccd1 _22028_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13247__B _22365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17942__B _23529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17082__A2 _16451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14850_ _23270_/D _14749_/X _14849_/Y vssd1 vssd1 vccd1 vccd1 _14850_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19359__A1 _18673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13801_ _13394_/A _21744_/C _13355_/A _13783_/B vssd1 vssd1 vccd1 vccd1 _13803_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA_input18_A wb_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14781_ _14781_/A _14781_/B vssd1 vssd1 vccd1 vccd1 _14788_/C sky130_fd_sc_hd__nand2_1
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11993_ _11757_/A _18812_/B _11608_/A vssd1 vssd1 vccd1 vccd1 _12121_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__13643__A2 _13642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ _16522_/A _16522_/B _16519_/Y vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__a21oi_1
XFILLER_95_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13263__A _23322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13732_ _13732_/A _13732_/B _13732_/C vssd1 vssd1 vccd1 vccd1 _13732_/X sky130_fd_sc_hd__or3_1
XFILLER_56_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16451_ _16458_/A _16451_/B _16451_/C vssd1 vssd1 vccd1 vccd1 _16451_/X sky130_fd_sc_hd__or3_1
XFILLER_32_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13663_ _13663_/A _22562_/B _13663_/C _21882_/B vssd1 vssd1 vccd1 vccd1 _13663_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17790__B1 _17792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15402_ _15402_/A _15402_/B _15442_/D _15442_/C vssd1 vssd1 vccd1 vccd1 _15439_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ _18984_/B _19309_/A _19158_/Y _19162_/B vssd1 vssd1 vccd1 vccd1 _19172_/B
+ sky130_fd_sc_hd__o211ai_4
X_12614_ _23448_/Q vssd1 vssd1 vccd1 vccd1 _20784_/C sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _16382_/A vssd1 vssd1 vccd1 vccd1 _17285_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13594_ _13698_/A _13698_/B _13593_/X vssd1 vssd1 vccd1 vccd1 _13594_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18334__A2 _17723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18121_ _18123_/A _18123_/B _18123_/C _18133_/B vssd1 vssd1 vccd1 vccd1 _18134_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_169_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19531__A1 _18859_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19531__B2 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15333_ _15279_/B _15292_/X _15332_/X vssd1 vssd1 vccd1 vccd1 _15395_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20527__C _23454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12545_ _18571_/A _18571_/B _12557_/A vssd1 vssd1 vccd1 vccd1 _12545_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_184_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18052_ _17922_/X _17924_/X _17930_/Y _17957_/Y _18049_/B vssd1 vssd1 vccd1 vccd1
+ _18138_/A sky130_fd_sc_hd__o221ai_2
X_15264_ _15350_/C _15409_/A _15419_/A _15260_/X _15259_/Y vssd1 vssd1 vccd1 vccd1
+ _15264_/Y sky130_fd_sc_hd__a32oi_1
X_12476_ _18945_/C _19485_/A _12177_/Y _12475_/X vssd1 vssd1 vccd1 vccd1 _12478_/C
+ sky130_fd_sc_hd__a31o_2
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17003_ _17003_/A _17003_/B vssd1 vssd1 vccd1 vccd1 _17003_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18098__A1 _16478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14215_ _14220_/A _14220_/B _14221_/B vssd1 vssd1 vccd1 vccd1 _14215_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_172_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23091__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15195_ _15195_/A _15195_/B _15195_/C vssd1 vssd1 vccd1 vccd1 _15201_/A sky130_fd_sc_hd__and3_1
XFILLER_125_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output86_A _23262_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _14222_/A _14222_/B _14217_/C _14218_/A vssd1 vssd1 vccd1 vccd1 _14148_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21358__C _21358_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14659__A1 _15338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18954_ _18938_/X _18952_/Y _18953_/X vssd1 vssd1 vccd1 vccd1 _18954_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14077_ _14124_/A _23357_/Q _14077_/C vssd1 vssd1 vccd1 vccd1 _14864_/B sky130_fd_sc_hd__nor3_2
XANTENNA__12342__A _19512_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12134__A2 _11849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17905_ _17905_/A _17905_/B _17905_/C vssd1 vssd1 vccd1 vccd1 _17916_/C sky130_fd_sc_hd__nand3_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13028_ _20556_/A _20556_/B vssd1 vssd1 vccd1 vccd1 _13028_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18885_ _18868_/X _18870_/Y _18864_/Y _18866_/Y vssd1 vssd1 vccd1 vccd1 _18885_/Y
+ sky130_fd_sc_hd__a2bb2oi_4
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17836_ _17540_/X _17686_/A _17832_/D _17835_/X vssd1 vssd1 vccd1 vccd1 _17836_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_120_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18007__D1 _17723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17767_ _17611_/X _17763_/X _17710_/X _17876_/B _17754_/Y vssd1 vssd1 vccd1 vccd1
+ _17767_/X sky130_fd_sc_hd__o311a_1
XFILLER_94_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14979_ _14178_/Y _14097_/X _14089_/Y _15488_/C vssd1 vssd1 vccd1 vccd1 _14979_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19506_ _19504_/X _19505_/X _12040_/X _18481_/B _19502_/A vssd1 vssd1 vccd1 vccd1
+ _19649_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_63_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16718_ _16722_/A _16950_/A _16722_/B _16722_/C vssd1 vssd1 vccd1 vccd1 _16718_/Y
+ sky130_fd_sc_hd__nand4_2
X_17698_ _17698_/A _17698_/B vssd1 vssd1 vccd1 vccd1 _17703_/B sky130_fd_sc_hd__nor2_2
XFILLER_23_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19770__A1 _19380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19437_ _19437_/A vssd1 vssd1 vccd1 vccd1 _19638_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16649_ _16649_/A _16649_/B vssd1 vssd1 vccd1 vccd1 _16650_/B sky130_fd_sc_hd__nand2_1
XFILLER_179_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19368_ _19363_/Y _19540_/A _19365_/Y _19900_/D _19705_/A vssd1 vssd1 vccd1 vccd1
+ _19369_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_50_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18319_ _18319_/A _18319_/B _18319_/C _18319_/D vssd1 vssd1 vccd1 vccd1 _18319_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21865__C1 _21971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20132__A2 _20055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19299_ _19094_/A _19094_/B _19442_/A vssd1 vssd1 vccd1 vccd1 _19299_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_198_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23580__CLK _23588_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21330_ _21330_/A _21330_/B _21330_/C vssd1 vssd1 vccd1 vccd1 _21331_/C sky130_fd_sc_hd__nand3_1
XFILLER_136_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18089__B2 _18211_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21261_ _23564_/Q _21144_/B _21249_/Y _21257_/Y _21258_/Y vssd1 vssd1 vccd1 vccd1
+ _21262_/B sky130_fd_sc_hd__o2111ai_2
XANTENNA__23082__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15828__A _16315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23000_ _23000_/A vssd1 vssd1 vccd1 vccd1 _23331_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__23467__D _23479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20212_ _20212_/A _20287_/A _20212_/C _20212_/D vssd1 vssd1 vccd1 vccd1 _20222_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_117_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21192_ _21493_/A _21493_/B _21295_/B vssd1 vssd1 vccd1 vccd1 _21192_/Y sky130_fd_sc_hd__nand3_4
XFILLER_190_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15847__B1 _15682_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20143_ _20146_/C _20146_/D _20138_/X vssd1 vssd1 vccd1 vccd1 _20143_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19038__B1 _19148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13322__A1 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12125__A2 _11841_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20074_ _19977_/Y _19974_/Y _19986_/B _20073_/X vssd1 vssd1 vccd1 vccd1 _20074_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1044 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16811__A2 _15766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22099__C _22099_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ _20978_/A _20978_/B vssd1 vssd1 vccd1 vccd1 _20984_/A sky130_fd_sc_hd__xor2_1
XFILLER_198_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19761__A1 _19554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22715_ _22716_/D _22564_/A _22564_/B _22789_/A _22716_/C vssd1 vssd1 vccd1 vccd1
+ _22717_/C sky130_fd_sc_hd__a32o_1
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22646_ _22646_/A vssd1 vssd1 vccd1 vccd1 _22830_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_1113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19513__A1 _16437_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20659__B1 _20894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22577_ _22577_/A _22577_/B vssd1 vssd1 vccd1 vccd1 _22577_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12330_ _12323_/X _12324_/X _12327_/Y _12329_/X vssd1 vssd1 vccd1 vccd1 _12330_/X
+ sky130_fd_sc_hd__o31a_1
X_21528_ _21528_/A _21528_/B _21528_/C vssd1 vssd1 vccd1 vccd1 _21529_/A sky130_fd_sc_hd__nand3_1
XFILLER_166_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15738__A _15738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ _18673_/A _11898_/X _12260_/Y vssd1 vssd1 vccd1 vccd1 _12273_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__23073__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21459_ _21377_/B _21378_/C _21455_/Y vssd1 vssd1 vccd1 vccd1 _21460_/B sky130_fd_sc_hd__a21o_1
XANTENNA__20363__B _20363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14000_ _23503_/Q vssd1 vssd1 vccd1 vccd1 _14162_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18485__D1 _19846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ _12281_/A _17642_/A _12178_/Y vssd1 vssd1 vccd1 vccd1 _12192_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14361__B _14980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15838__B1 _16062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput53 _23599_/X vssd1 vssd1 vccd1 vccd1 wb_ack_o sky130_fd_sc_hd__buf_2
X_23129_ _23129_/A vssd1 vssd1 vccd1 vccd1 _23388_/D sky130_fd_sc_hd__clkbuf_1
Xoutput64 _14676_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput75 _14714_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[29] sky130_fd_sc_hd__buf_2
Xoutput86 _23262_/Q vssd1 vssd1 vccd1 vccd1 y[0] sky130_fd_sc_hd__buf_2
Xoutput97 _23580_/Q vssd1 vssd1 vccd1 vccd1 y[9] sky130_fd_sc_hd__buf_2
X_15951_ _15946_/Y _15947_/X _15949_/X _15950_/Y vssd1 vssd1 vccd1 vccd1 _16002_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_89_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14902_ _14588_/X _14050_/X _14061_/X _14901_/X _14980_/A vssd1 vssd1 vccd1 vccd1
+ _14903_/B sky130_fd_sc_hd__o311a_1
XFILLER_62_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18670_ _18670_/A _18670_/B vssd1 vssd1 vccd1 vccd1 _18670_/Y sky130_fd_sc_hd__nor2_1
X_15882_ _15882_/A vssd1 vssd1 vccd1 vccd1 _15882_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_768 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17391__C _17391_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17621_ _17612_/X _17614_/X _17609_/A _17609_/B vssd1 vssd1 vccd1 vccd1 _17622_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_5_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14833_ _15195_/B vssd1 vssd1 vccd1 vccd1 _15054_/A sky130_fd_sc_hd__buf_2
XFILLER_64_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23453__CLK _23462_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14089__A _23495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _17549_/A _17393_/A _17550_/X _17551_/X vssd1 vssd1 vccd1 vccd1 _17791_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_14764_ _14764_/A _14764_/B vssd1 vssd1 vccd1 vccd1 _15301_/A sky130_fd_sc_hd__nand2_2
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _11902_/A _11902_/B _11902_/C _11912_/B _11912_/A vssd1 vssd1 vccd1 vccd1
+ _11976_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_440 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16503_ _15855_/Y _15856_/Y _16528_/B _16500_/Y _16501_/X vssd1 vssd1 vccd1 vccd1
+ _16503_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13715_ _13727_/A _13715_/B vssd1 vssd1 vccd1 vccd1 _13715_/X sky130_fd_sc_hd__or2_1
XFILLER_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17483_ _17483_/A vssd1 vssd1 vccd1 vccd1 _17497_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14695_ _23342_/Q _14689_/X _14694_/X _23310_/Q _14678_/X vssd1 vssd1 vccd1 vccd1
+ _14695_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_624 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19222_ _19219_/X _19220_/Y _19205_/X _19221_/Y vssd1 vssd1 vccd1 vccd1 _19222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16434_ _16572_/B _16428_/X _16433_/X vssd1 vssd1 vccd1 vccd1 _16435_/C sky130_fd_sc_hd__o21ai_2
X_13646_ _13646_/A _13646_/B _13646_/C vssd1 vssd1 vccd1 vccd1 _13671_/A sky130_fd_sc_hd__nand3_1
XANTENNA__22639__A1 _22644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12588__C1 _14655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16365_ _16365_/A _16821_/A _18481_/B vssd1 vssd1 vccd1 vccd1 _16366_/B sky130_fd_sc_hd__nand3_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ _19157_/A vssd1 vssd1 vccd1 vccd1 _19502_/A sky130_fd_sc_hd__clkbuf_4
X_13577_ _13569_/Y _13575_/Y _13576_/Y vssd1 vssd1 vccd1 vccd1 _13577_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_188_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18104_ _18104_/A _18104_/B _18179_/A vssd1 vssd1 vccd1 vccd1 _18179_/B sky130_fd_sc_hd__nand3_2
XFILLER_157_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15316_ _15316_/A vssd1 vssd1 vccd1 vccd1 _15419_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12528_ _12528_/A _12528_/B _12537_/B vssd1 vssd1 vccd1 vccd1 _12529_/C sky130_fd_sc_hd__nand3_1
XFILLER_158_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19084_ _19076_/Y _19080_/X _19091_/C _19083_/X vssd1 vssd1 vccd1 vccd1 _19094_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_145_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16296_ _16340_/C _16340_/A vssd1 vssd1 vccd1 vccd1 _16296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18035_ _17916_/B _17916_/C _17916_/A vssd1 vssd1 vccd1 vccd1 _18036_/B sky130_fd_sc_hd__a21boi_1
X_15247_ _15249_/A _15246_/Y _15187_/C vssd1 vssd1 vccd1 vccd1 _15247_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ _12104_/X _12107_/A _12110_/Y vssd1 vssd1 vccd1 vccd1 _12469_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__21075__B1 _20969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15178_ _15179_/B _15179_/C _15179_/A vssd1 vssd1 vccd1 vccd1 _15250_/A sky130_fd_sc_hd__a21o_1
XFILLER_158_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14271__B _14760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18959__A _18959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14129_ _14116_/X _14118_/X _14183_/A _14121_/Y _15082_/B vssd1 vssd1 vccd1 vccd1
+ _14130_/C sky130_fd_sc_hd__o2111ai_1
X_19986_ _19986_/A _19986_/B vssd1 vssd1 vccd1 vccd1 _19987_/C sky130_fd_sc_hd__nand2_1
XFILLER_140_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17582__B _18778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18937_ _18500_/X _18604_/X _18942_/A vssd1 vssd1 vccd1 vccd1 _19141_/A sky130_fd_sc_hd__o21ai_1
XFILLER_140_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16479__A _16479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21917__A3 _22270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11866__A1 _11864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18868_ _18868_/A _18868_/B _18868_/C vssd1 vssd1 vccd1 vccd1 _18868_/X sky130_fd_sc_hd__and3_2
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20050__A1 _20209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17819_ _18072_/D _18072_/C vssd1 vssd1 vccd1 vccd1 _18253_/A sky130_fd_sc_hd__nand2_2
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14804__A1 _14207_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18799_ _18799_/A _18799_/B vssd1 vssd1 vccd1 vccd1 _18800_/B sky130_fd_sc_hd__nand2_1
XFILLER_82_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20830_ _20961_/A _12648_/X _20529_/B _20678_/A _20829_/X vssd1 vssd1 vccd1 vccd1
+ _20887_/B sky130_fd_sc_hd__o32a_1
XFILLER_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20761_ _23561_/Q _20761_/B _20761_/C vssd1 vssd1 vccd1 vccd1 _20763_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__16557__A1 _16530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14727__A _23595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22500_ _22500_/A _22500_/B _22500_/C vssd1 vssd1 vccd1 vccd1 _22541_/C sky130_fd_sc_hd__nand3_1
XFILLER_51_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23480_ _23492_/CLK hold7/X vssd1 vssd1 vccd1 vccd1 _23480_/Q sky130_fd_sc_hd__dfxtp_2
X_20692_ _20691_/Y _20492_/B _20518_/X vssd1 vssd1 vccd1 vccd1 _20695_/A sky130_fd_sc_hd__a21boi_1
X_22431_ _22237_/A _21892_/X _22264_/Y vssd1 vssd1 vccd1 vccd1 _22434_/D sky130_fd_sc_hd__o21ai_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22362_ _22362_/A _22362_/B vssd1 vssd1 vccd1 vccd1 _22362_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16661__B _19308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21313_ _21312_/X _21195_/X _21386_/B _21307_/D vssd1 vssd1 vccd1 vccd1 _21317_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_190_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22293_ _22293_/A vssd1 vssd1 vccd1 vccd1 _22476_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__20183__B _20183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21244_ _21019_/C _21244_/B _21244_/C _21244_/D vssd1 vssd1 vccd1 vccd1 _21255_/A
+ sky130_fd_sc_hd__nand4b_1
XFILLER_105_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21175_ _21037_/A _21279_/C _21174_/Y vssd1 vssd1 vccd1 vccd1 _21179_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14099__A2 _14203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16493__B1 _16458_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20126_ _20201_/A _20201_/B _20310_/C _20201_/C vssd1 vssd1 vccd1 vccd1 _20128_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15835__A3 _17057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23476__CLK _23492_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20057_ _19807_/X _20045_/Y _19973_/X vssd1 vssd1 vccd1 vccd1 _20058_/B sky130_fd_sc_hd__o21ai_1
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _11830_/A vssd1 vssd1 vccd1 vccd1 _16027_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18537__A2 _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_771 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _18756_/B vssd1 vssd1 vccd1 vccd1 _12183_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20344__A2 _20295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20959_ _12689_/X _12850_/B _12815_/B _12692_/Y vssd1 vssd1 vccd1 vccd1 _20959_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_92_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16548__B2 _16549_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13500_ _23475_/Q vssd1 vssd1 vccd1 vccd1 _22064_/C sky130_fd_sc_hd__clkbuf_2
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14559__B1 _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14446_/Y _14452_/X _14441_/Y vssd1 vssd1 vccd1 vccd1 _14486_/C sky130_fd_sc_hd__a21boi_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _23586_/Q vssd1 vssd1 vccd1 vccd1 _11860_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_41_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _13431_/A vssd1 vssd1 vccd1 vccd1 _13431_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22629_ _22629_/A _22629_/B _22629_/C vssd1 vssd1 vccd1 vccd1 _22813_/A sky130_fd_sc_hd__nand3_1
XFILLER_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16150_ _16614_/A vssd1 vssd1 vccd1 vccd1 _16598_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13362_ _21767_/A _22039_/C vssd1 vssd1 vccd1 vccd1 _13362_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12294__A2_N _12297_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ _14860_/Y _15112_/B _14632_/X _13937_/X vssd1 vssd1 vccd1 vccd1 _15102_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_194_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12313_ _19653_/A vssd1 vssd1 vccd1 vccd1 _16529_/C sky130_fd_sc_hd__buf_2
XFILLER_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16081_ _16081_/A _16081_/B vssd1 vssd1 vccd1 vccd1 _16084_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15468__A _15538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13293_ _22562_/B vssd1 vssd1 vccd1 vccd1 _22361_/C sky130_fd_sc_hd__buf_2
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15032_ _15030_/X _15031_/Y _15035_/A _15035_/B vssd1 vssd1 vccd1 vccd1 _15033_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_181_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12244_ _11815_/X _16523_/A _16523_/B _16458_/A _12243_/X vssd1 vssd1 vccd1 vccd1
+ _12244_/X sky130_fd_sc_hd__o32a_1
XFILLER_6_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19840_ _19840_/A _20046_/A _20047_/A vssd1 vssd1 vccd1 vccd1 _19848_/A sky130_fd_sc_hd__nand3_1
XFILLER_122_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12175_ _12175_/A vssd1 vssd1 vccd1 vccd1 _12175_/X sky130_fd_sc_hd__buf_2
XFILLER_123_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19771_ _19932_/A _19771_/B _19771_/C _19932_/B vssd1 vssd1 vccd1 vccd1 _19771_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_150_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16983_ _16988_/A _16983_/B _16983_/C _17026_/B vssd1 vssd1 vccd1 vccd1 _16983_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18722_ _18722_/A vssd1 vssd1 vccd1 vccd1 _18722_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15934_ _16781_/B _15933_/Y _17137_/C vssd1 vssd1 vccd1 vccd1 _17885_/A sky130_fd_sc_hd__o21a_2
XFILLER_7_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12620__A _14655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18653_ _18798_/A _23394_/Q _18653_/C vssd1 vssd1 vccd1 vccd1 _18973_/B sky130_fd_sc_hd__nand3_2
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _15861_/X _16523_/C _12518_/X _16064_/A vssd1 vssd1 vccd1 vccd1 _15866_/B
+ sky130_fd_sc_hd__o22a_2
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_844 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _19709_/C vssd1 vssd1 vccd1 vccd1 _20055_/D sky130_fd_sc_hd__buf_4
XANTENNA__18945__C _18945_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14816_ _14816_/A _14816_/B _14816_/C _14816_/D vssd1 vssd1 vccd1 vccd1 _14825_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18584_ _18584_/A _18584_/B vssd1 vssd1 vccd1 vccd1 _18584_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _15796_/A _15796_/B _15796_/C vssd1 vssd1 vccd1 vccd1 _15894_/A sky130_fd_sc_hd__nand3_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23570__D _23570_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ _17535_/A vssd1 vssd1 vccd1 vccd1 _18207_/A sky130_fd_sc_hd__buf_2
XFILLER_33_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11959_ _11959_/A vssd1 vssd1 vccd1 vccd1 _16808_/A sky130_fd_sc_hd__buf_4
X_14747_ _15338_/A _23506_/Q vssd1 vssd1 vccd1 vccd1 _14961_/A sky130_fd_sc_hd__xor2_1
XFILLER_32_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17466_ _12088_/A _17465_/X _17460_/A vssd1 vssd1 vccd1 vccd1 _17562_/A sky130_fd_sc_hd__o21ai_1
X_14678_ _23040_/D vssd1 vssd1 vccd1 vccd1 _14678_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_616 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19205_ _19203_/X _17408_/X _19204_/X _19018_/X vssd1 vssd1 vccd1 vccd1 _19205_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_34_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16417_ _16421_/A _16475_/C _16418_/A vssd1 vssd1 vccd1 vccd1 _16472_/A sky130_fd_sc_hd__a21o_1
X_13629_ _21883_/A _22064_/C _21883_/C vssd1 vssd1 vccd1 vccd1 _13630_/B sky130_fd_sc_hd__nand3_2
XFILLER_158_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17397_ _17397_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17397_/Y sky130_fd_sc_hd__nand2_1
X_19136_ _19133_/A _19133_/B _19134_/A vssd1 vssd1 vccd1 vccd1 _19140_/A sky130_fd_sc_hd__o21ai_1
XFILLER_192_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16348_ _16348_/A _16348_/B _16348_/C vssd1 vssd1 vccd1 vccd1 _16581_/B sky130_fd_sc_hd__nand3_1
XFILLER_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19067_ _19065_/X _19066_/Y _19057_/D _19060_/B vssd1 vssd1 vccd1 vccd1 _19069_/B
+ sky130_fd_sc_hd__o211ai_4
X_16279_ _16281_/A _16281_/B _16281_/C _16281_/D vssd1 vssd1 vccd1 vccd1 _16282_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18018_ _18075_/A _18075_/B _18114_/A _18014_/B vssd1 vssd1 vccd1 vccd1 _18018_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17593__A _17593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19661__B1 _19846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19969_ _19969_/A vssd1 vssd1 vccd1 vccd1 _20268_/C sky130_fd_sc_hd__buf_2
XFILLER_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18216__A1 _17959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18216__B2 _18219_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11839__A1 _11834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22980_ _22980_/A vssd1 vssd1 vccd1 vccd1 _23322_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__19016__C _19148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21931_ _21939_/A _21939_/B _21940_/B vssd1 vssd1 vccd1 vccd1 _21936_/A sky130_fd_sc_hd__a21o_1
XFILLER_27_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21771__A1 _13642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12249__D1 _19180_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21862_ _21859_/A _21859_/B _22107_/D _22455_/A vssd1 vssd1 vccd1 vccd1 _21864_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_55_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20813_ _20957_/A _12862_/A _20805_/A vssd1 vssd1 vccd1 vccd1 _20819_/C sky130_fd_sc_hd__o21ai_1
XFILLER_24_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21793_ _21793_/A _21793_/B _21793_/C _21878_/A vssd1 vssd1 vccd1 vccd1 _21793_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13361__A _23471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23532_ _23538_/CLK _23532_/D vssd1 vssd1 vccd1 vccd1 _23532_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18684__A2_N _12185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20744_ _21008_/C _20577_/Y _20593_/C _20740_/Y _20743_/Y vssd1 vssd1 vccd1 vccd1
+ _21157_/A sky130_fd_sc_hd__o2111ai_2
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22079__A2 _21994_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23463_ _23559_/CLK _23475_/Q vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20675_ _20675_/A _20675_/B _23453_/Q vssd1 vssd1 vccd1 vccd1 _20676_/B sky130_fd_sc_hd__nand3_2
XFILLER_10_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22414_ _22383_/X _22389_/Y _22394_/Y vssd1 vssd1 vccd1 vccd1 _22414_/X sky130_fd_sc_hd__o21a_1
XFILLER_183_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23394_ _23395_/CLK _23394_/D vssd1 vssd1 vccd1 vccd1 _23394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23028__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22345_ _22344_/Y _22246_/Y _22439_/A vssd1 vssd1 vccd1 vccd1 _22445_/D sky130_fd_sc_hd__o21bai_1
XFILLER_136_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22276_ _22276_/A vssd1 vssd1 vccd1 vccd1 _22656_/B sky130_fd_sc_hd__buf_2
XFILLER_163_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11966__D _19334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21227_ _21165_/X _21162_/Y _21166_/Y _21221_/B _21221_/C vssd1 vssd1 vccd1 vccd1
+ _21228_/D sky130_fd_sc_hd__o2111ai_4
XANTENNA__21737__B _23326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21158_ _21158_/A _21158_/B _21158_/C _21241_/C vssd1 vssd1 vccd1 vccd1 _21158_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_78_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20109_ _20111_/A _20111_/D vssd1 vssd1 vccd1 vccd1 _20110_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16481__A3 _16451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13980_ _23502_/Q vssd1 vssd1 vccd1 vccd1 _14791_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_4_4_0_bq_clk_i_A clkbuf_4_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23200__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21089_ _21089_/A _21095_/A vssd1 vssd1 vccd1 vccd1 _21089_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12440__A _16661_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20014__A1 _19040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12931_ _20773_/C _12941_/A _20773_/A vssd1 vssd1 vccd1 vccd1 _13113_/C sky130_fd_sc_hd__nand3_2
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13255__B _13660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12862_ _12862_/A vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__clkbuf_4
X_15650_ _17098_/B _15928_/A _16677_/B _16661_/C vssd1 vssd1 vccd1 vccd1 _15650_/Y
+ sky130_fd_sc_hd__nand4_4
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20369__A _20369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _12144_/A vssd1 vssd1 vccd1 vccd1 _11814_/A sky130_fd_sc_hd__clkbuf_4
X_14601_ _23580_/Q _14551_/A _14587_/X _14188_/A vssd1 vssd1 vccd1 vccd1 _14601_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15581_ _23511_/Q _15585_/D _15586_/C vssd1 vssd1 vccd1 vccd1 _15582_/B sky130_fd_sc_hd__o21ai_1
XFILLER_73_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _12788_/B _12915_/A _12668_/X _12667_/B vssd1 vssd1 vccd1 vccd1 _13051_/C
+ sky130_fd_sc_hd__o211ai_2
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17320_ _18211_/D _16480_/X _17326_/C _17326_/B vssd1 vssd1 vccd1 vccd1 _17322_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14550_/A vssd1 vssd1 vccd1 vccd1 _14532_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _23382_/Q _11656_/B _11758_/A vssd1 vssd1 vccd1 vccd1 _11746_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__19877__B _19888_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17251_ _17249_/X _17250_/X _16308_/C _17569_/A vssd1 vssd1 vccd1 vccd1 _17433_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12007__A1 _12004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14463_ _13965_/X _13966_/X _15118_/A _13972_/X _14462_/Y vssd1 vssd1 vccd1 vccd1
+ _14463_/Y sky130_fd_sc_hd__o2111ai_2
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11675_ _11754_/A vssd1 vssd1 vccd1 vccd1 _11686_/B sky130_fd_sc_hd__buf_2
XFILLER_169_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13414_ _13414_/A _13414_/B _13414_/C vssd1 vssd1 vccd1 vccd1 _13460_/D sky130_fd_sc_hd__nand3_2
X_16202_ _15634_/C _15618_/A _15682_/B _15706_/A _15652_/A vssd1 vssd1 vccd1 vccd1
+ _16202_/Y sky130_fd_sc_hd__o2111ai_4
X_17182_ _16946_/X _16942_/X _17187_/A _17186_/A vssd1 vssd1 vccd1 vccd1 _17182_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14394_ _13890_/A _13890_/B _14105_/A vssd1 vssd1 vccd1 vccd1 _14395_/B sky130_fd_sc_hd__a21o_1
X_16133_ _16121_/Y _16610_/A _16124_/X vssd1 vssd1 vccd1 vccd1 _16135_/B sky130_fd_sc_hd__a21o_1
X_13345_ _13358_/A vssd1 vssd1 vccd1 vccd1 _21744_/C sky130_fd_sc_hd__buf_2
XANTENNA__23019__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _16064_/A vssd1 vssd1 vccd1 vccd1 _16066_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13276_ _23476_/Q vssd1 vssd1 vccd1 vccd1 _13642_/A sky130_fd_sc_hd__inv_2
XANTENNA__15901__C1 _16856_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22778__B1 _22858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15015_ _15015_/A _15015_/B _15015_/C vssd1 vssd1 vccd1 vccd1 _15035_/B sky130_fd_sc_hd__nand3_2
XFILLER_142_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12227_ _12227_/A _12227_/B _12227_/C vssd1 vssd1 vccd1 vccd1 _12532_/B sky130_fd_sc_hd__and3_1
XFILLER_170_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23565__D _23565_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12191__B1 _19485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19823_ _19823_/A _19823_/B vssd1 vssd1 vccd1 vccd1 _19823_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__21450__B1 _21376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12158_ _12158_/A vssd1 vssd1 vccd1 vccd1 _12199_/A sky130_fd_sc_hd__buf_2
XFILLER_190_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19754_ _19588_/Y _19570_/X _19733_/Y _19743_/X _19747_/A vssd1 vssd1 vccd1 vccd1
+ _19757_/B sky130_fd_sc_hd__o2111ai_1
X_16966_ _17899_/B vssd1 vssd1 vccd1 vccd1 _18161_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12089_ _12089_/A vssd1 vssd1 vccd1 vccd1 _12090_/A sky130_fd_sc_hd__clkbuf_2
X_18705_ _18707_/A _18707_/B _18706_/A _18892_/A vssd1 vssd1 vccd1 vccd1 _18709_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19946__A1 _18435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15917_ _11738_/X _11740_/X _11741_/Y _15668_/A _17233_/A vssd1 vssd1 vccd1 vccd1
+ _15917_/Y sky130_fd_sc_hd__o2111ai_4
X_19685_ _19685_/A _19685_/B _19685_/C vssd1 vssd1 vccd1 vccd1 _19688_/B sky130_fd_sc_hd__nand3_2
XANTENNA__17860__B _20142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16897_ _16054_/A _16055_/A _15922_/A _15937_/A vssd1 vssd1 vccd1 vccd1 _16913_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16757__A _16757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17421__A2 _16741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18675__C _18675_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18636_ _16044_/A _18461_/B _18460_/A _18635_/Y vssd1 vssd1 vccd1 vccd1 _18804_/A
+ sky130_fd_sc_hd__o31ai_4
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _16311_/A vssd1 vssd1 vccd1 vccd1 _16370_/A sky130_fd_sc_hd__buf_2
XFILLER_25_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18567_ _18545_/Y _18548_/Y _18557_/B _18728_/A vssd1 vssd1 vccd1 vccd1 _18568_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15779_ _16593_/D vssd1 vssd1 vccd1 vccd1 _17066_/C sky130_fd_sc_hd__buf_2
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19174__A2 _18455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17518_ _17353_/Y _17357_/Y _17362_/Y vssd1 vssd1 vccd1 vccd1 _17519_/B sky130_fd_sc_hd__o21a_1
XFILLER_177_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18498_ _18482_/Y _18487_/X _18458_/Y _18465_/A vssd1 vssd1 vccd1 vccd1 _18499_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_36_1127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17588__A _20142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17449_ _17449_/A vssd1 vssd1 vccd1 vccd1 _19534_/B sky130_fd_sc_hd__buf_2
XFILLER_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20460_ _12987_/Y _20459_/Y _13208_/B vssd1 vssd1 vccd1 vccd1 _20465_/A sky130_fd_sc_hd__a21o_1
XFILLER_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19119_ _17591_/A _17593_/A _12283_/Y _12282_/X _17595_/A vssd1 vssd1 vccd1 vccd1
+ _19119_/Y sky130_fd_sc_hd__o221ai_4
X_20391_ _23555_/Q vssd1 vssd1 vccd1 vccd1 _20393_/A sky130_fd_sc_hd__inv_2
XFILLER_119_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22130_ _22130_/A _22130_/B _22130_/C _22130_/D vssd1 vssd1 vccd1 vccd1 _22139_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_161_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22061_ _22061_/A _22061_/B _22061_/C vssd1 vssd1 vccd1 vccd1 _22061_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__19308__A _19652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18212__A _18277_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20461__B _23458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21012_ _21012_/A vssd1 vssd1 vccd1 vccd1 _21012_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13356__A _23326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12260__A _12306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22963_ _22963_/A vssd1 vssd1 vccd1 vccd1 _23315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22388__B _22388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19043__A _19043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21914_ _22040_/A vssd1 vssd1 vccd1 vccd1 _22045_/B sky130_fd_sc_hd__buf_2
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22894_ _22895_/A _22895_/B vssd1 vssd1 vccd1 vccd1 _23577_/D sky130_fd_sc_hd__nor2_1
XFILLER_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0_0_bq_clk_i clkbuf_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_167_1035 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21845_ _21843_/Y _21844_/X _21834_/Y vssd1 vssd1 vccd1 vccd1 _21847_/A sky130_fd_sc_hd__o21bai_1
XFILLER_71_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_730 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21776_ _13339_/X _22141_/A _21744_/B vssd1 vssd1 vccd1 vccd1 _21777_/B sky130_fd_sc_hd__o21ai_2
XFILLER_23_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23515_ _23518_/CLK input51/X vssd1 vssd1 vccd1 vccd1 _23515_/Q sky130_fd_sc_hd__dfxtp_1
X_20727_ _20886_/A _20726_/D _20862_/A _20707_/Y vssd1 vssd1 vccd1 vccd1 _20727_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23446_ _23492_/CLK _23446_/D vssd1 vssd1 vccd1 vccd1 _23446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20658_ _12792_/A _12722_/A _12754_/A _20645_/Y _20647_/Y vssd1 vssd1 vccd1 vccd1
+ _20666_/A sky130_fd_sc_hd__o221a_1
XFILLER_7_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_87 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18676__B2 _18474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23377_ _23377_/CLK _23377_/D vssd1 vssd1 vccd1 vccd1 _23377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20589_ _20589_/A _20736_/A _20589_/C vssd1 vssd1 vccd1 vccd1 _20589_/X sky130_fd_sc_hd__and3_1
XFILLER_180_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13130_ _21121_/A _13121_/C _12979_/A _13124_/C vssd1 vssd1 vccd1 vccd1 _13133_/A
+ sky130_fd_sc_hd__a31o_1
X_22328_ _22260_/X _22231_/A _22325_/Y _22327_/Y vssd1 vssd1 vccd1 vccd1 _22357_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_944 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_966 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _12887_/C _12894_/B _12894_/C vssd1 vssd1 vccd1 vccd1 _13061_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__19218__A _19218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22259_ _21850_/A _21850_/B _22117_/Y _22243_/Y _22246_/Y vssd1 vssd1 vccd1 vccd1
+ _22346_/B sky130_fd_sc_hd__a221o_1
XFILLER_151_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20371__B _20371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16439__B1 _16064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ _19157_/C vssd1 vssd1 vccd1 vccd1 _12306_/A sky130_fd_sc_hd__buf_4
XFILLER_2_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input48_A x[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16820_ _17050_/A _16819_/X _15863_/A vssd1 vssd1 vccd1 vccd1 _17041_/C sky130_fd_sc_hd__a21oi_1
XFILLER_94_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13266__A _23475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18776__B _18966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12601__C _12601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12476__A1 _18945_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16751_ _16585_/Y _16587_/Y _16744_/Y _16750_/Y vssd1 vssd1 vccd1 vccd1 _16778_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_111_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13963_ _13948_/X _14191_/A _14191_/B vssd1 vssd1 vccd1 vccd1 _14331_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__22932__A0 _20902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18495__C _18495_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15702_ _11625_/A _11741_/A _11733_/Y _12147_/A vssd1 vssd1 vccd1 vccd1 _15704_/A
+ sky130_fd_sc_hd__a31o_4
X_19470_ _19470_/A vssd1 vssd1 vccd1 vccd1 _19470_/Y sky130_fd_sc_hd__inv_2
X_12914_ _13101_/C _13101_/B vssd1 vssd1 vccd1 vccd1 _12985_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13894_ _14459_/A vssd1 vssd1 vccd1 vccd1 _14835_/C sky130_fd_sc_hd__clkbuf_2
X_16682_ _16911_/A _16911_/B _16900_/A _17149_/A _17420_/B vssd1 vssd1 vccd1 vccd1
+ _16682_/Y sky130_fd_sc_hd__o2111ai_4
X_18421_ _18430_/A _18420_/X _18407_/C _18408_/B vssd1 vssd1 vccd1 vccd1 _18423_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15633_ _15630_/Y _15631_/Y _15713_/B vssd1 vssd1 vccd1 vccd1 _15634_/B sky130_fd_sc_hd__o21ai_1
X_12845_ _12845_/A _12845_/B _12845_/C vssd1 vssd1 vccd1 vccd1 _12901_/B sky130_fd_sc_hd__nand3_2
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15965__A2 _17456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14097__A _14097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _18293_/A _18293_/B _18355_/A _18355_/B _18314_/C vssd1 vssd1 vccd1 vccd1
+ _18394_/B sky130_fd_sc_hd__o221ai_4
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15564_ _15564_/A _15564_/B vssd1 vssd1 vccd1 vccd1 _15564_/Y sky130_fd_sc_hd__nor2_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12776_/A _12776_/B vssd1 vssd1 vccd1 vccd1 _12779_/A sky130_fd_sc_hd__nand2_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17303_/A vssd1 vssd1 vccd1 vccd1 _18211_/D sky130_fd_sc_hd__buf_2
XFILLER_9_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14515_ input3/X vssd1 vssd1 vccd1 vccd1 _14633_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_42_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11727_ _18805_/A vssd1 vssd1 vccd1 vccd1 _16661_/C sky130_fd_sc_hd__clkbuf_4
X_18283_ _18324_/A _18335_/C _18324_/C _18339_/A vssd1 vssd1 vccd1 vccd1 _18284_/B
+ sky130_fd_sc_hd__a22oi_2
X_15495_ _15497_/B _15496_/A _15494_/X vssd1 vssd1 vccd1 vccd1 _15498_/A sky130_fd_sc_hd__a21boi_1
XFILLER_30_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17234_ _19494_/D _17766_/B _17766_/C _17236_/B _17236_/C vssd1 vssd1 vccd1 vccd1
+ _17238_/A sky130_fd_sc_hd__a32o_1
X_14446_ _14446_/A _14446_/B _14446_/C vssd1 vssd1 vccd1 vccd1 _14446_/Y sky130_fd_sc_hd__nand3_1
X_11658_ _23385_/Q _23384_/Q vssd1 vssd1 vccd1 vccd1 _11823_/B sky130_fd_sc_hd__nor2_4
XFILLER_70_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22999__A0 _23331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18016__B _18016_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17165_ _17166_/A _17166_/B _17350_/A _17170_/B vssd1 vssd1 vccd1 vccd1 _17167_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18667__A1 _18627_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14377_ _14377_/A _15082_/D _14377_/C vssd1 vssd1 vccd1 vccd1 _14492_/C sky130_fd_sc_hd__and3_1
XFILLER_70_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12345__A _18778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11589_ _11634_/A vssd1 vssd1 vccd1 vccd1 _12510_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16116_ _18169_/A vssd1 vssd1 vccd1 vccd1 _18219_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13328_ _21764_/C vssd1 vssd1 vccd1 vccd1 _22276_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12951__A2 _12637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17096_ _17096_/A vssd1 vssd1 vccd1 vccd1 _17096_/X sky130_fd_sc_hd__buf_2
XFILLER_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16047_ _16047_/A vssd1 vssd1 vccd1 vccd1 _16451_/C sky130_fd_sc_hd__clkbuf_4
X_13259_ _13259_/A vssd1 vssd1 vccd1 vccd1 _13377_/D sky130_fd_sc_hd__clkinv_2
XANTENNA__17890__A2 _17635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11911__B1 _11912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19806_ _17593_/X _17591_/X _17595_/X _20055_/A _20055_/B vssd1 vssd1 vccd1 vccd1
+ _19807_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23537__CLK _23538_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12080__A _18778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15094__C _15094_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17998_ _17852_/Y _17848_/X _17850_/Y _17867_/Y vssd1 vssd1 vccd1 vccd1 _17999_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15653__A1 _15621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19737_ _19734_/Y _19735_/Y _19736_/Y vssd1 vssd1 vccd1 vccd1 _19742_/A sky130_fd_sc_hd__o21ai_1
XFILLER_42_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16949_ _16953_/A _17173_/A _16953_/B _16953_/C vssd1 vssd1 vccd1 vccd1 _16949_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_38_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22923__A0 _14615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19668_ _19668_/A vssd1 vssd1 vccd1 vccd1 _19668_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18619_ _18619_/A _18619_/B _18619_/C vssd1 vssd1 vccd1 vccd1 _18715_/B sky130_fd_sc_hd__nand3_1
XFILLER_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19599_ _19755_/A _19755_/B _19609_/B _19598_/Y vssd1 vssd1 vccd1 vccd1 _19605_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21630_ _21630_/A _21630_/B vssd1 vssd1 vccd1 vccd1 _21631_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23113__A _23169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21561_ _21561_/A _21561_/B vssd1 vssd1 vccd1 vccd1 _21561_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15708__A2 _16802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14735__A _14735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23300_ _23300_/CLK _23300_/D vssd1 vssd1 vccd1 vccd1 _23300_/Q sky130_fd_sc_hd__dfxtp_4
X_20512_ _20512_/A _20512_/B vssd1 vssd1 vccd1 vccd1 _20515_/A sky130_fd_sc_hd__nand2_1
XFILLER_193_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21492_ _21561_/A _21561_/B _21491_/C vssd1 vssd1 vccd1 vccd1 _21495_/A sky130_fd_sc_hd__a21o_1
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23231_ _23434_/Q input19/X _23239_/S vssd1 vssd1 vccd1 vccd1 _23232_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14392__A1 _14433_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20443_ _20455_/A _20442_/B _20442_/C vssd1 vssd1 vccd1 vccd1 _20444_/B sky130_fd_sc_hd__o21a_1
XFILLER_193_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18658__A1 _11848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23162_ _23162_/A vssd1 vssd1 vccd1 vccd1 _23403_/D sky130_fd_sc_hd__clkbuf_1
X_20374_ _20322_/A _20322_/B _20269_/X vssd1 vssd1 vccd1 vccd1 _20428_/C sky130_fd_sc_hd__a21oi_2
XFILLER_173_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19870__A3 _17546_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22113_ _22113_/A _22451_/A vssd1 vssd1 vccd1 vccd1 _22115_/A sky130_fd_sc_hd__or2b_2
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23093_ _23373_/Q input22/X _23095_/S vssd1 vssd1 vccd1 vccd1 _23094_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14470__A _14819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22044_ _22035_/X _22041_/Y _22061_/C vssd1 vssd1 vccd1 vccd1 _22044_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_47_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19980__B _20146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17094__B1 _16591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_67 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22914__A0 _12675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_855 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22946_ _22946_/A vssd1 vssd1 vccd1 vccd1 _23307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_674 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21453__D _21453_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22390__A1 _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22877_ _22868_/B _22868_/A _22865_/B _22861_/X vssd1 vssd1 vccd1 vccd1 _22878_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_71_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12630_ _12604_/Y _12945_/B _12627_/X _12654_/A vssd1 vssd1 vccd1 vccd1 _12718_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_188_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21828_ _22420_/A vssd1 vssd1 vccd1 vccd1 _21829_/A sky130_fd_sc_hd__buf_2
XFILLER_71_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12561_ _12561_/A vssd1 vssd1 vccd1 vccd1 _19090_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16357__C1 _14735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21759_ _21759_/A _21759_/B _21759_/C vssd1 vssd1 vccd1 vccd1 _21760_/A sky130_fd_sc_hd__nand3_1
XFILLER_93_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20366__B _20366_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14300_ _14469_/D _15075_/B _14298_/A vssd1 vssd1 vccd1 vccd1 _14310_/C sky130_fd_sc_hd__a21o_1
XFILLER_54_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15280_ _15292_/A _15292_/B vssd1 vssd1 vccd1 vccd1 _15392_/A sky130_fd_sc_hd__nor2_1
X_12492_ _12491_/Y _12139_/Y _12157_/B vssd1 vssd1 vccd1 vccd1 _12492_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14231_ _14227_/A _14227_/B _14228_/A vssd1 vssd1 vccd1 vccd1 _14826_/B sky130_fd_sc_hd__o21ai_1
XFILLER_109_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23429_ _23429_/CLK _23429_/D vssd1 vssd1 vccd1 vccd1 _23429_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_153_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19874__C _20003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19310__A2 _19307_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14162_ _14167_/A _14162_/B _14360_/A _14167_/D vssd1 vssd1 vccd1 vccd1 _14162_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16124__A2 _11972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13113_ _13113_/A _13113_/B _13113_/C vssd1 vssd1 vccd1 vccd1 _13126_/C sky130_fd_sc_hd__nand3_1
XFILLER_166_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14093_ _14070_/X _13927_/A _15114_/B _14193_/C vssd1 vssd1 vccd1 vccd1 _14184_/A
+ sky130_fd_sc_hd__o211ai_4
X_18970_ _18796_/X _18790_/X _18792_/Y _18806_/B vssd1 vssd1 vccd1 vccd1 _18983_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_124_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17921_ _18045_/A vssd1 vssd1 vccd1 vccd1 _17922_/A sky130_fd_sc_hd__inv_2
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13044_/A _13044_/B vssd1 vssd1 vccd1 vccd1 _13044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17852_ _17750_/B _17745_/Y _17840_/B _17840_/A vssd1 vssd1 vccd1 vccd1 _17852_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__18821__A1 _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater102_A _23497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21925__B _21925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16803_ _16807_/A _16815_/D vssd1 vssd1 vccd1 vccd1 _16804_/B sky130_fd_sc_hd__and2_1
XFILLER_38_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17783_ _17747_/X _17758_/Y _17768_/Y _17771_/Y vssd1 vssd1 vccd1 vccd1 _17783_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15923__B _16198_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14995_ _14995_/A _14995_/B vssd1 vssd1 vccd1 vccd1 _15104_/A sky130_fd_sc_hd__nand2_1
XANTENNA__22905__A0 _12678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19522_ _19522_/A _19577_/B vssd1 vssd1 vccd1 vccd1 _19523_/A sky130_fd_sc_hd__nand2_1
X_16734_ _16268_/A _16268_/B _16268_/D _16260_/Y vssd1 vssd1 vccd1 vccd1 _16739_/A
+ sky130_fd_sc_hd__a31o_1
X_13946_ _13946_/A vssd1 vssd1 vccd1 vccd1 _14094_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19453_ _19451_/X _19453_/B _23545_/Q vssd1 vssd1 vccd1 vccd1 _19461_/A sky130_fd_sc_hd__nand3b_1
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16665_ _16665_/A vssd1 vssd1 vccd1 vccd1 _16665_/X sky130_fd_sc_hd__buf_2
X_13877_ _23350_/Q vssd1 vssd1 vccd1 vccd1 _14863_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__15938__A2 _17625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18404_ _18402_/Y _18403_/Y _18319_/Y _18264_/B _18367_/Y vssd1 vssd1 vccd1 vccd1
+ _18407_/D sky130_fd_sc_hd__o221ai_4
XFILLER_50_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15616_ _23417_/Q vssd1 vssd1 vccd1 vccd1 _15624_/A sky130_fd_sc_hd__inv_2
X_19384_ _19387_/B _19568_/A _19569_/A vssd1 vssd1 vccd1 vccd1 _19385_/C sky130_fd_sc_hd__nand3_1
X_12828_ _20532_/A _20532_/B _20528_/C vssd1 vssd1 vccd1 vccd1 _12828_/Y sky130_fd_sc_hd__nand3_1
X_16596_ _16601_/B _16601_/C _16595_/X vssd1 vssd1 vccd1 vccd1 _16597_/C sky130_fd_sc_hd__a21o_1
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18335_ _18378_/C _18335_/B _18335_/C _18335_/D vssd1 vssd1 vccd1 vccd1 _18378_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12082__C1 _16807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15547_ _15525_/B _15525_/A _15548_/A vssd1 vssd1 vccd1 vccd1 _15547_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12621__A1 _12667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _23451_/Q vssd1 vssd1 vccd1 vccd1 _20801_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_187_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18266_ _23534_/Q vssd1 vssd1 vccd1 vccd1 _18309_/A sky130_fd_sc_hd__inv_2
XFILLER_187_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_574 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15478_ _15478_/A _15527_/A _15478_/C vssd1 vssd1 vccd1 vccd1 _15479_/B sky130_fd_sc_hd__or3_1
X_17217_ _17217_/A vssd1 vssd1 vccd1 vccd1 _17535_/A sky130_fd_sc_hd__clkbuf_2
X_14429_ _14429_/A vssd1 vssd1 vccd1 vccd1 _15238_/C sky130_fd_sc_hd__buf_2
X_18197_ _18069_/Y _18070_/Y _18072_/B _18059_/A vssd1 vssd1 vccd1 vccd1 _18252_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__20447__A1 _20031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17148_ _17148_/A vssd1 vssd1 vccd1 vccd1 _17712_/D sky130_fd_sc_hd__buf_4
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17079_ _17089_/A _17089_/B _17079_/C _17079_/D vssd1 vssd1 vccd1 vccd1 _17221_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12803__A _13051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19065__A1 _19046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20090_ _20090_/A _20090_/B _20078_/A vssd1 vssd1 vccd1 vccd1 _20175_/C sky130_fd_sc_hd__nor3b_2
XFILLER_131_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22012__A _22564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22800_ _22800_/A _22800_/B _22800_/C vssd1 vssd1 vccd1 vccd1 _22800_/X sky130_fd_sc_hd__and3_1
XFILLER_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20992_ _20989_/A _20989_/B _20990_/A vssd1 vssd1 vccd1 vccd1 _20995_/A sky130_fd_sc_hd__o21ai_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22731_ _22731_/A _22731_/B vssd1 vssd1 vccd1 vccd1 _22731_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16051__A1 _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19321__A _19321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22662_ _22565_/Y _22572_/Y _22582_/X vssd1 vssd1 vccd1 vccd1 _22663_/C sky130_fd_sc_hd__o21ai_1
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21613_ _21630_/B vssd1 vssd1 vccd1 vccd1 _21666_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_179_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22593_ _22549_/A _22549_/B _22598_/A _22591_/A vssd1 vssd1 vccd1 vccd1 _22594_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17000__B1 _23522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21544_ _21544_/A _21512_/B vssd1 vssd1 vccd1 vccd1 _21566_/A sky130_fd_sc_hd__or2b_1
XFILLER_139_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17551__A1 _12279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14184__B _14184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21475_ _21404_/B _21404_/A _21335_/A _21354_/X vssd1 vssd1 vccd1 vccd1 _21477_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_14_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23214_ _23214_/A vssd1 vssd1 vccd1 vccd1 _23426_/D sky130_fd_sc_hd__clkbuf_1
X_20426_ _16816_/Y _16796_/X _16794_/B _17050_/X _20368_/D vssd1 vssd1 vccd1 vccd1
+ _20426_/X sky130_fd_sc_hd__a221o_1
XFILLER_107_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23145_ _23396_/Q input12/X _23145_/S vssd1 vssd1 vccd1 vccd1 _23146_/A sky130_fd_sc_hd__mux2_1
X_20357_ _23554_/Q vssd1 vssd1 vccd1 vccd1 _20357_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15727__C _16798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12128__B1 _12051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15865__A1 _15861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15865__B2 _16064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23076_ _15338_/A input13/X _23084_/S vssd1 vssd1 vccd1 vccd1 _23077_/A sky130_fd_sc_hd__mux2_1
X_20288_ _20287_/A _20287_/B _20287_/C _20284_/X vssd1 vssd1 vccd1 vccd1 _20288_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22027_ _22039_/B vssd1 vssd1 vccd1 vccd1 _22381_/B sky130_fd_sc_hd__buf_2
XFILLER_49_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13247__C _13523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_195_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17082__A3 _16451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19359__A2 _17846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13800_ _13430_/A _13410_/A _13797_/A vssd1 vssd1 vccd1 vccd1 _13812_/A sky130_fd_sc_hd__o21ai_2
XFILLER_17_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14780_ _14245_/A _14773_/Y _14775_/Y _14779_/X vssd1 vssd1 vccd1 vccd1 _14781_/B
+ sky130_fd_sc_hd__o211ai_1
X_11992_ _18468_/A vssd1 vssd1 vccd1 vccd1 _12099_/D sky130_fd_sc_hd__clkinv_2
XFILLER_112_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13731_ _13741_/B _13741_/C _13701_/Y _13415_/X vssd1 vssd1 vccd1 vccd1 _13731_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22929_ _23300_/Q input12/X _22929_/S vssd1 vssd1 vccd1 vccd1 _22930_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16450_ _16441_/Y _16507_/A _16448_/X _16449_/X vssd1 vssd1 vccd1 vccd1 _16450_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_16_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13662_ _13243_/Y _13658_/Y _22564_/C _13497_/A _13661_/Y vssd1 vssd1 vccd1 vccd1
+ _13666_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_72_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _15442_/C _15401_/B vssd1 vssd1 vccd1 vccd1 _23278_/D sky130_fd_sc_hd__xor2_1
X_12613_ _20528_/B vssd1 vssd1 vccd1 vccd1 _13121_/B sky130_fd_sc_hd__buf_2
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16381_ _16404_/A _16404_/B _16380_/Y vssd1 vssd1 vccd1 vccd1 _16381_/Y sky130_fd_sc_hd__a21oi_1
X_13593_ _13755_/A _13755_/B _13755_/C vssd1 vssd1 vccd1 vccd1 _13593_/X sky130_fd_sc_hd__and3_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _18132_/B vssd1 vssd1 vccd1 vccd1 _18133_/B sky130_fd_sc_hd__inv_2
XANTENNA__18334__A3 _17723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19531__A2 _17443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12544_ _12541_/Y _12542_/Y _12398_/C _12543_/Y vssd1 vssd1 vccd1 vccd1 _12557_/A
+ sky130_fd_sc_hd__o22ai_4
X_15332_ _15332_/A _15332_/B vssd1 vssd1 vccd1 vccd1 _15332_/X sky130_fd_sc_hd__xor2_2
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20141__A3 _20080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_73 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18051_ _18058_/D _18139_/B _17933_/X _18058_/A _18050_/Y vssd1 vssd1 vccd1 vccd1
+ _18051_/Y sky130_fd_sc_hd__a41oi_1
X_12475_ _18859_/A _12475_/B _19659_/C _18531_/A vssd1 vssd1 vccd1 vccd1 _12475_/X
+ sky130_fd_sc_hd__and4_1
X_15263_ _15263_/A vssd1 vssd1 vccd1 vccd1 _15409_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17002_ _16989_/A _16762_/Y _16776_/Y _17376_/A vssd1 vssd1 vccd1 vccd1 _17003_/B
+ sky130_fd_sc_hd__a22o_1
X_14214_ _14219_/C _14219_/D vssd1 vssd1 vccd1 vccd1 _14221_/B sky130_fd_sc_hd__nand2_2
XANTENNA__18098__A2 _17465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ _15193_/B _15193_/C _15193_/A vssd1 vssd1 vccd1 vccd1 _15203_/B sky130_fd_sc_hd__a21o_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14145_ _14090_/X _14098_/X _14084_/X _14101_/Y vssd1 vssd1 vccd1 vccd1 _14222_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_141_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18953_ _11834_/A _11834_/B _17966_/A _17966_/B vssd1 vssd1 vccd1 vccd1 _18953_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output79_A _14567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14076_ _14796_/A _14312_/D _14790_/C vssd1 vssd1 vccd1 vccd1 _14163_/B sky130_fd_sc_hd__and3_1
XFILLER_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13438__B _13810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21929__A1 _13469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17904_ _17868_/Y _17873_/Y _17901_/A _17901_/B _17881_/Y vssd1 vssd1 vccd1 vccd1
+ _17905_/C sky130_fd_sc_hd__o221ai_1
XFILLER_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22051__B1 _13453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ _13027_/A _13027_/B vssd1 vssd1 vccd1 vccd1 _20556_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12134__A3 _19308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18884_ _18884_/A _18884_/B vssd1 vssd1 vccd1 vccd1 _18884_/Y sky130_fd_sc_hd__nor2_2
XFILLER_94_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16749__B _18157_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17835_ _17705_/B _17680_/C _17834_/Y vssd1 vssd1 vccd1 vccd1 _17835_/X sky130_fd_sc_hd__a21o_1
XFILLER_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18007__C1 _17712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17766_ _17960_/A _17766_/B _17766_/C vssd1 vssd1 vccd1 vccd1 _17876_/B sky130_fd_sc_hd__and3_1
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14978_ _14978_/A vssd1 vssd1 vccd1 vccd1 _15488_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19505_ _19505_/A vssd1 vssd1 vccd1 vccd1 _19505_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16717_ _16957_/A _16956_/A _16956_/B vssd1 vssd1 vccd1 vccd1 _16722_/C sky130_fd_sc_hd__nand3_1
XANTENNA__12842__A1 _13131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13929_ _14172_/B vssd1 vssd1 vccd1 vccd1 _15353_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__20346__B1_N _23554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17697_ _17951_/D _17951_/A vssd1 vssd1 vccd1 vccd1 _23587_/D sky130_fd_sc_hd__xor2_2
XFILLER_179_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19436_ _19428_/A _19616_/A _19616_/B vssd1 vssd1 vccd1 vccd1 _19436_/X sky130_fd_sc_hd__a21o_1
X_16648_ _16853_/A _16649_/B _16644_/A vssd1 vssd1 vccd1 vccd1 _16648_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14595__A1 _14070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19367_ _19040_/X _17763_/A _19371_/A vssd1 vssd1 vccd1 vccd1 _19369_/B sky130_fd_sc_hd__o21ai_1
X_16579_ _16582_/C _16351_/Y _16765_/A _17009_/B vssd1 vssd1 vccd1 vccd1 _17026_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__14595__B2 _12121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18318_ _18318_/A _18318_/B vssd1 vssd1 vccd1 vccd1 _23594_/D sky130_fd_sc_hd__xnor2_1
XFILLER_148_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19298_ _19298_/A _19298_/B vssd1 vssd1 vccd1 vccd1 _19298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20132__A3 _20055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18249_ _18241_/Y _18243_/Y _18293_/A _18267_/A vssd1 vssd1 vccd1 vccd1 _18295_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_814 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21260_ _21249_/Y _21257_/Y _21259_/X vssd1 vssd1 vccd1 vccd1 _21260_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20211_ _18100_/A _20320_/B _20320_/C _20268_/C _18218_/A vssd1 vssd1 vccd1 vccd1
+ _20212_/C sky130_fd_sc_hd__a32o_1
XFILLER_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13570__A2 _22380_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21191_ _20906_/X _20907_/X _13131_/A _20908_/X vssd1 vssd1 vccd1 vccd1 _21191_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_132_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15847__A1 _15920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20142_ _20142_/A _20142_/B _20142_/C _20142_/D vssd1 vssd1 vccd1 vccd1 _20146_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19038__A1 _19148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22042__B1 _21913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13322__A2 _13226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20073_ _20073_/A _20073_/B _20073_/C vssd1 vssd1 vccd1 vccd1 _20073_/X sky130_fd_sc_hd__and3_1
XFILLER_131_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23483__D _23495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_9_0_bq_clk_i_A clkbuf_4_9_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18549__B1 _18526_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20975_ _20975_/A _20975_/B vssd1 vssd1 vccd1 vccd1 _20978_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17757__D1 _20217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19761__A2 _19534_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22714_ _22713_/C _22392_/A _22392_/B _22713_/D _22713_/A vssd1 vssd1 vccd1 vccd1
+ _22716_/C sky130_fd_sc_hd__a32o_1
XFILLER_198_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17772__A1 _17747_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22645_ _22830_/A _22461_/X _22641_/A vssd1 vssd1 vccd1 vccd1 _22649_/A sky130_fd_sc_hd__o21ai_1
XFILLER_41_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19201__D _19847_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19513__A2 _19858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12597__B1 _12601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22576_ _22559_/X _22478_/X _22565_/Y _22572_/Y _22663_/B vssd1 vssd1 vccd1 vccd1
+ _22584_/B sky130_fd_sc_hd__o221ai_1
XFILLER_178_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21527_ _21342_/Y _21343_/Y _21346_/A vssd1 vssd1 vccd1 vccd1 _21528_/A sky130_fd_sc_hd__a21oi_1
XFILLER_142_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12349__B1 _12348_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ _12306_/A _17149_/A _12260_/C _12260_/D vssd1 vssd1 vccd1 vccd1 _12260_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21458_ _21513_/A _21456_/Y _21460_/C vssd1 vssd1 vccd1 vccd1 _21463_/C sky130_fd_sc_hd__o21bai_1
XFILLER_119_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20409_ _20409_/A _20409_/B vssd1 vssd1 vccd1 vccd1 _20411_/C sky130_fd_sc_hd__or2_1
XANTENNA__18485__C1 _15704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ _11935_/X _12171_/Y _19485_/A _12308_/A _12177_/Y vssd1 vssd1 vccd1 vccd1
+ _12191_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21389_ _21389_/A _21389_/B vssd1 vssd1 vccd1 vccd1 _21391_/C sky130_fd_sc_hd__nor2_1
XFILLER_162_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21178__D _21279_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23128_ _11665_/A input35/X _23134_/S vssd1 vssd1 vccd1 vccd1 _23129_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput54 _14542_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_96_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput65 _14556_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput76 _14561_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput87 _23581_/Q vssd1 vssd1 vccd1 vccd1 y[10] sky130_fd_sc_hd__buf_2
XFILLER_110_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23059_ _23059_/A vssd1 vssd1 vccd1 vccd1 _23357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15950_ _15948_/A _16246_/B _15948_/C vssd1 vssd1 vccd1 vccd1 _15950_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12521__B1 _12522_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A wb_dat_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14901_ _14901_/A vssd1 vssd1 vccd1 vccd1 _14901_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15881_ _15750_/Y _15754_/X _15759_/X vssd1 vssd1 vccd1 vccd1 _15886_/B sky130_fd_sc_hd__a21bo_1
XFILLER_23_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17620_ _17609_/A _17609_/B _17618_/X _17619_/X vssd1 vssd1 vccd1 vccd1 _17622_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14832_ _23505_/Q vssd1 vssd1 vccd1 vccd1 _15195_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23182__S _23182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17551_ _12279_/X _17506_/A _17891_/A _17546_/C vssd1 vssd1 vccd1 vccd1 _17551_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11627__A2 _16619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14763_ _14756_/Y _14757_/Y _14754_/X vssd1 vssd1 vccd1 vccd1 _14766_/A sky130_fd_sc_hd__o21ai_1
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _11902_/B _11902_/C _11902_/A vssd1 vssd1 vccd1 vccd1 _11975_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _12346_/A _15974_/C _15682_/D _16500_/Y _16501_/X vssd1 vssd1 vccd1 vccd1
+ _16502_/X sky130_fd_sc_hd__a32o_1
XFILLER_44_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13714_ _13585_/A _22553_/D _13582_/B _22465_/D vssd1 vssd1 vccd1 vccd1 _13715_/B
+ sky130_fd_sc_hd__a22oi_1
X_17482_ _17482_/A _17482_/B _17482_/C vssd1 vssd1 vccd1 vccd1 _17483_/A sky130_fd_sc_hd__nand3_1
XFILLER_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14694_ _22896_/D vssd1 vssd1 vccd1 vccd1 _14694_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19221_ _19221_/A _19221_/B _19221_/C vssd1 vssd1 vccd1 vccd1 _19221_/Y sky130_fd_sc_hd__nand3_1
XFILLER_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14817__B _23505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16433_ _16757_/C vssd1 vssd1 vccd1 vccd1 _16433_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14577__A1 _23267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14577__B2 _12608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13645_ _13645_/A _13645_/B _13645_/C vssd1 vssd1 vccd1 vccd1 _13646_/C sky130_fd_sc_hd__nand3_2
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12588__B1 _12678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19152_ _18975_/X _18978_/B _18984_/Y vssd1 vssd1 vccd1 vccd1 _19167_/A sky130_fd_sc_hd__a21oi_1
X_16364_ _16364_/A _16364_/B _17041_/B vssd1 vssd1 vccd1 vccd1 _16364_/X sky130_fd_sc_hd__and3_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13576_ _13569_/B _13569_/C _13569_/A vssd1 vssd1 vccd1 vccd1 _13576_/Y sky130_fd_sc_hd__a21oi_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _18098_/X _18103_/B _18103_/C vssd1 vssd1 vccd1 vccd1 _18179_/A sky130_fd_sc_hd__nand3b_2
XFILLER_173_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15315_ _15237_/A _15237_/B _15245_/C vssd1 vssd1 vccd1 vccd1 _15315_/X sky130_fd_sc_hd__a21o_1
X_19083_ _19087_/A _19087_/B _19082_/X vssd1 vssd1 vccd1 vccd1 _19083_/X sky130_fd_sc_hd__a21o_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ _12527_/A vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16295_ _16326_/A _16096_/A _16097_/Y _16091_/Y vssd1 vssd1 vccd1 vccd1 _16340_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__23568__D _23568_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18034_ _18037_/B _18037_/C vssd1 vssd1 vccd1 vccd1 _18036_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_847 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15246_ _15179_/B _15179_/C _15179_/A vssd1 vssd1 vccd1 vccd1 _15246_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12458_ _12490_/A _12490_/B vssd1 vssd1 vccd1 vccd1 _12481_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13449__A _23475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21075__B2 _12722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12353__A _12353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12389_ _11908_/A _11908_/B _12061_/Y _12388_/Y vssd1 vssd1 vccd1 vccd1 _12396_/A
+ sky130_fd_sc_hd__o22ai_4
X_15177_ _15000_/B _15096_/Y _15107_/C vssd1 vssd1 vccd1 vccd1 _15179_/A sky130_fd_sc_hd__o21ai_1
XFILLER_126_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14271__C _14777_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15829__A1 _11766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18959__B _18959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14128_ _14128_/A vssd1 vssd1 vccd1 vccd1 _15082_/B sky130_fd_sc_hd__clkbuf_2
X_19985_ _19985_/A _19985_/B vssd1 vssd1 vccd1 vccd1 _19986_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18678__C _18859_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15664__A _15664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18936_ _18755_/Y _18934_/Y _18938_/A vssd1 vssd1 vccd1 vccd1 _18942_/A sky130_fd_sc_hd__o21ai_1
X_14059_ _14058_/X _13943_/X _13954_/Y vssd1 vssd1 vccd1 vccd1 _14284_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__17582__C _18778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18867_ _18782_/X _18786_/Y _18864_/Y _18866_/Y vssd1 vssd1 vccd1 vccd1 _18867_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11866__A2 _11865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20050__A2 _17600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13184__A _13184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17818_ _17686_/X _17541_/Y _17680_/C _17821_/B vssd1 vssd1 vccd1 vccd1 _18072_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__17451__B1 _16479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16198__C _16198_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13068__A1 _13131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18798_ _18798_/A _18798_/B vssd1 vssd1 vccd1 vccd1 _18799_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14804__A2 _14212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17749_ _17285_/X _17980_/A _17840_/A _17840_/B _17745_/Y vssd1 vssd1 vccd1 vccd1
+ _17751_/B sky130_fd_sc_hd__o221ai_1
XFILLER_78_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20760_ _20751_/Y _20754_/X _21542_/A _20759_/X vssd1 vssd1 vccd1 vccd1 _20761_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_165_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19419_ _19406_/A _19422_/B _19410_/X _19409_/X vssd1 vssd1 vccd1 vccd1 _19423_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_168_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14568__A1 input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14568__B2 _12601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20691_ _20501_/X _20520_/Y _20521_/Y vssd1 vssd1 vccd1 vccd1 _20691_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22430_ _22430_/A _22430_/B _22430_/C vssd1 vssd1 vccd1 vccd1 _22524_/A sky130_fd_sc_hd__nand3_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22361_ _22564_/A _22564_/B _22361_/C vssd1 vssd1 vccd1 vccd1 _22362_/B sky130_fd_sc_hd__nand3_4
XFILLER_175_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18215__A _19967_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_836 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21312_ _21365_/A _21455_/A _21435_/C _21497_/A vssd1 vssd1 vccd1 vccd1 _21312_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__16661__C _16661_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22292_ _22292_/A vssd1 vssd1 vccd1 vccd1 _22476_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21243_ _21243_/A _21243_/B vssd1 vssd1 vccd1 vccd1 _21244_/D sky130_fd_sc_hd__nand2_1
XFILLER_191_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20813__A1 _20957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21174_ _21174_/A _21174_/B _21174_/C vssd1 vssd1 vccd1 vccd1 _21174_/Y sky130_fd_sc_hd__nand3_1
XFILLER_105_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20125_ _20121_/X _20124_/X _23550_/Q _20119_/Y vssd1 vssd1 vccd1 vccd1 _20201_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_131_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16493__B2 _16478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22015__B1 _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21295__B _21295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12503__B1 _11721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20056_ _20056_/A _20056_/B vssd1 vssd1 vccd1 vccd1 _20060_/A sky130_fd_sc_hd__nand2_1
XFILLER_133_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11607__A _23397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12806__A1 _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11760_/A _11760_/B vssd1 vssd1 vccd1 vccd1 _18756_/B sky130_fd_sc_hd__nor2_4
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ _20957_/X _12862_/X _12877_/Y _21278_/A vssd1 vssd1 vccd1 vccd1 _20973_/B
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__17745__A1 _16479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16548__A2 _16549_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14559__A1 _23264_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11691_ _18849_/C vssd1 vssd1 vccd1 vccd1 _18859_/B sky130_fd_sc_hd__buf_2
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14559__B2 _15662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15756__B1 _15762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20889_ _20769_/A _13121_/A _13121_/B _21121_/B _21121_/C vssd1 vssd1 vccd1 vccd1
+ _21124_/A sky130_fd_sc_hd__a32o_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13430_ _13430_/A vssd1 vssd1 vccd1 vccd1 _13732_/A sky130_fd_sc_hd__buf_2
X_22628_ _22628_/A vssd1 vssd1 vccd1 vccd1 _23567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13361_ _23471_/Q vssd1 vssd1 vccd1 vccd1 _22039_/C sky130_fd_sc_hd__buf_2
XANTENNA__15749__A _15749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22559_ _22716_/A _22756_/B _22700_/D _22700_/C vssd1 vssd1 vccd1 vccd1 _22559_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_195_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14653__A _22028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15100_ _13937_/X _14870_/Y _14632_/X vssd1 vssd1 vccd1 vccd1 _15102_/A sky130_fd_sc_hd__o21ai_1
XFILLER_181_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12312_ _17149_/A vssd1 vssd1 vccd1 vccd1 _19653_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11996__B _12187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16080_ _15889_/X _15890_/Y _15867_/Y _15891_/Y vssd1 vssd1 vccd1 vccd1 _16081_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_13292_ _23477_/Q vssd1 vssd1 vccd1 vccd1 _22562_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_181_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16720__A2 _16176_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12243_ _18675_/B vssd1 vssd1 vccd1 vccd1 _12243_/X sky130_fd_sc_hd__buf_2
X_15031_ _15077_/A _15030_/B _15030_/C vssd1 vssd1 vccd1 vccd1 _15031_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_142_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_774 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_711 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12174_ _12174_/A vssd1 vssd1 vccd1 vccd1 _12174_/X sky130_fd_sc_hd__buf_2
XFILLER_174_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19770_ _19380_/X _19764_/Y _19621_/X _19769_/Y _19620_/X vssd1 vssd1 vccd1 vccd1
+ _19770_/X sky130_fd_sc_hd__o311a_1
X_16982_ _17365_/C _17026_/C _17026_/D _17369_/A vssd1 vssd1 vccd1 vccd1 _16982_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18721_ _18721_/A _18721_/B vssd1 vssd1 vccd1 vccd1 _18722_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_584 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15933_ _15604_/X _15605_/A _15599_/X _15921_/C vssd1 vssd1 vccd1 vccd1 _15933_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_114_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1092 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18652_ _18972_/B vssd1 vssd1 vccd1 vccd1 _20046_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _15864_/A vssd1 vssd1 vccd1 vccd1 _16064_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22309__A1 _22045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _17761_/B vssd1 vssd1 vccd1 vccd1 _19709_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14815_ _14227_/A _14227_/B _14215_/Y _14218_/Y vssd1 vssd1 vccd1 vccd1 _14816_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_92_856 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18583_ _18571_/Y _18572_/X _12563_/Y _12561_/A vssd1 vssd1 vccd1 vccd1 _18586_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15795_ _15782_/Y _15785_/Y _15946_/A _15794_/Y vssd1 vssd1 vccd1 vccd1 _15796_/C
+ sky130_fd_sc_hd__o211ai_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _17534_/A _17534_/B vssd1 vssd1 vccd1 vccd1 _23586_/D sky130_fd_sc_hd__xnor2_2
XFILLER_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13732__A _13732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14746_ _11633_/Y _23256_/A _14738_/A vssd1 vssd1 vccd1 vccd1 _23269_/D sky130_fd_sc_hd__a21oi_1
X_11958_ _11625_/A _11711_/B _16802_/B _16141_/A _16800_/A vssd1 vssd1 vccd1 vccd1
+ _11958_/X sky130_fd_sc_hd__a41o_1
XANTENNA__21371__D _21440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22190__C1 _21853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_254 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17465_ _17465_/A vssd1 vssd1 vccd1 vccd1 _17465_/X sky130_fd_sc_hd__buf_2
X_14677_ _14698_/A vssd1 vssd1 vccd1 vccd1 _14677_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11889_ _12016_/A _12016_/B _12032_/A vssd1 vssd1 vccd1 vccd1 _11891_/A sky130_fd_sc_hd__o21ai_2
XFILLER_189_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19204_ _19196_/A _19218_/A _15882_/X _19803_/A vssd1 vssd1 vccd1 vccd1 _19204_/X
+ sky130_fd_sc_hd__o22a_1
X_16416_ _16517_/B _16476_/D vssd1 vssd1 vccd1 vccd1 _16416_/X sky130_fd_sc_hd__and2_1
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19489__A1 _11926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13628_ _13621_/Y _13625_/X _13626_/Y _13627_/Y vssd1 vssd1 vccd1 vccd1 _13645_/B
+ sky130_fd_sc_hd__o211ai_4
X_17396_ _17810_/C _17810_/D _17810_/A vssd1 vssd1 vccd1 vccd1 _17806_/A sky130_fd_sc_hd__and3_2
XFILLER_158_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19135_ _19409_/A _19409_/B _19409_/C vssd1 vssd1 vccd1 vccd1 _19135_/Y sky130_fd_sc_hd__nand3_1
XFILLER_146_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16347_ _16347_/A _16347_/B _16347_/C vssd1 vssd1 vccd1 vccd1 _16348_/C sky130_fd_sc_hd__nand3_1
XFILLER_158_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13559_ _13634_/B vssd1 vssd1 vccd1 vccd1 _21988_/B sky130_fd_sc_hd__buf_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19066_ _19066_/A _19066_/B vssd1 vssd1 vccd1 vccd1 _19066_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18700__A3 _18499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_bq_clk_i clkbuf_2_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_157_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16278_ _16106_/Y _16350_/A _16273_/X vssd1 vssd1 vccd1 vccd1 _16278_/Y sky130_fd_sc_hd__o21ai_2
X_18017_ _18163_/B _18017_/B _18017_/C _18017_/D vssd1 vssd1 vccd1 vccd1 _18075_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_172_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15229_ _15227_/Y _15228_/X _14834_/A _15388_/C vssd1 vssd1 vccd1 vccd1 _15293_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19968_ _19967_/D _19967_/B _19203_/X _18097_/A vssd1 vssd1 vccd1 vccd1 _19985_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_141_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18216__A2 _17959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18919_ _19443_/A vssd1 vssd1 vccd1 vccd1 _18919_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11839__A2 _11834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19899_ _20017_/A _20017_/B _20017_/C vssd1 vssd1 vccd1 vccd1 _19899_/Y sky130_fd_sc_hd__nand3_2
XFILLER_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16227__A1 _16225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_983 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21930_ _21938_/A _21938_/B vssd1 vssd1 vccd1 vccd1 _21940_/B sky130_fd_sc_hd__nand2_2
XFILLER_95_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12249__C1 _18945_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21861_ _23271_/Q _21861_/B _21861_/C vssd1 vssd1 vccd1 vccd1 _21861_/Y sky130_fd_sc_hd__nand3b_2
XANTENNA__14738__A _14738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20812_ _20812_/A _20812_/B _20812_/C vssd1 vssd1 vccd1 vccd1 _20836_/A sky130_fd_sc_hd__nand3_1
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21792_ _13520_/A _13492_/A _21791_/Y vssd1 vssd1 vccd1 vccd1 _21792_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_23_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23531_ _23538_/CLK _23531_/D vssd1 vssd1 vccd1 vccd1 _23531_/Q sky130_fd_sc_hd__dfxtp_2
X_20743_ _20743_/A _20747_/C vssd1 vssd1 vccd1 vccd1 _20743_/Y sky130_fd_sc_hd__nand2_1
XFILLER_169_939 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19967__C _19967_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23462_ _23462_/CLK _23474_/Q vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dfxtp_1
XFILLER_184_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20674_ _12640_/A _12637_/X _23454_/Q _12724_/A vssd1 vssd1 vccd1 vccd1 _20674_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_50_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22413_ _22410_/Y _22411_/X _22541_/A _22400_/D vssd1 vssd1 vccd1 vccd1 _22417_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23393_ _23396_/CLK _23393_/D vssd1 vssd1 vccd1 vccd1 _23393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22344_ _22439_/B vssd1 vssd1 vccd1 vccd1 _22344_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16702__A2 _16663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22275_ _22289_/A _22289_/B vssd1 vssd1 vccd1 vccd1 _22288_/A sky130_fd_sc_hd__nand2_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21226_ _21216_/A _21221_/C _21225_/X vssd1 vssd1 vccd1 vccd1 _21228_/C sky130_fd_sc_hd__a21o_1
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21737__C _23325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21157_ _21157_/A _21157_/B _21157_/C _21157_/D vssd1 vssd1 vccd1 vccd1 _21158_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__23593__CLK _23598_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20108_ _20108_/A _20108_/B vssd1 vssd1 vccd1 vccd1 _20111_/D sky130_fd_sc_hd__nand2_1
XFILLER_120_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21088_ _21089_/A _21095_/A _21083_/Y _21087_/Y vssd1 vssd1 vccd1 vccd1 _21088_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_59_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20014__A2 _18373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20039_ _20039_/A _20039_/B vssd1 vssd1 vccd1 vccd1 _20040_/B sky130_fd_sc_hd__nand2_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19504__A _19504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12930_ _12930_/A vssd1 vssd1 vccd1 vccd1 _20773_/A sky130_fd_sc_hd__buf_2
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12861_ _12723_/X _12725_/X _12733_/B _12728_/Y vssd1 vssd1 vccd1 vccd1 _12867_/A
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14648__A _23429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13552__A _13552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14600_ input52/X _14549_/X _14647_/A _14599_/X vssd1 vssd1 vccd1 vccd1 _14600_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11812_ _11853_/A _11807_/X _15682_/B vssd1 vssd1 vccd1 vccd1 _12144_/A sky130_fd_sc_hd__o21ai_2
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15580_ _15580_/A _15580_/B vssd1 vssd1 vccd1 vccd1 _23499_/D sky130_fd_sc_hd__nor2_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12792_ _12792_/A vssd1 vssd1 vccd1 vccd1 _20957_/A sky130_fd_sc_hd__buf_2
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14531_/A vssd1 vssd1 vccd1 vccd1 _14550_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17959__A _17959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11743_/A vssd1 vssd1 vccd1 vccd1 _11746_/A sky130_fd_sc_hd__inv_2
XFILLER_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12168__A _12168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_224 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17250_ _17250_/A vssd1 vssd1 vccd1 vccd1 _17250_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_786 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12007__A2 _12006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14462_ _14461_/A _14461_/C _14472_/B vssd1 vssd1 vccd1 vccd1 _14462_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _23397_/Q vssd1 vssd1 vccd1 vccd1 _11754_/A sky130_fd_sc_hd__clkinv_2
X_16201_ _11822_/A _16319_/A _15797_/A _11848_/X vssd1 vssd1 vccd1 vccd1 _16201_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_186_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13413_ _13407_/Y _13410_/X _22264_/B _22388_/B _13433_/A vssd1 vssd1 vccd1 vccd1
+ _13414_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_155_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17181_ _17181_/A _17181_/B _17181_/C vssd1 vssd1 vccd1 vccd1 _17186_/A sky130_fd_sc_hd__nand3_1
X_14393_ _14393_/A _14393_/B _14433_/D _14407_/D vssd1 vssd1 vccd1 vccd1 _14438_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_183_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16132_ _16132_/A _16132_/B vssd1 vssd1 vccd1 vccd1 _16135_/A sky130_fd_sc_hd__nand2_1
XFILLER_155_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16154__B1 _15971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13344_ _13344_/A _13377_/B _21901_/D _13377_/C vssd1 vssd1 vccd1 vccd1 _13358_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16063_ _16062_/B _16073_/B _16073_/A vssd1 vssd1 vccd1 vccd1 _16063_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13275_ _13498_/B vssd1 vssd1 vccd1 vccd1 _13741_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15901__B1 _16856_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20238__C1 _20237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15014_ _14968_/A _14968_/B _14968_/C _14967_/X vssd1 vssd1 vccd1 vccd1 _15015_/C
+ sky130_fd_sc_hd__a31oi_1
X_12226_ _12532_/A vssd1 vssd1 vccd1 vccd1 _12540_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17103__C1 _19659_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12191__A1 _11935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19822_ _19822_/A _19823_/A _19823_/B vssd1 vssd1 vccd1 vccd1 _19835_/A sky130_fd_sc_hd__nand3_2
X_12157_ _12157_/A _12157_/B _12157_/C vssd1 vssd1 vccd1 vccd1 _12158_/A sky130_fd_sc_hd__nand3_1
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19753_ _19733_/Y _19743_/A _19744_/X vssd1 vssd1 vccd1 vccd1 _19757_/A sky130_fd_sc_hd__a21o_1
X_12088_ _12088_/A vssd1 vssd1 vccd1 vccd1 _12088_/X sky130_fd_sc_hd__clkbuf_4
X_16965_ _17388_/A vssd1 vssd1 vccd1 vccd1 _17899_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_84_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18704_ _18706_/B vssd1 vssd1 vccd1 vccd1 _18892_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15916_ _15916_/A _15916_/B _15916_/C vssd1 vssd1 vccd1 vccd1 _16237_/A sky130_fd_sc_hd__nand3_1
X_19684_ _19684_/A _19684_/B vssd1 vssd1 vccd1 vccd1 _19685_/C sky130_fd_sc_hd__and2_1
X_16896_ _15918_/C _15610_/X _11830_/A _15659_/A vssd1 vssd1 vccd1 vccd1 _16908_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_64_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18635_ _15904_/A _15905_/A _18445_/A _18447_/B vssd1 vssd1 vccd1 vccd1 _18635_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _15920_/A _15678_/Y _15682_/D vssd1 vssd1 vccd1 vccd1 _16311_/A sky130_fd_sc_hd__o21ai_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18566_ _18728_/A _18562_/Y _12522_/C _18559_/X vssd1 vssd1 vccd1 vccd1 _18568_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_18_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _15821_/A _16047_/A vssd1 vssd1 vccd1 vccd1 _16593_/D sky130_fd_sc_hd__nor2_2
XFILLER_80_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17517_ _17522_/B _17522_/C _17522_/D vssd1 vssd1 vccd1 vccd1 _17699_/A sky130_fd_sc_hd__nand3_2
XANTENNA__13181__B _13181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19174__A3 _18461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14729_ _14729_/A _16144_/B vssd1 vssd1 vccd1 vccd1 _14730_/D sky130_fd_sc_hd__nor2_1
XANTENNA__12078__A _20142_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18497_ _18497_/A _18497_/B vssd1 vssd1 vccd1 vccd1 _18499_/B sky130_fd_sc_hd__nand2_2
XFILLER_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17448_ _17269_/X _17248_/Y _17271_/X vssd1 vssd1 vccd1 vccd1 _17453_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17379_ _17379_/A _17379_/B vssd1 vssd1 vccd1 vccd1 _17380_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19331__B1 _19847_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19118_ _12246_/Y _12247_/Y _19363_/C _19363_/D vssd1 vssd1 vccd1 vccd1 _19118_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11710__A _23587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20390_ _20392_/A _20392_/B _23555_/Q vssd1 vssd1 vccd1 vccd1 _20420_/B sky130_fd_sc_hd__a21o_1
XFILLER_173_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19049_ _19046_/Y _19048_/Y _19037_/A vssd1 vssd1 vccd1 vccd1 _19052_/A sky130_fd_sc_hd__o21ai_1
XFILLER_160_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22060_ _13552_/A _22059_/X _22037_/X _22153_/A _22040_/Y vssd1 vssd1 vccd1 vccd1
+ _22061_/B sky130_fd_sc_hd__o221ai_1
XFILLER_126_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19308__B _19308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21011_ _21011_/A _21011_/B _21011_/C vssd1 vssd1 vccd1 vccd1 _21012_/A sky130_fd_sc_hd__nand3_1
XFILLER_102_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16448__A1 _16360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16448__B2 _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12260__B _17149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22962_ _23315_/Q input28/X _22962_/S vssd1 vssd1 vccd1 vccd1 _22963_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21913_ _21913_/A _21913_/B vssd1 vssd1 vccd1 vccd1 _21934_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22893_ _22895_/A _22895_/B vssd1 vssd1 vccd1 vccd1 _23576_/D sky130_fd_sc_hd__nor2_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13372__A _23326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21844_ _21844_/A _21844_/B _21844_/C vssd1 vssd1 vccd1 vccd1 _21844_/X sky130_fd_sc_hd__and3_1
XFILLER_130_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21775_ _13348_/X _21744_/A _21738_/C _22028_/B vssd1 vssd1 vccd1 vccd1 _21777_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20726_ _20862_/A _20707_/Y _20886_/A _20726_/D vssd1 vssd1 vccd1 vccd1 _20862_/B
+ sky130_fd_sc_hd__and4bb_2
XFILLER_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23514_ _23518_/CLK input50/X vssd1 vssd1 vccd1 vccd1 _23514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23445_ _23445_/CLK _23445_/D vssd1 vssd1 vccd1 vccd1 _23445_/Q sky130_fd_sc_hd__dfxtp_1
X_20657_ _20624_/A _20631_/A _20636_/A vssd1 vssd1 vccd1 vccd1 _20667_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12716__A _21039_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23376_ _23443_/CLK _23376_/D vssd1 vssd1 vccd1 vccd1 _23376_/Q sky130_fd_sc_hd__dfxtp_1
X_20588_ _20589_/A _20736_/A _20589_/C vssd1 vssd1 vccd1 vccd1 _20588_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_99 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22327_ _22327_/A _22332_/C vssd1 vssd1 vccd1 vccd1 _22327_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13060_ _13056_/X _12796_/A _13058_/Y _13059_/X vssd1 vssd1 vccd1 vccd1 _13060_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19086__C1 _20317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22258_ _22249_/A _22249_/B _21980_/A vssd1 vssd1 vccd1 vccd1 _22346_/A sky130_fd_sc_hd__o21ai_1
XFILLER_180_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22224__A3 _21988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16439__A1 _11882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ _12011_/A vssd1 vssd1 vccd1 vccd1 _12011_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17636__B1 _17410_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17097__D1 _15807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21209_ _21187_/A _21173_/X _21290_/C _21210_/B vssd1 vssd1 vccd1 vccd1 _21212_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__13547__A _13547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22189_ _13339_/X _22141_/C _23331_/Q _22168_/X _22144_/A vssd1 vssd1 vccd1 vccd1
+ _22191_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_155_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21983__A2 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15762__A _15762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16750_ _16744_/A _16744_/B _16749_/X _16194_/Y vssd1 vssd1 vccd1 vccd1 _16750_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_98_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13962_ _14001_/A _13945_/X _14865_/A _13977_/B vssd1 vssd1 vccd1 vccd1 _14331_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__12476__A2 _19485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22932__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14870__B1 _14621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15701_ _15783_/A _15785_/B vssd1 vssd1 vccd1 vccd1 _15723_/A sky130_fd_sc_hd__nand2_2
XANTENNA__18061__B1 _23530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ _12905_/Y _12909_/Y _12910_/Y _12912_/X vssd1 vssd1 vccd1 vccd1 _13101_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_73_130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16681_ _16679_/Y _16680_/Y _16202_/Y vssd1 vssd1 vccd1 vccd1 _16900_/A sky130_fd_sc_hd__o21ai_4
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13893_ _14430_/A vssd1 vssd1 vccd1 vccd1 _14459_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14378__A _15017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18420_ _23537_/Q _18420_/B _18420_/C vssd1 vssd1 vccd1 vccd1 _18420_/X sky130_fd_sc_hd__and3b_1
XANTENNA__13282__A _23474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15632_ _23429_/Q vssd1 vssd1 vccd1 vccd1 _15713_/B sky130_fd_sc_hd__buf_2
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _12991_/A _12988_/A _12988_/B vssd1 vssd1 vccd1 vccd1 _12911_/B sky130_fd_sc_hd__nand3_1
XFILLER_15_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _18349_/A _18349_/B _18349_/C vssd1 vssd1 vccd1 vccd1 _18355_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__21499__A1 _21548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15563_ _15439_/C _15561_/A _15561_/B vssd1 vssd1 vccd1 vccd1 _15563_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _13138_/C _12776_/B _12775_/C _12775_/D vssd1 vssd1 vccd1 vccd1 _12975_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__16593__A _16593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17302_/A _17302_/B vssd1 vssd1 vccd1 vccd1 _17327_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ input4/X vssd1 vssd1 vccd1 vccd1 _14633_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _18324_/A _18335_/C _18324_/C _18339_/A vssd1 vssd1 vccd1 vccd1 _18284_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11726_/A _11726_/B vssd1 vssd1 vccd1 vccd1 _18805_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16375__B1 _17454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15494_ _15462_/B _15462_/C _15462_/A vssd1 vssd1 vccd1 vccd1 _15494_/X sky130_fd_sc_hd__o21ba_1
XFILLER_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17233_ _17233_/A vssd1 vssd1 vccd1 vccd1 _17766_/C sky130_fd_sc_hd__clkbuf_4
X_14445_ _14446_/A _14446_/B _14446_/C _14465_/C vssd1 vssd1 vccd1 vccd1 _14445_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_35_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11657_ _11823_/A vssd1 vssd1 vccd1 vccd1 _11980_/A sky130_fd_sc_hd__buf_2
XFILLER_11_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22999__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18016__C _18016_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17164_ _17179_/C vssd1 vssd1 vccd1 vccd1 _17170_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14376_ _14371_/Y _14393_/B _14393_/A vssd1 vssd1 vccd1 vccd1 _14377_/C sky130_fd_sc_hd__a21boi_1
XFILLER_31_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11588_ _12497_/A _11960_/B _11593_/C vssd1 vssd1 vccd1 vccd1 _11971_/A sky130_fd_sc_hd__a21o_1
XFILLER_6_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16115_ _17969_/D vssd1 vssd1 vccd1 vccd1 _18169_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13327_ _13269_/X _13313_/X _22392_/C _13320_/X _13561_/A vssd1 vssd1 vccd1 vccd1
+ _13474_/A sky130_fd_sc_hd__o2111ai_4
XANTENNA__15937__A _15937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17095_ _17095_/A _17095_/B vssd1 vssd1 vccd1 vccd1 _17096_/A sky130_fd_sc_hd__nand2_1
XFILLER_142_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16046_ _16194_/A _16315_/A _16045_/Y vssd1 vssd1 vccd1 vccd1 _16046_/Y sky130_fd_sc_hd__o21ai_4
X_13258_ _23320_/Q _23318_/Q vssd1 vssd1 vccd1 vccd1 _13377_/A sky130_fd_sc_hd__nor2_2
XFILLER_124_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17088__D1 _17454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ _16066_/C _11815_/X _12177_/A _11952_/Y _11937_/X vssd1 vssd1 vccd1 vccd1
+ _12211_/C sky130_fd_sc_hd__o32a_1
XFILLER_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18683__A2_N _19491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13189_ _20583_/A _13162_/A _13178_/X _13188_/X vssd1 vssd1 vccd1 vccd1 _13189_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_111_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19805_ _19805_/A vssd1 vssd1 vccd1 vccd1 _20055_/B sky130_fd_sc_hd__buf_2
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13176__B _21182_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17997_ _17999_/B _18085_/B _17996_/X _17869_/Y vssd1 vssd1 vccd1 vccd1 _18022_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__23176__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16850__A1 _15861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15653__A2 _15618_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19736_ _19475_/X _19527_/Y _19571_/Y _19574_/X vssd1 vssd1 vccd1 vccd1 _19736_/Y
+ sky130_fd_sc_hd__o22ai_2
X_16948_ _16948_/A _16948_/B _16948_/C vssd1 vssd1 vccd1 vccd1 _16953_/C sky130_fd_sc_hd__nand3_2
XANTENNA__22518__A4 _22756_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22923__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19667_ _19667_/A _19667_/B _19675_/A _19667_/D vssd1 vssd1 vccd1 vccd1 _19682_/B
+ sky130_fd_sc_hd__nand4_2
X_16879_ _16879_/A _16879_/B _16879_/C vssd1 vssd1 vccd1 vccd1 _16879_/X sky130_fd_sc_hd__and3_1
XFILLER_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11705__A _19363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18618_ _18931_/A _18615_/Y _18617_/X vssd1 vssd1 vccd1 vccd1 _18619_/C sky130_fd_sc_hd__a21o_1
X_19598_ _19598_/A _19598_/B _19598_/C vssd1 vssd1 vccd1 vccd1 _19598_/Y sky130_fd_sc_hd__nand3_1
XFILLER_80_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19001__C1 _19163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18549_ _18519_/Y _18523_/Y _18526_/Y vssd1 vssd1 vccd1 vccd1 _18549_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21560_ _21508_/A _21559_/X _21557_/Y vssd1 vssd1 vccd1 vccd1 _21564_/C sky130_fd_sc_hd__a21o_1
XFILLER_61_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18760__D1 _12260_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16905__A2 _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20511_ _20501_/X _20507_/X _20510_/Y vssd1 vssd1 vccd1 vccd1 _20512_/B sky130_fd_sc_hd__o21ai_2
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21491_ _21561_/A _21561_/B _21491_/C vssd1 vssd1 vccd1 vccd1 _21495_/C sky130_fd_sc_hd__nand3_1
XFILLER_21_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23100__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23230_ _23241_/A vssd1 vssd1 vccd1 vccd1 _23239_/S sky130_fd_sc_hd__clkbuf_2
X_20442_ _20455_/A _20442_/B _20442_/C vssd1 vssd1 vccd1 vccd1 _20444_/A sky130_fd_sc_hd__nor3_1
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21849__A _21852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_912 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23161_ _23403_/Q input20/X _23167_/S vssd1 vssd1 vccd1 vccd1 _23162_/A sky130_fd_sc_hd__mux2_1
X_20373_ _20373_/A _20373_/B vssd1 vssd1 vccd1 vccd1 _20428_/B sky130_fd_sc_hd__nand2_1
XFILLER_161_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23486__D _23498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22112_ _22112_/A _23273_/Q vssd1 vssd1 vccd1 vccd1 _22451_/A sky130_fd_sc_hd__nand2_1
XFILLER_161_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23092_ _23092_/A vssd1 vssd1 vccd1 vccd1 _23372_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17618__B1 _17606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22043_ _22043_/A _22043_/B vssd1 vssd1 vccd1 vccd1 _22061_/C sky130_fd_sc_hd__nand2_1
XFILLER_125_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23167__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22914__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_867 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22945_ _23307_/Q input20/X _22951_/S vssd1 vssd1 vccd1 vccd1 _22946_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11615__A _23397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13407__A1 _13349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22876_ _22876_/A vssd1 vssd1 vccd1 vccd1 _23573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21827_ _21844_/A _21844_/B _21844_/C vssd1 vssd1 vccd1 vccd1 _21827_/Y sky130_fd_sc_hd__nand3_1
XFILLER_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12560_ _23539_/Q _18733_/A vssd1 vssd1 vccd1 vccd1 _12567_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12091__B1 _12088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16357__B1 _18172_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21758_ _13797_/B _13793_/Y _21916_/A _13616_/B vssd1 vssd1 vccd1 vccd1 _21759_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_54_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20709_ _20703_/Y _20705_/X _20708_/X vssd1 vssd1 vccd1 vccd1 _20853_/B sky130_fd_sc_hd__o21ai_4
XFILLER_196_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12491_ _12491_/A _12491_/B vssd1 vssd1 vccd1 vccd1 _12491_/Y sky130_fd_sc_hd__nor2_1
X_21689_ _21689_/A _21688_/Y vssd1 vssd1 vccd1 vccd1 _21690_/A sky130_fd_sc_hd__or2b_1
X_14230_ _14230_/A _14302_/B vssd1 vssd1 vccd1 vccd1 _14826_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23428_ _23428_/CLK _23428_/D vssd1 vssd1 vccd1 vccd1 _23428_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_172_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17306__C1 _17712_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19874__D _19888_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16860__B _16860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14083__D _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14161_ _14162_/B _14360_/A _14167_/A _14167_/D vssd1 vssd1 vccd1 vccd1 _14161_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_125_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23359_ _23359_/CLK _23359_/D vssd1 vssd1 vccd1 vccd1 _23359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13112_ _13113_/A _13113_/B _13113_/C vssd1 vssd1 vccd1 vccd1 _13126_/B sky130_fd_sc_hd__a21o_1
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14092_ _23359_/Q vssd1 vssd1 vccd1 vccd1 _14193_/C sky130_fd_sc_hd__inv_2
XFILLER_4_966 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21197__C _21358_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17920_ _17920_/A _17920_/B _17920_/C vssd1 vssd1 vccd1 vccd1 _18045_/A sky130_fd_sc_hd__nand3_4
XFILLER_140_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22602__B1 _22505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043_ _13041_/X _13042_/X _13032_/X _13038_/Y vssd1 vssd1 vccd1 vccd1 _13048_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15195__C _15195_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17085__A1 _12509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17851_ _17840_/Y _17842_/Y _17848_/X _17850_/Y vssd1 vssd1 vccd1 vccd1 _17880_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21925__C _22510_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16802_ _16802_/A _16802_/B _16816_/B _16802_/D vssd1 vssd1 vccd1 vccd1 _16804_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17782_ _17782_/A _17782_/B _17782_/C vssd1 vssd1 vccd1 vccd1 _17782_/Y sky130_fd_sc_hd__nand3_1
XFILLER_94_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14994_ _13937_/X _14860_/Y _14621_/X vssd1 vssd1 vccd1 vccd1 _14995_/B sky130_fd_sc_hd__o21ai_2
XFILLER_59_480 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22905__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19521_ _19522_/A _19521_/B _19521_/C vssd1 vssd1 vccd1 vccd1 _19526_/A sky130_fd_sc_hd__nand3_1
X_16733_ _16733_/A vssd1 vssd1 vccd1 vccd1 _16744_/A sky130_fd_sc_hd__clkbuf_2
X_13945_ _14863_/D vssd1 vssd1 vccd1 vccd1 _13945_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16045__C1 _17414_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19452_ _19295_/X _19293_/A _19778_/D vssd1 vssd1 vccd1 vccd1 _19453_/B sky130_fd_sc_hd__a21o_1
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16664_ _16458_/A _16928_/A _16662_/Y _16663_/X vssd1 vssd1 vccd1 vccd1 _16939_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_62_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13876_ _13876_/A vssd1 vssd1 vccd1 vccd1 _23559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15938__A3 _17625_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18990__D1 _15928_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18403_ _18403_/A _18403_/B vssd1 vssd1 vccd1 vccd1 _18403_/Y sky130_fd_sc_hd__nand2_1
X_15615_ _15615_/A vssd1 vssd1 vccd1 vccd1 _15631_/B sky130_fd_sc_hd__clkbuf_2
X_19383_ _19573_/A _19573_/B vssd1 vssd1 vccd1 vccd1 _19387_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22756__C _22756_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ _12827_/A vssd1 vssd1 vccd1 vccd1 _20961_/A sky130_fd_sc_hd__clkbuf_2
X_16595_ _11971_/X _11972_/X _16319_/A vssd1 vssd1 vccd1 vccd1 _16595_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22133__A2 _22126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18334_ _20369_/A _17723_/A _17723_/B _20320_/A _18157_/C vssd1 vssd1 vccd1 vccd1
+ _18335_/D sky130_fd_sc_hd__a32o_1
X_15546_ _15558_/A _15546_/B vssd1 vssd1 vccd1 vccd1 _15548_/A sky130_fd_sc_hd__or2_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12872_/A _12874_/B vssd1 vssd1 vccd1 vccd1 _12864_/B sky130_fd_sc_hd__nand2_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12621__A2 _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16899__A1 _11822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18265_ _18265_/A _18265_/B vssd1 vssd1 vccd1 vccd1 _23593_/D sky130_fd_sc_hd__xor2_1
XFILLER_188_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16899__B2 _11848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11709_ _11647_/B _11649_/X _11708_/Y _16619_/A vssd1 vssd1 vccd1 vccd1 _11713_/A
+ sky130_fd_sc_hd__o211ai_4
X_15477_ _15478_/A _15478_/C _15527_/A vssd1 vssd1 vccd1 vccd1 _15479_/A sky130_fd_sc_hd__o21ai_1
X_12689_ _12850_/A vssd1 vssd1 vccd1 vccd1 _12689_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17216_ _17216_/A _17216_/B vssd1 vssd1 vccd1 vccd1 _23584_/D sky130_fd_sc_hd__xnor2_4
XANTENNA__12909__B1 _12902_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14428_ _13978_/A _13978_/B _14181_/A vssd1 vssd1 vccd1 vccd1 _14428_/X sky130_fd_sc_hd__a21o_1
X_18196_ _18122_/Y _18192_/Y _18195_/Y vssd1 vssd1 vccd1 vccd1 _18196_/X sky130_fd_sc_hd__o21a_1
XFILLER_116_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ _16908_/X _17138_/A _17146_/X _17140_/Y vssd1 vssd1 vccd1 vccd1 _17151_/B
+ sky130_fd_sc_hd__o211ai_1
X_14359_ _14251_/Y _14245_/Y _14347_/C vssd1 vssd1 vccd1 vccd1 _14359_/X sky130_fd_sc_hd__o21a_1
XFILLER_183_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20292__B _20295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17078_ _12509_/X _16377_/X _17068_/X _17069_/X _17070_/X vssd1 vssd1 vccd1 vccd1
+ _17079_/D sky130_fd_sc_hd__o221ai_2
XFILLER_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16029_ _16029_/A _16029_/B vssd1 vssd1 vccd1 vccd1 _16089_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19065__A2 _19048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12522__C _12522_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20408__A_N _20407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16498__A _17248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13637__A1 _13495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21554__D _21554_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22012__B _22564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19719_ _19719_/A _19719_/B _19719_/C vssd1 vssd1 vccd1 vccd1 _19719_/Y sky130_fd_sc_hd__nand3_2
X_20991_ _20981_/Y _20985_/X _20986_/Y _20990_/Y vssd1 vssd1 vccd1 vccd1 _20997_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_81_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22730_ _22730_/A _22730_/B vssd1 vssd1 vccd1 vccd1 _22731_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16587__B1 _16275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14047__D1 _14858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16051__A2 _15800_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22661_ _22661_/A _22661_/B _22710_/A vssd1 vssd1 vccd1 vccd1 _22720_/A sky130_fd_sc_hd__nand3_1
XFILLER_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21612_ _21568_/A _21612_/B _21612_/C vssd1 vssd1 vccd1 vccd1 _21630_/B sky130_fd_sc_hd__nand3b_1
XFILLER_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22592_ _22599_/B _22598_/A _22676_/A vssd1 vssd1 vccd1 vccd1 _22594_/B sky130_fd_sc_hd__nand3_1
XFILLER_52_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21543_ _21526_/A _21577_/B _21529_/A vssd1 vssd1 vccd1 vccd1 _21631_/C sky130_fd_sc_hd__a21oi_2
XFILLER_166_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15011__B1 _15371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21474_ _21474_/A _21474_/B vssd1 vssd1 vccd1 vccd1 _21474_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19694__D _19900_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20425_ _20405_/A _20405_/B _20403_/A _20401_/X vssd1 vssd1 vccd1 vccd1 _20430_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_135_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23213_ _16191_/A input10/X _23217_/S vssd1 vssd1 vccd1 vccd1 _23214_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20356_ _20356_/A _20356_/B vssd1 vssd1 vccd1 vccd1 _20356_/Y sky130_fd_sc_hd__nand2_1
XFILLER_161_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23144_ _23144_/A vssd1 vssd1 vccd1 vccd1 _23395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_978 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15865__A2 _16523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23075_ _23097_/A vssd1 vssd1 vccd1 vccd1 _23084_/S sky130_fd_sc_hd__clkbuf_2
X_20287_ _20287_/A _20287_/B _20287_/C vssd1 vssd1 vccd1 vccd1 _20287_/X sky130_fd_sc_hd__and3_1
XFILLER_122_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22026_ _22026_/A vssd1 vssd1 vccd1 vccd1 _22381_/A sky130_fd_sc_hd__buf_2
XFILLER_103_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22060__A1 _13552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22899__A0 _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11991_ _11980_/Y _12121_/B _14646_/A _11838_/A vssd1 vssd1 vccd1 vccd1 _12187_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_17_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19512__A _19868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _13730_/A _13730_/B _13730_/C vssd1 vssd1 vccd1 vccd1 _13730_/Y sky130_fd_sc_hd__nand3_1
XFILLER_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22928_ _22928_/A vssd1 vssd1 vccd1 vccd1 _23299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ _13520_/A _13659_/Y _13660_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Y sky130_fd_sc_hd__o21ai_2
X_22859_ _22859_/A vssd1 vssd1 vccd1 vccd1 _22859_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13560__A _22159_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15400_ _15442_/B _15442_/D _15478_/A vssd1 vssd1 vccd1 vccd1 _15401_/B sky130_fd_sc_hd__a21o_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _20527_/B vssd1 vssd1 vccd1 vccd1 _20528_/B sky130_fd_sc_hd__clkbuf_2
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _16369_/A _16369_/B _16369_/C vssd1 vssd1 vccd1 vccd1 _16380_/Y sky130_fd_sc_hd__a21oi_2
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13800__A1 _13430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13592_ _13755_/C _13755_/B _13755_/A vssd1 vssd1 vccd1 vccd1 _13698_/A sky130_fd_sc_hd__a21o_1
XFILLER_197_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15331_ _15331_/A _15331_/B vssd1 vssd1 vccd1 vccd1 _15332_/B sky130_fd_sc_hd__xnor2_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19531__A3 _17444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12543_ _18437_/D _12542_/B _12542_/A vssd1 vssd1 vccd1 vccd1 _12543_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__14806__D _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23527__CLK _23588_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18050_ _17535_/A _17536_/A _18072_/B _18059_/A vssd1 vssd1 vccd1 vccd1 _18050_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__23076__A0 _15338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15262_ _15262_/A vssd1 vssd1 vccd1 vccd1 _15350_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13159__A3 _21177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ _12474_/A vssd1 vssd1 vccd1 vccd1 _19659_/C sky130_fd_sc_hd__buf_4
XFILLER_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17001_ _17217_/A _17218_/A _16776_/Y _16989_/A _16762_/Y vssd1 vssd1 vccd1 vccd1
+ _17003_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_177_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14213_ _14207_/Y _14212_/X _14800_/A _14934_/A vssd1 vssd1 vccd1 vccd1 _14219_/D
+ sky130_fd_sc_hd__o211ai_2
XFILLER_172_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15193_ _15193_/A _15193_/B _15193_/C vssd1 vssd1 vccd1 vccd1 _15277_/A sky130_fd_sc_hd__nand3_2
XANTENNA__18098__A3 _20210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ _14083_/Y _14084_/X _14101_/Y vssd1 vssd1 vccd1 vccd1 _14222_/A sky130_fd_sc_hd__a21o_1
XFILLER_126_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18952_ _19530_/D _19703_/B _19123_/B _18952_/D vssd1 vssd1 vccd1 vccd1 _18952_/Y
+ sky130_fd_sc_hd__nand4_2
X_14075_ _14075_/A vssd1 vssd1 vccd1 vccd1 _14796_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21936__B _21936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17903_ _17782_/A _17782_/B _17784_/Y vssd1 vssd1 vccd1 vccd1 _17905_/B sky130_fd_sc_hd__a21o_1
X_13026_ _12792_/A _12936_/A _12952_/A _13025_/X _13022_/Y vssd1 vssd1 vccd1 vccd1
+ _13027_/B sky130_fd_sc_hd__o221ai_2
X_18883_ _18782_/X _18786_/Y _18864_/Y vssd1 vssd1 vccd1 vccd1 _18884_/B sky130_fd_sc_hd__o21ai_4
XFILLER_117_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17834_ _17924_/A _17924_/B _17814_/C vssd1 vssd1 vccd1 vccd1 _17834_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_120_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16749__C _16749_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16111__A _17860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18007__B1 _17712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17765_ _17610_/X _17752_/X _17760_/Y _17764_/X vssd1 vssd1 vccd1 vccd1 _17765_/X
+ sky130_fd_sc_hd__o22a_1
X_14977_ _15316_/A _15317_/A vssd1 vssd1 vccd1 vccd1 _14978_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19504_ _19504_/A vssd1 vssd1 vccd1 vccd1 _19504_/X sky130_fd_sc_hd__clkbuf_4
X_16716_ _16700_/A _16956_/A _16712_/B _16712_/A vssd1 vssd1 vccd1 vccd1 _16722_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_13928_ _14173_/B vssd1 vssd1 vccd1 vccd1 _14172_/B sky130_fd_sc_hd__buf_2
X_17696_ _23526_/Q _17529_/B _17533_/B _17695_/Y vssd1 vssd1 vccd1 vccd1 _17951_/A
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19435_ _19259_/A _19259_/B _19259_/C _19431_/A vssd1 vssd1 vccd1 vccd1 _19435_/Y
+ sky130_fd_sc_hd__a31oi_1
X_16647_ _16647_/A _16647_/B _16647_/C vssd1 vssd1 vccd1 vccd1 _16647_/X sky130_fd_sc_hd__and3_1
X_13859_ _13857_/A _13857_/B _13853_/A _13853_/B vssd1 vssd1 vccd1 vccd1 _13861_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_179_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19507__B1 _19649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13470__A _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19366_ _19363_/Y _19540_/A _19365_/Y vssd1 vssd1 vccd1 vccd1 _19371_/A sky130_fd_sc_hd__o21ai_1
X_16578_ _16486_/Y _16492_/Y _16768_/B _17010_/A vssd1 vssd1 vccd1 vccd1 _17009_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15792__A1 _11792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18317_ _18265_/B _18319_/B _18319_/A vssd1 vssd1 vccd1 vccd1 _18318_/B sky130_fd_sc_hd__a21boi_1
XFILLER_188_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15529_ _15478_/A _15528_/C _15528_/B vssd1 vssd1 vccd1 vccd1 _15530_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__21865__A1 _21861_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19297_ _19297_/A _19297_/B _19431_/A vssd1 vssd1 vccd1 vccd1 _19297_/X sky130_fd_sc_hd__and3_1
XFILLER_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1086 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16781__A _18435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23067__A0 _14879_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ _18134_/C _18298_/C _18194_/A _18210_/Y vssd1 vssd1 vccd1 vccd1 _18296_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_124_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18179_ _18179_/A _18179_/B _18227_/B _18179_/D vssd1 vssd1 vccd1 vccd1 _18180_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_156_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20210_ _20210_/A _20265_/B _20210_/C _20210_/D vssd1 vssd1 vccd1 vccd1 _20287_/A
+ sky130_fd_sc_hd__or4_2
X_21190_ _13019_/Y _13014_/Y _20957_/X _13021_/Y vssd1 vssd1 vccd1 vccd1 _21190_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20141_ _20137_/Y _19953_/A _20080_/A _20138_/X _20146_/D vssd1 vssd1 vccd1 vccd1
+ _20141_/X sky130_fd_sc_hd__o311a_1
XFILLER_132_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22042__A1 _22045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20072_ _20068_/Y _20160_/B _20072_/C vssd1 vssd1 vccd1 vccd1 _20172_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__11869__B1 _11741_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13322__A3 _13523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15860__A _16821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20974_ _20974_/A _20974_/B _21101_/A vssd1 vssd1 vccd1 vccd1 _20975_/B sky130_fd_sc_hd__nand3_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22713_ _22713_/A _22756_/B _22713_/C _22713_/D vssd1 vssd1 vccd1 vccd1 _22789_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_14_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22644_ _22644_/A vssd1 vssd1 vccd1 vccd1 _22830_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22575_ _22565_/Y _22573_/Y _22574_/Y vssd1 vssd1 vccd1 vccd1 _22663_/B sky130_fd_sc_hd__o21ai_2
XFILLER_90_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23058__A0 _14588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21526_ _21526_/A _21577_/B vssd1 vssd1 vccd1 vccd1 _21614_/D sky130_fd_sc_hd__nand2_1
XFILLER_139_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21457_ _20906_/X _20907_/X _21493_/C _20908_/X vssd1 vssd1 vccd1 vccd1 _21460_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20408_ _20407_/B _20408_/B vssd1 vssd1 vccd1 vccd1 _20409_/B sky130_fd_sc_hd__and2b_1
XANTENNA__18485__B1 _12149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12190_ _17098_/C vssd1 vssd1 vccd1 vccd1 _19485_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22281__A1 _13465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21388_ _21514_/A _21387_/B _21387_/D _21387_/A vssd1 vssd1 vccd1 vccd1 _21389_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_107_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14361__D _14819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23127_ _23127_/A vssd1 vssd1 vccd1 vccd1 _23387_/D sky130_fd_sc_hd__clkbuf_1
X_20339_ _20339_/A vssd1 vssd1 vccd1 vccd1 _20384_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput55 _14609_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[10] sky130_fd_sc_hd__buf_2
XANTENNA__13849__A1 _22220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput66 _14681_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_150_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput77 _14717_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput88 _23582_/Q vssd1 vssd1 vccd1 vccd1 y[11] sky130_fd_sc_hd__buf_2
X_23058_ _14588_/X input36/X _23062_/S vssd1 vssd1 vccd1 vccd1 _23059_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14900_ _14900_/A _14900_/B _14900_/C vssd1 vssd1 vccd1 vccd1 _14966_/A sky130_fd_sc_hd__nand3_2
X_22009_ _22218_/A _22220_/D _22218_/B vssd1 vssd1 vccd1 vccd1 _22203_/B sky130_fd_sc_hd__and3_1
XFILLER_62_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15880_ _16070_/C _15746_/B _16070_/B vssd1 vssd1 vccd1 vccd1 _15886_/A sky130_fd_sc_hd__a21boi_1
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input23_A wb_dat_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ _14831_/A _14831_/B _14831_/C vssd1 vssd1 vccd1 vccd1 _14831_/Y sky130_fd_sc_hd__nor3_1
Xclkbuf_3_4_0_bq_clk_i clkbuf_3_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_64_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14274__A1 _15231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16866__A _16866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _12323_/X _17303_/A _17888_/A _19862_/A vssd1 vssd1 vccd1 vccd1 _17550_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ _14766_/C _14762_/B _14762_/C vssd1 vssd1 vccd1 vccd1 _14788_/A sky130_fd_sc_hd__nand3b_2
XFILLER_56_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ _11968_/A _11969_/A _12289_/A _11942_/Y vssd1 vssd1 vccd1 vccd1 _12200_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16501_ _16526_/D _16526_/C _16536_/B _16526_/A vssd1 vssd1 vccd1 vccd1 _16501_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _22566_/C vssd1 vssd1 vccd1 vccd1 _22465_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17481_ _17487_/A _17487_/B _17481_/C _17481_/D vssd1 vssd1 vccd1 vccd1 _17482_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_147_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14693_ _14693_/A vssd1 vssd1 vccd1 vccd1 _14693_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13290__A _13523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19220_ _19012_/B _19210_/Y _19013_/X _19201_/Y vssd1 vssd1 vccd1 vccd1 _19220_/Y
+ sky130_fd_sc_hd__o211ai_2
X_16432_ _16426_/Y _16432_/B _16432_/C vssd1 vssd1 vccd1 vccd1 _16757_/C sky130_fd_sc_hd__nand3b_1
X_13644_ _13632_/X _13641_/Y _13643_/Y vssd1 vssd1 vccd1 vccd1 _13645_/C sky130_fd_sc_hd__o21a_1
XFILLER_71_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19151_ _19149_/Y _19150_/X _19052_/B vssd1 vssd1 vccd1 vccd1 _19151_/Y sky130_fd_sc_hd__a21oi_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16389_/A _16322_/B _16323_/A _16499_/A _16462_/B vssd1 vssd1 vccd1 vccd1
+ _16369_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_13_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13756_/B _13575_/B vssd1 vssd1 vccd1 vccd1 _13575_/Y sky130_fd_sc_hd__nor2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18102_ _17766_/B _18100_/A _17766_/C _18101_/B _18101_/D vssd1 vssd1 vccd1 vccd1
+ _18103_/C sky130_fd_sc_hd__a32o_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23049__A0 _14188_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15314_ _15348_/A _15312_/Y _15302_/X _15303_/X vssd1 vssd1 vccd1 vccd1 _15324_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_40_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19082_ _19082_/A _19082_/B _20368_/B _20368_/A vssd1 vssd1 vccd1 vccd1 _19082_/X
+ sky130_fd_sc_hd__or4_4
X_12526_ _12536_/A vssd1 vssd1 vccd1 vccd1 _12528_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16294_ _16294_/A vssd1 vssd1 vccd1 vccd1 _16576_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_185_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18033_ _18033_/A _18033_/B _18033_/C vssd1 vssd1 vccd1 vccd1 _18037_/C sky130_fd_sc_hd__nand3_1
X_15245_ _15245_/A _15245_/B _15245_/C vssd1 vssd1 vccd1 vccd1 _15250_/D sky130_fd_sc_hd__nand3_1
X_12457_ _12451_/Y _18497_/B _12484_/B _12484_/A vssd1 vssd1 vccd1 vccd1 _12490_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_173_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12634__A _12709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output91_A _23265_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15176_ _15095_/X _15170_/Y _15172_/Y _15175_/X vssd1 vssd1 vccd1 vccd1 _15179_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_193_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12388_ _12388_/A _12388_/B _12388_/C vssd1 vssd1 vccd1 vccd1 _12388_/Y sky130_fd_sc_hd__nor3_1
XFILLER_4_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14127_ _14094_/X _14125_/Y _14126_/Y vssd1 vssd1 vccd1 vccd1 _14128_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__15829__A2 _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20822__A2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19984_ _19974_/Y _19977_/Y _19982_/Y vssd1 vssd1 vccd1 vccd1 _19986_/A sky130_fd_sc_hd__o21ai_1
XFILLER_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23584__D _23584_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18935_ _11875_/A _15861_/A _18932_/B vssd1 vssd1 vccd1 vccd1 _18938_/A sky130_fd_sc_hd__o21ai_2
XFILLER_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14058_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14058_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18678__D _18859_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13465__A _13465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ _23296_/Q vssd1 vssd1 vccd1 vccd1 _20494_/D sky130_fd_sc_hd__inv_2
X_18866_ _18863_/A _18863_/B _18865_/Y vssd1 vssd1 vccd1 vccd1 _18866_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17817_ _17817_/A _17817_/B vssd1 vssd1 vccd1 vccd1 _17821_/B sky130_fd_sc_hd__and2_1
XANTENNA__17451__B2 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18797_ _18799_/B _18798_/A _19156_/C vssd1 vssd1 vccd1 vccd1 _18800_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__14265__B2 _15231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17748_ _17566_/X _17575_/X _17583_/B _17571_/Y vssd1 vssd1 vccd1 vccd1 _17751_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_82_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20889__A2 _13121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17679_ _17539_/X _17541_/Y _17832_/C vssd1 vssd1 vccd1 vccd1 _17682_/A sky130_fd_sc_hd__o21ai_1
XFILLER_39_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17754__A2 _17613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11713__A _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19418_ _19416_/Y _19417_/Y _19254_/A _19245_/X vssd1 vssd1 vccd1 vccd1 _19423_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20690_ _20690_/A vssd1 vssd1 vccd1 vccd1 _20718_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19349_ _19230_/B _19189_/X _19179_/Y _19176_/Y vssd1 vssd1 vccd1 vccd1 _19353_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22360_ _22332_/B _22332_/C _22359_/Y vssd1 vssd1 vccd1 vccd1 _22430_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__22663__D _22663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21311_ _21311_/A _21327_/D vssd1 vssd1 vccd1 vccd1 _21311_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22291_ _22288_/Y _22289_/Y _22290_/Y _22166_/Y vssd1 vssd1 vccd1 vccd1 _22291_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_117_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21279__D _21279_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21242_ _21003_/X _21020_/Y _21140_/C vssd1 vssd1 vccd1 vccd1 _21244_/C sky130_fd_sc_hd__o21ai_1
XFILLER_102_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19327__A _19805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21173_ _21187_/B vssd1 vssd1 vccd1 vccd1 _21173_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20124_ _20118_/X _20113_/B _20025_/B _20117_/X vssd1 vssd1 vccd1 vccd1 _20124_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21295__C _21358_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20055_ _20055_/A _20055_/B _20055_/C _20055_/D vssd1 vssd1 vccd1 vccd1 _20056_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11857__A3 _19218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21592__A _21592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12806__A2 _20969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20639__C _20639_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ _20957_/A vssd1 vssd1 vccd1 vccd1 _20957_/X sky130_fd_sc_hd__buf_2
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17745__A2 _18096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _12282_/B _11686_/Y _11689_/Y vssd1 vssd1 vccd1 vccd1 _18849_/C sky130_fd_sc_hd__a21oi_4
X_20888_ _21121_/A _21121_/B _21121_/C _21268_/A vssd1 vssd1 vccd1 vccd1 _20890_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_198_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22627_ _22627_/A _22694_/B vssd1 vssd1 vccd1 vccd1 _22628_/A sky130_fd_sc_hd__and2_1
XFILLER_195_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17310__A _17388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ _13796_/B vssd1 vssd1 vccd1 vccd1 _21767_/A sky130_fd_sc_hd__buf_2
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15749__B _15749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22558_ _22558_/A vssd1 vssd1 vccd1 vccd1 _22700_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12311_ _12311_/A vssd1 vssd1 vccd1 vccd1 _12379_/A sky130_fd_sc_hd__clkbuf_2
X_21509_ _21509_/A _21559_/C vssd1 vssd1 vccd1 vccd1 _21544_/A sky130_fd_sc_hd__xnor2_1
X_13291_ _13712_/A vssd1 vssd1 vccd1 vccd1 _13585_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22489_ _22489_/A _22489_/B _22489_/C vssd1 vssd1 vccd1 vccd1 _22493_/B sky130_fd_sc_hd__nand3_1
XFILLER_170_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15030_ _15077_/A _15030_/B _15030_/C vssd1 vssd1 vccd1 vccd1 _15030_/X sky130_fd_sc_hd__and3_1
XFILLER_142_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12242_ _16225_/A vssd1 vssd1 vccd1 vccd1 _16458_/A sky130_fd_sc_hd__buf_2
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12173_ _12173_/A vssd1 vssd1 vccd1 vccd1 _12173_/X sky130_fd_sc_hd__buf_2
XFILLER_3_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16981_ _17365_/B vssd1 vssd1 vccd1 vccd1 _17369_/A sky130_fd_sc_hd__buf_2
XFILLER_111_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17980__A _17980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18720_ _18914_/A _18914_/B _18914_/C vssd1 vssd1 vccd1 vccd1 _18725_/C sky130_fd_sc_hd__a21bo_1
XFILLER_122_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15932_ _15932_/A vssd1 vssd1 vccd1 vccd1 _16781_/B sky130_fd_sc_hd__buf_2
XFILLER_7_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21765__B1 _13469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11702__C1 _11677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15863_ _15863_/A vssd1 vssd1 vccd1 vccd1 _16523_/C sky130_fd_sc_hd__buf_2
X_18651_ _18973_/A vssd1 vssd1 vccd1 vccd1 _18972_/B sky130_fd_sc_hd__buf_2
XANTENNA__18630__B1 _16360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _19709_/B vssd1 vssd1 vccd1 vccd1 _20055_/C sky130_fd_sc_hd__buf_4
X_14814_ _14814_/A _14814_/B _14814_/C vssd1 vssd1 vccd1 vccd1 _14816_/C sky130_fd_sc_hd__nand3_1
XANTENNA__12258__B1 _12260_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18582_ _18912_/B _18569_/A _12546_/B _18571_/Y vssd1 vssd1 vccd1 vccd1 _18586_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_15794_ _15793_/Y _15650_/Y _15651_/Y vssd1 vssd1 vccd1 vccd1 _15794_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _17533_/A _17533_/B vssd1 vssd1 vccd1 vccd1 _17534_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13732__B _13732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14745_ _23256_/A _16815_/A _14738_/A vssd1 vssd1 vccd1 vccd1 _23268_/D sky130_fd_sc_hd__a21o_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _11966_/A _11966_/B _11915_/A _17642_/A vssd1 vssd1 vccd1 vccd1 _11967_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12629__A _13052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15650__D _16661_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19700__A _19700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17464_ _17276_/B _17258_/Y _17268_/C vssd1 vssd1 vccd1 vccd1 _17471_/B sky130_fd_sc_hd__o21ai_1
X_14676_ _23401_/Q _14672_/X _14647_/X _23433_/Q _14675_/X vssd1 vssd1 vccd1 vccd1
+ _14676_/X sky130_fd_sc_hd__a221o_1
XFILLER_189_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11888_ _11760_/A _11885_/Y _12022_/A vssd1 vssd1 vccd1 vccd1 _12032_/A sky130_fd_sc_hd__o21ai_2
XFILLER_149_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19203_ _19203_/A vssd1 vssd1 vccd1 vccd1 _19203_/X sky130_fd_sc_hd__clkbuf_2
X_16415_ _16517_/C _16415_/B vssd1 vssd1 vccd1 vccd1 _16476_/D sky130_fd_sc_hd__nand2_1
X_13627_ _13627_/A _22269_/C _13816_/A vssd1 vssd1 vccd1 vccd1 _13627_/Y sky130_fd_sc_hd__nand3_2
XFILLER_38_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17395_ _17810_/C _17810_/D _17810_/A vssd1 vssd1 vccd1 vccd1 _17395_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19134_ _19134_/A _19354_/A vssd1 vssd1 vccd1 vccd1 _19409_/C sky130_fd_sc_hd__nand2_1
XFILLER_34_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16346_ _16077_/X _16340_/A _16340_/C vssd1 vssd1 vccd1 vccd1 _16348_/B sky130_fd_sc_hd__a21bo_1
XFILLER_160_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13558_ _13634_/A vssd1 vssd1 vccd1 vccd1 _21988_/A sky130_fd_sc_hd__buf_2
XFILLER_121_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19065_ _19046_/Y _19048_/Y _19052_/B _19037_/A vssd1 vssd1 vccd1 vccd1 _19065_/X
+ sky130_fd_sc_hd__o211a_1
X_12509_ _12509_/A vssd1 vssd1 vccd1 vccd1 _12509_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_121_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16277_ _16108_/A _16108_/B _16108_/C _16581_/C vssd1 vssd1 vccd1 vccd1 _16350_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_146_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13489_ _13400_/Y _13482_/A _13440_/Y vssd1 vssd1 vccd1 vccd1 _13490_/A sky130_fd_sc_hd__o21ai_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18016_ _18161_/C _18016_/B _18016_/C _18016_/D vssd1 vssd1 vccd1 vccd1 _18075_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_173_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15228_ _15228_/A _15228_/B vssd1 vssd1 vccd1 vccd1 _15228_/X sky130_fd_sc_hd__and2_1
XFILLER_160_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20256__B1 _20031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19110__B2 _19082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15159_ _15159_/A _15228_/A vssd1 vssd1 vccd1 vccd1 _15162_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19967_ _19967_/A _19967_/B _19967_/C _19967_/D vssd1 vssd1 vccd1 vccd1 _19985_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_45_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18918_ _18918_/A _18918_/B vssd1 vssd1 vccd1 vccd1 _19443_/A sky130_fd_sc_hd__nand2_1
XFILLER_45_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19898_ _19749_/Y _19750_/Y _19744_/X _19743_/X vssd1 vssd1 vccd1 vccd1 _20017_/C
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_132_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18621__B1 _18617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1166 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18849_ _19017_/A _19364_/A _18849_/C _19017_/D vssd1 vssd1 vccd1 vccd1 _18856_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_68_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12249__B1 _16372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21860_ _22107_/D _22455_/A _22107_/A vssd1 vssd1 vccd1 vccd1 _21861_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__15841__C _16612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19177__A1 _19186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20811_ _20624_/X _20631_/X _20636_/X _20653_/Y vssd1 vssd1 vccd1 vccd1 _20812_/C
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_36_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21791_ _21882_/A _21883_/B _21882_/C vssd1 vssd1 vccd1 vccd1 _21791_/Y sky130_fd_sc_hd__nand3_2
X_23530_ _23558_/CLK _23530_/D vssd1 vssd1 vccd1 vccd1 _23530_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20742_ _21455_/B _20726_/D _20565_/D _20565_/A _20566_/X vssd1 vssd1 vccd1 vccd1
+ _20747_/C sky130_fd_sc_hd__a41o_1
XANTENNA__15199__C1 _14777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23461_ _23559_/CLK _23473_/Q vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20673_ _20673_/A _20673_/B vssd1 vssd1 vccd1 vccd1 _20678_/A sky130_fd_sc_hd__nand2_1
XFILLER_177_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23489__D _23501_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22412_ _22412_/A vssd1 vssd1 vccd1 vccd1 _22541_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23392_ _23395_/CLK _23392_/D vssd1 vssd1 vccd1 vccd1 _23392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22343_ _22246_/A _22246_/B _22439_/B _22439_/A vssd1 vssd1 vccd1 vccd1 _22445_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_164_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22274_ _22474_/C _22269_/Y _22271_/Y _22160_/Y _22183_/Y vssd1 vssd1 vccd1 vccd1
+ _22289_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21225_ _21162_/Y _21165_/X _21166_/Y vssd1 vssd1 vccd1 vccd1 _21225_/X sky130_fd_sc_hd__o21a_1
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21156_ _21014_/X _21002_/Y _20999_/X vssd1 vssd1 vccd1 vccd1 _21158_/B sky130_fd_sc_hd__a21oi_1
XFILLER_144_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_990 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20107_ _20111_/B _20111_/C vssd1 vssd1 vccd1 vccd1 _20110_/A sky130_fd_sc_hd__nand2_1
X_21087_ _21095_/A _21212_/B _21097_/A vssd1 vssd1 vccd1 vccd1 _21087_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12440__C _19193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20038_ _20042_/B _20042_/A _20034_/Y vssd1 vssd1 vccd1 vccd1 _20039_/B sky130_fd_sc_hd__a21o_1
XFILLER_74_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18612__B1 _18080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _12860_/A vssd1 vssd1 vccd1 vccd1 _12900_/A sky130_fd_sc_hd__buf_2
XFILLER_170_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20369__C _20369_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11811_ _15707_/B vssd1 vssd1 vccd1 vccd1 _15682_/B sky130_fd_sc_hd__clkbuf_4
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _13119_/A _13119_/B _20669_/C vssd1 vssd1 vccd1 vccd1 _12815_/C sky130_fd_sc_hd__nand3_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21989_ _21989_/A _21989_/B _21989_/C vssd1 vssd1 vccd1 vccd1 _22086_/A sky130_fd_sc_hd__and3_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14530_ _22968_/D vssd1 vssd1 vccd1 vccd1 _14531_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_732 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _23385_/Q vssd1 vssd1 vccd1 vccd1 _11743_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17959__B _17959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23042__A _23110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14461_ _14461_/A _14472_/B _14461_/C vssd1 vssd1 vccd1 vccd1 _14461_/X sky130_fd_sc_hd__or3_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11618_/C _11606_/X _11828_/B _11672_/Y vssd1 vssd1 vccd1 vccd1 _11851_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_186_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_798 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16200_ _16200_/A vssd1 vssd1 vccd1 vccd1 _16319_/A sky130_fd_sc_hd__buf_2
X_13412_ _22270_/C vssd1 vssd1 vccd1 vccd1 _22388_/B sky130_fd_sc_hd__buf_2
X_17180_ _17121_/A _17335_/A _17178_/Y _17179_/X vssd1 vssd1 vccd1 vccd1 _17181_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_169_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14392_ _14433_/D _14407_/D _14393_/A _14393_/B vssd1 vssd1 vccd1 vccd1 _14438_/A
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__12412__B1 _18997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_984 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23268__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16131_ _16119_/A _16153_/A _15998_/A vssd1 vssd1 vccd1 vccd1 _16132_/B sky130_fd_sc_hd__o21ai_1
XFILLER_195_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17975__A _17975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13343_ _23324_/Q vssd1 vssd1 vccd1 vccd1 _21901_/D sky130_fd_sc_hd__clkinv_2
XFILLER_167_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12184__A _12184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16062_ _16073_/A _16062_/B _16073_/B vssd1 vssd1 vccd1 vccd1 _16062_/Y sky130_fd_sc_hd__nand3_1
XFILLER_154_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13274_ _13366_/B _13732_/B _13228_/X vssd1 vssd1 vccd1 vccd1 _13498_/B sky130_fd_sc_hd__o21ai_2
XFILLER_182_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15013_ _15013_/A _15013_/B _15013_/C _15013_/D vssd1 vssd1 vccd1 vccd1 _15015_/B
+ sky130_fd_sc_hd__nand4_1
X_12225_ _12227_/A _12059_/A _12227_/C vssd1 vssd1 vccd1 vccd1 _12532_/A sky130_fd_sc_hd__a21oi_1
XFILLER_108_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21986__B1 _21992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19821_ _19992_/A _19992_/B _19992_/C vssd1 vssd1 vccd1 vccd1 _19823_/B sky130_fd_sc_hd__nand3_1
XFILLER_97_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12156_ _12143_/Y _12152_/X _12217_/B _12217_/C vssd1 vssd1 vccd1 vccd1 _12157_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_586 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19752_ _19746_/Y _19609_/A _19751_/Y vssd1 vssd1 vccd1 vccd1 _19752_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_96_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12087_ _17610_/A vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__clkbuf_2
X_16964_ _16964_/A _16964_/B _16964_/C vssd1 vssd1 vccd1 vccd1 _16969_/B sky130_fd_sc_hd__nand3_1
XFILLER_111_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18703_ _18528_/Y _18700_/Y _18701_/Y _18702_/Y vssd1 vssd1 vccd1 vccd1 _18706_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA_output54_A _14542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15915_ _15899_/X _15910_/X _15902_/Y _12262_/B _17098_/B vssd1 vssd1 vccd1 vccd1
+ _15916_/C sky130_fd_sc_hd__o2111ai_1
X_19683_ _19503_/X _19647_/Y _19650_/X _19653_/X vssd1 vssd1 vccd1 vccd1 _19684_/A
+ sky130_fd_sc_hd__o211ai_1
X_16895_ _16895_/A _16895_/B _16895_/C vssd1 vssd1 vccd1 vccd1 _17173_/A sky130_fd_sc_hd__nand3_2
XFILLER_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18634_ _18634_/A _18634_/B vssd1 vssd1 vccd1 vccd1 _18830_/B sky130_fd_sc_hd__nand2_2
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _15753_/B _15975_/A _15991_/A _15993_/A _16443_/C vssd1 vssd1 vccd1 vccd1
+ _15943_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16090__B1 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18565_ _18565_/A _18571_/B vssd1 vssd1 vccd1 vccd1 _18568_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _23456_/Q _13181_/B vssd1 vssd1 vccd1 vccd1 _12991_/C sky130_fd_sc_hd__nand2_1
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15777_ _15656_/X _15648_/A _15664_/A vssd1 vssd1 vccd1 vccd1 _16047_/A sky130_fd_sc_hd__a21oi_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17516_ _17385_/Y _17372_/B _17515_/X vssd1 vssd1 vccd1 vccd1 _17537_/A sky130_fd_sc_hd__o21bai_2
X_14728_ _16815_/C vssd1 vssd1 vccd1 vccd1 _16144_/B sky130_fd_sc_hd__inv_2
X_18496_ _18458_/Y _18465_/X _18670_/A _18670_/B vssd1 vssd1 vccd1 vccd1 _18499_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17447_ _17271_/X _17432_/X _17441_/Y _17446_/Y vssd1 vssd1 vccd1 vccd1 _17473_/C
+ sky130_fd_sc_hd__o211ai_4
X_14659_ _15338_/A _14635_/X _14658_/X vssd1 vssd1 vccd1 vccd1 _14659_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20295__B _20295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_707 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20726__D _20726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17378_ _23525_/Q _17379_/A _17379_/B vssd1 vssd1 vccd1 vccd1 _17382_/B sky130_fd_sc_hd__nand3b_1
X_19117_ _18953_/X _18952_/Y _18938_/X vssd1 vssd1 vccd1 vccd1 _19125_/A sky130_fd_sc_hd__a21boi_1
XFILLER_192_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_943 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17885__A _17885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16329_ _16475_/C vssd1 vssd1 vccd1 vccd1 _16422_/B sky130_fd_sc_hd__inv_2
XFILLER_185_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17893__A1 _17644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048_ _18872_/A _18871_/Y _18872_/B _19047_/Y vssd1 vssd1 vccd1 vccd1 _19048_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_160_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12822__A _23455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_851 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19308__C _19308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21010_ _13202_/A _13208_/A _20605_/A _20465_/C vssd1 vssd1 vccd1 vccd1 _21011_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16448__A2 _16447_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22961_ _22961_/A vssd1 vssd1 vccd1 vccd1 _23314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_770 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21912_ _21912_/A vssd1 vssd1 vccd1 vccd1 _21939_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22892_ _22895_/B _22892_/B vssd1 vssd1 vccd1 vccd1 _23575_/D sky130_fd_sc_hd__nor2_4
XFILLER_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21843_ _21844_/A _21844_/B _21844_/C vssd1 vssd1 vccd1 vccd1 _21843_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21774_ _22014_/A vssd1 vssd1 vccd1 vccd1 _22487_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17030__C1 _23428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_776 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23513_ _23518_/CLK input49/X vssd1 vssd1 vccd1 vccd1 _23513_/Q sky130_fd_sc_hd__dfxtp_1
X_20725_ _20725_/A vssd1 vssd1 vccd1 vccd1 _20862_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_184_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23444_ _23444_/CLK _23444_/D vssd1 vssd1 vccd1 vccd1 _23444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20656_ _20512_/B _20655_/X _20518_/X vssd1 vssd1 vccd1 vccd1 _20699_/A sky130_fd_sc_hd__o21ai_2
XFILLER_177_770 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23375_ _23377_/CLK _23375_/D vssd1 vssd1 vccd1 vccd1 _23375_/Q sky130_fd_sc_hd__dfxtp_1
X_20587_ _20577_/Y _20580_/X _21008_/C vssd1 vssd1 vccd1 vccd1 _20597_/A sky130_fd_sc_hd__o21ai_1
XFILLER_99_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22326_ _22332_/A _22332_/B vssd1 vssd1 vccd1 vccd1 _22327_/A sky130_fd_sc_hd__nand2_1
XFILLER_180_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21110__A _21159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22257_ _22253_/Y _22355_/A _22256_/X vssd1 vssd1 vccd1 vccd1 _23563_/D sky130_fd_sc_hd__o21ba_1
XFILLER_151_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _12016_/B _12010_/B vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17636__A1 _16408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21208_ _21208_/A _21208_/B vssd1 vssd1 vccd1 vccd1 _21218_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16439__A2 _11883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22188_ _22553_/A vssd1 vssd1 vccd1 vccd1 _22700_/A sky130_fd_sc_hd__buf_2
XFILLER_120_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21983__A3 _21892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20640__B1 _20495_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21139_ _21123_/X _21129_/Y _21135_/Y vssd1 vssd1 vccd1 vccd1 _21140_/C sky130_fd_sc_hd__o21ai_1
XFILLER_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13961_ _14024_/B vssd1 vssd1 vccd1 vccd1 _14865_/A sky130_fd_sc_hd__buf_2
XFILLER_47_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17035__A _17326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ _12902_/C _12902_/D _12911_/Y vssd1 vssd1 vccd1 vccd1 _12912_/X sky130_fd_sc_hd__a21o_1
XFILLER_4_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15700_ _11764_/A _16315_/A _15699_/Y vssd1 vssd1 vccd1 vccd1 _15785_/B sky130_fd_sc_hd__o21ai_1
XFILLER_111_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16680_ _16032_/A _16033_/A _16677_/C vssd1 vssd1 vccd1 vccd1 _16680_/Y sky130_fd_sc_hd__o21ai_1
X_13892_ _14149_/A vssd1 vssd1 vccd1 vccd1 _14430_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22876__A _22876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16072__B1 _16469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12843_ _12991_/A _12988_/A _12988_/B vssd1 vssd1 vccd1 vccd1 _12911_/A sky130_fd_sc_hd__a21o_1
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15631_ _15712_/C _15631_/B vssd1 vssd1 vccd1 vccd1 _15631_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19888__C _20003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18350_ _18350_/A vssd1 vssd1 vccd1 vccd1 _18355_/A sky130_fd_sc_hd__inv_2
X_15562_ _15528_/A _15559_/B _15561_/B vssd1 vssd1 vccd1 vccd1 _23446_/D sky130_fd_sc_hd__o21bai_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12774_/A _12777_/A vssd1 vssd1 vccd1 vccd1 _12775_/D sky130_fd_sc_hd__nand2_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20396__A _20411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17301_/A _17301_/B vssd1 vssd1 vccd1 vccd1 _17302_/B sky130_fd_sc_hd__nand2_1
X_14513_ _14538_/A vssd1 vssd1 vccd1 vccd1 _14519_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _11916_/A _11838_/A _11798_/A vssd1 vssd1 vccd1 vccd1 _11726_/B sky130_fd_sc_hd__o21ai_1
X_18281_ _18279_/D _18279_/Y _18275_/X _18277_/X vssd1 vssd1 vccd1 vccd1 _18339_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__16375__A1 _16370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15493_ _15493_/A _15493_/B _15493_/C _15508_/C vssd1 vssd1 vccd1 vccd1 _15496_/A
+ sky130_fd_sc_hd__or4_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13189__A1 _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17232_ _17232_/A _17232_/B _17232_/C vssd1 vssd1 vccd1 vccd1 _17397_/A sky130_fd_sc_hd__nand3_2
X_14444_ _14438_/A _14438_/B _14439_/C _14442_/B vssd1 vssd1 vccd1 vccd1 _14446_/C
+ sky130_fd_sc_hd__o211ai_1
X_11656_ _23382_/Q _11656_/B vssd1 vssd1 vccd1 vccd1 _11823_/A sky130_fd_sc_hd__nor2_2
XFILLER_70_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19313__A1 _19304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17163_ _17163_/A _17163_/B _17163_/C vssd1 vssd1 vccd1 vccd1 _17179_/C sky130_fd_sc_hd__nand3_2
XANTENNA__18016__D _18016_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14375_ _15195_/A _14374_/D _15195_/C _14374_/C vssd1 vssd1 vccd1 vccd1 _14393_/A
+ sky130_fd_sc_hd__a31o_1
X_11587_ _11739_/A vssd1 vssd1 vccd1 vccd1 _11960_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_11_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16114_ _17420_/B vssd1 vssd1 vccd1 vccd1 _17969_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_156_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13326_ _13663_/A vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__buf_2
X_17094_ _15634_/C _15618_/X _16591_/B _16591_/A _15652_/A vssd1 vssd1 vccd1 vccd1
+ _17095_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_3_0_bq_clk_i_A clkbuf_3_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16045_ _11799_/X _11801_/X _17414_/C _17414_/D vssd1 vssd1 vccd1 vccd1 _16045_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_108_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ _13257_/A vssd1 vssd1 vccd1 vccd1 _13471_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16114__A _17420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17088__C1 _20049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ _12208_/A vssd1 vssd1 vccd1 vccd1 _16066_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_97_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21955__A _22089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13188_ _13191_/D _13188_/B _13191_/C vssd1 vssd1 vccd1 vccd1 _13188_/X sky130_fd_sc_hd__and3b_1
XFILLER_9_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19804_ _19804_/A vssd1 vssd1 vccd1 vccd1 _20055_/A sky130_fd_sc_hd__buf_2
XFILLER_123_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11911__A2 _11912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19425__A _19534_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _12123_/Y _12129_/Y _12153_/A vssd1 vssd1 vccd1 vccd1 _12139_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_96_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17996_ _17874_/A _17874_/B _17880_/A _17880_/B vssd1 vssd1 vccd1 vccd1 _17996_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__23592__D _23592_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12080__C _18163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19735_ _19735_/A _19735_/B vssd1 vssd1 vccd1 vccd1 _19735_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16850__A2 _16479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16947_ _16945_/Y _16946_/X _16948_/A vssd1 vssd1 vccd1 vccd1 _16953_/B sky130_fd_sc_hd__o21bai_2
XFILLER_42_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19666_ _19675_/A _19667_/D _19667_/A _19667_/B vssd1 vssd1 vccd1 vccd1 _19682_/A
+ sky130_fd_sc_hd__a22o_1
X_16878_ _16843_/Y _16836_/A _16853_/A vssd1 vssd1 vccd1 vccd1 _16878_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_25_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18617_ _16638_/X _16639_/X _11915_/A vssd1 vssd1 vccd1 vccd1 _18617_/X sky130_fd_sc_hd__a21o_2
XFILLER_53_827 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15829_ _11766_/B _16377_/A _15813_/A _15709_/A _15785_/A vssd1 vssd1 vccd1 vccd1
+ _15836_/B sky130_fd_sc_hd__o221ai_4
X_19597_ _19475_/X _19527_/Y _19583_/Y _19595_/Y _19596_/X vssd1 vssd1 vccd1 vccd1
+ _19598_/C sky130_fd_sc_hd__o2111ai_4
XANTENNA__12089__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19160__A _19308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19001__B1 _19308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18548_ _18562_/A _18562_/B vssd1 vssd1 vccd1 vccd1 _18548_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22151__A3 _22145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18479_ _18479_/A vssd1 vssd1 vccd1 vccd1 _19846_/A sky130_fd_sc_hd__buf_2
XFILLER_21_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23583__CLK _23588_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__A _11721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20510_ _20501_/A _20509_/Y _20506_/X vssd1 vssd1 vccd1 vccd1 _20510_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_193_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21490_ _21552_/A _21490_/B vssd1 vssd1 vccd1 vccd1 _21491_/C sky130_fd_sc_hd__nand2_1
XFILLER_119_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12536__B _12536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20441_ _23556_/Q _20419_/B _20440_/Y vssd1 vssd1 vccd1 vccd1 _20442_/C sky130_fd_sc_hd__o21ai_1
XFILLER_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17315__B1 _16908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21849__B _23482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23160_ _23160_/A vssd1 vssd1 vccd1 vccd1 _23402_/D sky130_fd_sc_hd__clkbuf_1
X_20372_ _20371_/B _20215_/B _20215_/C _20371_/A _20371_/D vssd1 vssd1 vccd1 vccd1
+ _20373_/B sky130_fd_sc_hd__a32o_1
XFILLER_118_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22111_ _23273_/Q _22112_/A vssd1 vssd1 vccd1 vccd1 _22113_/A sky130_fd_sc_hd__nor2_1
XFILLER_173_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23091_ _23372_/Q input21/X _23095_/S vssd1 vssd1 vccd1 vccd1 _23092_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22042_ _22045_/A _22045_/B _21913_/B vssd1 vssd1 vccd1 vccd1 _22043_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17094__A2 _15618_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13104__A1 _20464_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22944_ _22944_/A vssd1 vssd1 vccd1 vccd1 _23306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_304 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22875_ _22873_/Y _22875_/B vssd1 vssd1 vccd1 vccd1 _22876_/A sky130_fd_sc_hd__and2b_2
XFILLER_83_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15801__B1 _11741_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22678__A1 _22756_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21826_ _21844_/A _21844_/B _21844_/C vssd1 vssd1 vccd1 vccd1 _21826_/X sky130_fd_sc_hd__a21o_1
XFILLER_145_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21757_ _13793_/B _21906_/A _21753_/B _21750_/Y vssd1 vssd1 vccd1 vccd1 _21759_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_196_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12091__B2 _19082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11631__A _18947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20708_ _20775_/D _20704_/B _20725_/A _20707_/Y vssd1 vssd1 vccd1 vccd1 _20708_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12490_ _12490_/A _12490_/B _18524_/A _18524_/B vssd1 vssd1 vccd1 vccd1 _12494_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__15565__C1 _15559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21688_ _21688_/A _21688_/B _21688_/C _21688_/D vssd1 vssd1 vccd1 vccd1 _21688_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_133_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23427_ _23427_/CLK _23427_/D vssd1 vssd1 vccd1 vccd1 _23427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20639_ _20639_/A _20639_/B _20639_/C _20639_/D vssd1 vssd1 vccd1 vccd1 _20639_/Y
+ sky130_fd_sc_hd__nand4_2
XANTENNA__17306__B1 _17631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20663__B _21065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ _14791_/C _14791_/B _14396_/A _14795_/C vssd1 vssd1 vccd1 vccd1 _14167_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23358_ _23358_/CLK _23358_/D vssd1 vssd1 vccd1 vccd1 _23358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13111_ _13115_/A _13115_/B _21177_/B _13116_/C _13156_/A vssd1 vssd1 vccd1 vccd1
+ _13113_/B sky130_fd_sc_hd__a32o_1
X_22309_ _22045_/B _22040_/B _22051_/X vssd1 vssd1 vccd1 vccd1 _22309_/Y sky130_fd_sc_hd__a21oi_1
X_14091_ _14091_/A vssd1 vssd1 vccd1 vccd1 _15114_/B sky130_fd_sc_hd__buf_2
XFILLER_124_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23289_ _23298_/CLK _23289_/D vssd1 vssd1 vccd1 vccd1 _23289_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21197__D _21295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13042_ _13122_/B _12936_/X _12952_/X _13025_/X _13022_/Y vssd1 vssd1 vccd1 vccd1
+ _13042_/X sky130_fd_sc_hd__o221a_1
XFILLER_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12181__B _12181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17850_ _17855_/A _17853_/A _17982_/B vssd1 vssd1 vccd1 vccd1 _17850_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__17085__A2 _16377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16801_ _16815_/A _16815_/B _16815_/C vssd1 vssd1 vccd1 vccd1 _16802_/D sky130_fd_sc_hd__nor3_1
XFILLER_182_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17781_ _17781_/A _17781_/B vssd1 vssd1 vccd1 vccd1 _17782_/A sky130_fd_sc_hd__nand2_1
XFILLER_120_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14993_ _14879_/C _14864_/Y _15338_/A _15112_/B vssd1 vssd1 vccd1 vccd1 _14995_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19520_ _19494_/X _19335_/B _19328_/Y vssd1 vssd1 vccd1 vccd1 _19521_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__22102__C _22102_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19231__B1 _19048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16732_ _16732_/A _16732_/B _16732_/C vssd1 vssd1 vccd1 vccd1 _16733_/A sky130_fd_sc_hd__nand3_1
XFILLER_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13944_ _23352_/Q vssd1 vssd1 vccd1 vccd1 _13977_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__12854__B1 _20782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16045__B1 _17414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19451_ _19278_/C _19284_/C _19108_/A _19778_/D vssd1 vssd1 vccd1 vccd1 _19451_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16663_ _17142_/A _18461_/A _16194_/A _16194_/B vssd1 vssd1 vccd1 vccd1 _16663_/X
+ sky130_fd_sc_hd__o22a_2
X_13875_ _13875_/A _13875_/B vssd1 vssd1 vccd1 vccd1 _13876_/A sky130_fd_sc_hd__or2_1
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18402_ _23535_/Q vssd1 vssd1 vccd1 vccd1 _18402_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15614_ _15614_/A vssd1 vssd1 vccd1 vccd1 _15712_/C sky130_fd_sc_hd__clkbuf_1
X_12826_ _23454_/Q vssd1 vssd1 vccd1 vccd1 _12827_/A sky130_fd_sc_hd__inv_2
X_19382_ _19380_/X _19381_/X _19361_/A vssd1 vssd1 vccd1 vccd1 _19573_/B sky130_fd_sc_hd__o21ai_2
XFILLER_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16594_ _16382_/A _18675_/A _16601_/C _16601_/B vssd1 vssd1 vccd1 vccd1 _16597_/B
+ sky130_fd_sc_hd__o211ai_1
X_18333_ _20268_/D vssd1 vssd1 vccd1 vccd1 _20320_/A sky130_fd_sc_hd__buf_2
XANTENNA__17212__B _23524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12082__A1 _23256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15545_ _15544_/B _15545_/B vssd1 vssd1 vccd1 vccd1 _15546_/B sky130_fd_sc_hd__and2b_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _12874_/D _12682_/Y _20639_/C _12580_/A _13014_/A vssd1 vssd1 vccd1 vccd1
+ _12872_/A sky130_fd_sc_hd__a41oi_4
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16109__A _16549_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11708_ _12036_/B vssd1 vssd1 vccd1 vccd1 _11708_/Y sky130_fd_sc_hd__clkinv_2
X_18264_ _18264_/A _18264_/B _18264_/C vssd1 vssd1 vccd1 vccd1 _18265_/B sky130_fd_sc_hd__and3_1
X_15476_ _15476_/A _15476_/B vssd1 vssd1 vccd1 vccd1 _15527_/A sky130_fd_sc_hd__xor2_4
X_12688_ _12688_/A _12688_/B vssd1 vssd1 vccd1 vccd1 _12850_/A sky130_fd_sc_hd__nand2_1
X_17215_ _17019_/A _17019_/B _17019_/C _16996_/Y vssd1 vssd1 vccd1 vccd1 _17216_/B
+ sky130_fd_sc_hd__a31o_1
X_14427_ _14430_/D _14876_/B _14430_/A _15094_/C vssd1 vssd1 vccd1 vccd1 _14427_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__23230__A _23241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ _11936_/A vssd1 vssd1 vccd1 vccd1 _16604_/A sky130_fd_sc_hd__clkbuf_4
X_18195_ _18195_/A _18195_/B vssd1 vssd1 vccd1 vccd1 _18195_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__23587__D _23587_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358_ _14358_/A _14358_/B _14358_/C vssd1 vssd1 vccd1 vccd1 _14358_/Y sky130_fd_sc_hd__nand3_1
X_17146_ _11882_/X _11883_/X _16671_/A _16671_/B vssd1 vssd1 vccd1 vccd1 _17146_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13309_ _13308_/Y _22018_/A _23323_/Q vssd1 vssd1 vccd1 vccd1 _13318_/A sky130_fd_sc_hd__a21o_1
XFILLER_155_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17077_ _17077_/A _17077_/B vssd1 vssd1 vccd1 vccd1 _17079_/C sky130_fd_sc_hd__nand2_1
XFILLER_196_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14289_ _14349_/C _14349_/D vssd1 vssd1 vccd1 vccd1 _14358_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16028_ _16028_/A _16028_/B vssd1 vssd1 vccd1 vccd1 _16029_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15087__A1 _15488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16284__B1 _15713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17979_ _17986_/D _17986_/B _17978_/X vssd1 vssd1 vccd1 vccd1 _17994_/A sky130_fd_sc_hd__a21o_1
XFILLER_78_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19718_ _19722_/A _19723_/C vssd1 vssd1 vccd1 vccd1 _19719_/C sky130_fd_sc_hd__nand2_1
XANTENNA__11716__A _19323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20990_ _20990_/A _20994_/A vssd1 vssd1 vccd1 vccd1 _20990_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13634__C _21925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19649_ _19649_/A _19649_/B vssd1 vssd1 vccd1 vccd1 _19649_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21851__C _21858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17784__B1 _17771_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13931__A _23495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22660_ _22585_/Y _22587_/Y _22556_/X vssd1 vssd1 vccd1 vccd1 _22661_/A sky130_fd_sc_hd__a21oi_1
XFILLER_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14062__A2 _14050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21611_ _21611_/A _21611_/B vssd1 vssd1 vccd1 vccd1 _21612_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12073__A1 _11916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22591_ _22591_/A vssd1 vssd1 vccd1 vccd1 _22676_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16019__A _16019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21542_ _21542_/A vssd1 vssd1 vccd1 vccd1 _21542_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_6_0_bq_clk_i clkbuf_4_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _23492_/CLK
+ sky130_fd_sc_hd__clkbuf_8
X_21473_ _21473_/A _21524_/A _21474_/B vssd1 vssd1 vccd1 vccd1 _21482_/B sky130_fd_sc_hd__nand3_1
XFILLER_140_1040 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15562__A2 _15559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23212_ _23212_/A vssd1 vssd1 vccd1 vccd1 _23425_/D sky130_fd_sc_hd__clkbuf_1
X_20424_ _23557_/Q vssd1 vssd1 vccd1 vccd1 _20438_/A sky130_fd_sc_hd__inv_2
XFILLER_119_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22832__A1 _22861_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_648 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23143_ _19156_/B input11/X _23145_/S vssd1 vssd1 vccd1 vccd1 _23144_/A sky130_fd_sc_hd__mux2_1
X_20355_ _20255_/A _20354_/Y _20359_/A _20312_/C vssd1 vssd1 vccd1 vccd1 _20355_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16511__A1 _16510_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23074_ _23074_/A vssd1 vssd1 vccd1 vccd1 _23364_/D sky130_fd_sc_hd__clkbuf_1
X_20286_ _20283_/Y _20235_/X _20327_/A _20282_/Y vssd1 vssd1 vccd1 vccd1 _20287_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_103_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22025_ _22037_/A _22038_/A vssd1 vssd1 vccd1 vccd1 _22025_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__22060__A2 _22059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11626__A _11634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22899__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11990_ _18798_/B vssd1 vssd1 vccd1 vccd1 _14646_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22927_ _23299_/Q input11/X _22929_/S vssd1 vssd1 vccd1 vccd1 _22928_/A sky130_fd_sc_hd__mux2_1
XANTENNA__19512__B _20142_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13660_ _13660_/A _21883_/B _13660_/C vssd1 vssd1 vccd1 vccd1 _13660_/Y sky130_fd_sc_hd__nand3_1
XFILLER_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22858_ _22858_/A vssd1 vssd1 vccd1 vccd1 _22887_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _12601_/B _12601_/A _12875_/C _12608_/X vssd1 vssd1 vccd1 vccd1 _20527_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_71_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21809_ _13830_/Y _13820_/Y _13842_/B _21808_/Y vssd1 vssd1 vccd1 vccd1 _21809_/Y
+ sky130_fd_sc_hd__o22ai_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17032__B _17032_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13591_ _13578_/Y _13587_/Y _13590_/Y vssd1 vssd1 vccd1 vccd1 _13755_/A sky130_fd_sc_hd__a21bo_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22789_ _22789_/A _22789_/B _22789_/C vssd1 vssd1 vccd1 vccd1 _22789_/X sky130_fd_sc_hd__and3_2
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15330_/A _15330_/B vssd1 vssd1 vccd1 vccd1 _15331_/B sky130_fd_sc_hd__xnor2_1
XFILLER_197_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _12542_/A _12542_/B vssd1 vssd1 vccd1 vccd1 _12542_/Y sky130_fd_sc_hd__nand2_1
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15261_ _15262_/A _15419_/A _15263_/A _15156_/X vssd1 vssd1 vccd1 vccd1 _15261_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_40_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12473_ _12473_/A _12473_/B _12473_/C vssd1 vssd1 vccd1 vccd1 _12478_/B sky130_fd_sc_hd__nand3_4
XANTENNA__23076__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14672__A _14693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17000_ _17017_/A _17017_/B _23522_/Q vssd1 vssd1 vccd1 vccd1 _17019_/B sky130_fd_sc_hd__a21o_1
X_14212_ _14764_/A _14764_/B _14097_/A vssd1 vssd1 vccd1 vccd1 _14212_/X sky130_fd_sc_hd__a21o_4
XFILLER_172_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15192_ _15192_/A _15192_/B vssd1 vssd1 vccd1 vccd1 _15193_/C sky130_fd_sc_hd__nand2_1
XFILLER_153_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14143_ _14285_/C _14143_/B vssd1 vssd1 vccd1 vccd1 _14148_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16502__A1 _12346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18951_ _19410_/A _18944_/Y _18950_/Y vssd1 vssd1 vccd1 vccd1 _18951_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14074_ _14178_/A vssd1 vssd1 vccd1 vccd1 _15253_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17902_ _17902_/A _17902_/B vssd1 vssd1 vccd1 vccd1 _17905_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13025_ _13025_/A vssd1 vssd1 vccd1 vccd1 _13025_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18882_ _18882_/A _18882_/B _18774_/A vssd1 vssd1 vccd1 vccd1 _18882_/Y sky130_fd_sc_hd__nor3b_4
X_17833_ _17805_/Y _17708_/Y _17669_/X _17662_/A vssd1 vssd1 vccd1 vccd1 _17924_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18007__A1 _16665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19204__B1 _15882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19703__A _19703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17764_ _17644_/X _17613_/A _17465_/X _17763_/X vssd1 vssd1 vccd1 vccd1 _17764_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14976_ _14976_/A _14983_/A vssd1 vssd1 vccd1 vccd1 _14976_/Y sky130_fd_sc_hd__nor2_1
X_19503_ _20369_/B _20369_/C _19503_/C vssd1 vssd1 vccd1 vccd1 _19503_/X sky130_fd_sc_hd__and3_1
XFILLER_35_602 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16715_ _16722_/A _16950_/A _16713_/Y _16714_/X vssd1 vssd1 vccd1 vccd1 _16715_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13927_ _13927_/A _13939_/A _14124_/A vssd1 vssd1 vccd1 vccd1 _14173_/B sky130_fd_sc_hd__nand3_1
X_17695_ _17528_/A _17528_/B _23526_/Q _17380_/B _23525_/Q vssd1 vssd1 vccd1 vccd1
+ _17695_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_34_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19434_ _19434_/A _19434_/B _19434_/C vssd1 vssd1 vccd1 vccd1 _19434_/X sky130_fd_sc_hd__and3_1
XFILLER_63_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16646_ _16647_/A _16647_/C _16647_/B vssd1 vssd1 vccd1 vccd1 _16646_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13858_ _13853_/A _13853_/B _13857_/X vssd1 vssd1 vccd1 vccd1 _13861_/A sky130_fd_sc_hd__a21o_1
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19507__B2 _18656_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19365_ _19218_/A _15861_/X _19119_/Y vssd1 vssd1 vccd1 vccd1 _19365_/Y sky130_fd_sc_hd__o21ai_2
X_12809_ _12809_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _12810_/B sky130_fd_sc_hd__nand2_1
X_16577_ _16428_/X _16573_/Y _16755_/A _16755_/B vssd1 vssd1 vccd1 vccd1 _17010_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13789_ _13358_/X _21744_/A _21744_/B _13264_/B vssd1 vssd1 vccd1 vccd1 _22064_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__15792__A2 _11792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18316_ _18319_/C _18319_/D vssd1 vssd1 vccd1 vccd1 _18318_/A sky130_fd_sc_hd__nand2_1
XFILLER_194_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15528_ _15528_/A _15528_/B _15528_/C vssd1 vssd1 vccd1 vccd1 _15530_/A sky130_fd_sc_hd__or3_1
XFILLER_175_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19296_ _19261_/C _20320_/A _19261_/A _19263_/X vssd1 vssd1 vccd1 vccd1 _19431_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_163_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21865__A2 _21864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16781__B _16781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1098 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18247_ _18134_/C _18298_/C _18194_/A _18210_/Y _18246_/Y vssd1 vssd1 vccd1 vccd1
+ _18251_/A sky130_fd_sc_hd__o221ai_4
XANTENNA__23067__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15459_ _15459_/A _15459_/B _15353_/C vssd1 vssd1 vccd1 vccd1 _15460_/B sky130_fd_sc_hd__or3b_2
XFILLER_163_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18178_ _18179_/A _18179_/B _18227_/B _18179_/D vssd1 vssd1 vccd1 vccd1 _18180_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17129_ _17298_/B _17126_/X _17127_/Y _17128_/Y vssd1 vssd1 vccd1 vccd1 _17335_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_117_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20140_ _17600_/A _19953_/A _20139_/Y vssd1 vssd1 vccd1 vccd1 _20146_/D sky130_fd_sc_hd__o21ai_2
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20071_ _20071_/A _20160_/A _20071_/C vssd1 vssd1 vccd1 vccd1 _20160_/B sky130_fd_sc_hd__nand3_1
XFILLER_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22042__A2 _22045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11869__A1 _11738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19332__B _19332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20973_ _20973_/A _20973_/B vssd1 vssd1 vccd1 vccd1 _21101_/A sky130_fd_sc_hd__nand2_1
XFILLER_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21553__A1 _21554_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22712_ _22712_/A _22712_/B vssd1 vssd1 vccd1 vccd1 _22713_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22643_ _22643_/A vssd1 vssd1 vccd1 vccd1 _22713_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_638 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13794__A1 _13453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12597__A2 _12601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22574_ _22469_/X _22567_/Y _22468_/A vssd1 vssd1 vccd1 vccd1 _22574_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20494__A _20798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21525_ _21611_/A vssd1 vssd1 vccd1 vccd1 _21577_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23058__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20925__C _21174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21456_ _21377_/B _21378_/C _21455_/Y vssd1 vssd1 vccd1 vccd1 _21456_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12724__B _20966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20407_ _20408_/B _20407_/B vssd1 vssd1 vccd1 vccd1 _20409_/A sky130_fd_sc_hd__and2b_1
XFILLER_135_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_968 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21387_ _21387_/A _21387_/B _21387_/C _21387_/D vssd1 vssd1 vccd1 vccd1 _21389_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__22281__A2 _22059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16496__B1 _16529_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23126_ _12245_/X input34/X _23134_/S vssd1 vssd1 vccd1 vccd1 _23127_/A sky130_fd_sc_hd__mux2_1
X_20338_ _20337_/A _20298_/A _20336_/A _20336_/B vssd1 vssd1 vccd1 vccd1 _20339_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_134_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput56 _14619_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput67 _14684_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_89_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23057_ _23057_/A vssd1 vssd1 vccd1 vccd1 _23356_/D sky130_fd_sc_hd__clkbuf_1
Xoutput78 _14720_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[31] sky130_fd_sc_hd__buf_2
X_20269_ _20271_/A _20269_/B _20269_/C _20269_/D vssd1 vssd1 vccd1 vccd1 _20269_/X
+ sky130_fd_sc_hd__and4_1
Xoutput89 _23263_/Q vssd1 vssd1 vccd1 vccd1 y[1] sky130_fd_sc_hd__buf_2
XFILLER_103_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22008_ _22218_/A _22220_/D _22218_/B vssd1 vssd1 vccd1 vccd1 _22203_/A sky130_fd_sc_hd__a21oi_1
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14830_ _14830_/A vssd1 vssd1 vccd1 vccd1 _14831_/C sky130_fd_sc_hd__inv_2
XANTENNA__12767__A2_N _12770_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20669__A _20669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A wb_dat_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _11971_/X _11972_/X _12089_/A vssd1 vssd1 vccd1 vccd1 _12289_/A sky130_fd_sc_hd__a21o_2
XANTENNA__12285__A1 _12374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ _14756_/Y _14757_/Y _14760_/X vssd1 vssd1 vccd1 vccd1 _14762_/C sky130_fd_sc_hd__o21ai_1
XFILLER_5_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14667__A _14688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _16526_/A _16526_/C _16536_/B _16500_/D vssd1 vssd1 vccd1 vccd1 _16500_/Y
+ sky130_fd_sc_hd__nand4_4
XANTENNA__13571__A _22280_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _13712_/A _22566_/C _22553_/D _13712_/D vssd1 vssd1 vccd1 vccd1 _13727_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17480_ _17480_/A vssd1 vssd1 vccd1 vccd1 _17481_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14692_ _23405_/Q _14672_/X _14677_/X _23437_/Q _14691_/X vssd1 vssd1 vccd1 vccd1
+ _14692_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16431_ _16474_/B _16422_/B _16424_/Y _16425_/Y _16475_/B vssd1 vssd1 vccd1 vccd1
+ _16432_/C sky130_fd_sc_hd__o2111ai_1
X_13643_ _13492_/A _13642_/X _13630_/Y _13632_/A vssd1 vssd1 vccd1 vccd1 _13643_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_72_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12187__A _12187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19150_ _19047_/A _19047_/C _19007_/A _19007_/B vssd1 vssd1 vccd1 vccd1 _19150_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_198_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16362_ _16360_/X _15884_/X _16402_/A vssd1 vssd1 vccd1 vccd1 _16369_/A sky130_fd_sc_hd__o21ai_1
X_13574_ _13712_/A _13527_/X _13573_/D _13573_/A vssd1 vssd1 vccd1 vccd1 _13575_/B
+ sky130_fd_sc_hd__a22oi_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18101_ _18169_/A _18101_/B _18217_/A _18101_/D vssd1 vssd1 vccd1 vccd1 _18103_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_9_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ _12531_/A _12531_/B _12531_/C _12203_/Y _12231_/Y vssd1 vssd1 vccd1 vccd1
+ _12529_/B sky130_fd_sc_hd__a32oi_1
XFILLER_9_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15313_ _15302_/X _15303_/X _15348_/A _15312_/Y vssd1 vssd1 vccd1 vccd1 _15324_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19081_ _18901_/X _19077_/Y _19078_/Y _19079_/Y vssd1 vssd1 vccd1 vccd1 _19087_/A
+ sky130_fd_sc_hd__o211ai_4
X_16293_ _14735_/A _18172_/A _15802_/Y _16292_/X vssd1 vssd1 vccd1 vccd1 _16294_/A
+ sky130_fd_sc_hd__a31o_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__23049__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18032_ _18032_/A _18032_/B vssd1 vssd1 vccd1 vccd1 _18033_/C sky130_fd_sc_hd__nor2_1
XFILLER_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15244_ _15245_/A _15245_/B _15245_/C vssd1 vssd1 vccd1 vccd1 _15250_/C sky130_fd_sc_hd__a21o_1
X_12456_ _12445_/C _18497_/A _12454_/Y _12455_/X vssd1 vssd1 vccd1 vccd1 _12484_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_138_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15175_ _15233_/A _15233_/B _15175_/C vssd1 vssd1 vccd1 vccd1 _15175_/X sky130_fd_sc_hd__and3_1
X_12387_ _12387_/A _12387_/B _12059_/D vssd1 vssd1 vccd1 vccd1 _12388_/C sky130_fd_sc_hd__nor3b_1
XFILLER_153_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14126_ _13927_/A _14091_/A _14070_/X vssd1 vssd1 vccd1 vccd1 _14126_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_output84_A _14597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19983_ _19985_/A _19985_/B _19974_/Y _19977_/Y _19982_/Y vssd1 vssd1 vccd1 vccd1
+ _19987_/B sky130_fd_sc_hd__o221ai_1
XFILLER_114_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18934_ _12246_/Y _12247_/Y _17593_/A _17591_/A _17595_/A vssd1 vssd1 vccd1 vccd1
+ _18934_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__17218__A _17218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ _13933_/Y _13996_/Y _13953_/Y vssd1 vssd1 vccd1 vccd1 _14284_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__12650__A _13121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16122__A _16122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15664__C _15664_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17436__C1 _15974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18779__A2 _18615_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ _12999_/Y _13001_/X _13004_/X _13007_/Y vssd1 vssd1 vccd1 vccd1 _20556_/A
+ sky130_fd_sc_hd__o211ai_4
X_18865_ _18828_/Y _18840_/Y _18875_/C vssd1 vssd1 vccd1 vccd1 _18865_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_121_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17816_ _17821_/A _17832_/D vssd1 vssd1 vccd1 vccd1 _18072_/D sky130_fd_sc_hd__nand2_2
XFILLER_95_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18796_ _18796_/A vssd1 vssd1 vccd1 vccd1 _18796_/X sky130_fd_sc_hd__buf_2
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17747_ _17759_/A _17759_/B _17759_/C vssd1 vssd1 vccd1 vccd1 _17747_/X sky130_fd_sc_hd__and3_2
X_14959_ _15065_/A _15065_/B _14959_/C _15065_/C vssd1 vssd1 vccd1 vccd1 _14960_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_39_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17678_ _17680_/B _17680_/C vssd1 vssd1 vccd1 vccd1 _17832_/C sky130_fd_sc_hd__nand2_1
XANTENNA__20889__A3 _13121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19417_ _19239_/X _19240_/Y _19256_/C _19256_/A vssd1 vssd1 vccd1 vccd1 _19417_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16629_ _16064_/A _16147_/A _16625_/X _16628_/Y vssd1 vssd1 vccd1 vccd1 _16837_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_23_638 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11713__B _11713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16792__A _16792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19348_ _19471_/A _19471_/B _19470_/A vssd1 vssd1 vccd1 vccd1 _19401_/A sky130_fd_sc_hd__nand3_2
XANTENNA_clkbuf_4_13_0_bq_clk_i_A clkbuf_3_6_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_176_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19279_ _19279_/A vssd1 vssd1 vccd1 vccd1 _20120_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21310_ _21319_/A _21319_/B _21308_/Y _21309_/X vssd1 vssd1 vccd1 vccd1 _21327_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20464__D _20464_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22290_ _22290_/A _22290_/B vssd1 vssd1 vccd1 vccd1 _22290_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21241_ _21241_/A _21243_/B _21241_/C vssd1 vssd1 vccd1 vccd1 _21244_/B sky130_fd_sc_hd__nand3_1
XFILLER_85_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21172_ _21172_/A _21453_/D _21438_/A vssd1 vssd1 vccd1 vccd1 _21187_/B sky130_fd_sc_hd__and3_1
XANTENNA__19327__B _19327_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20123_ _20119_/Y _20122_/X _23550_/Q vssd1 vssd1 vccd1 vccd1 _20310_/C sky130_fd_sc_hd__a21o_1
XFILLER_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17690__A2 _18208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20054_ _20054_/A _20054_/B _20054_/C vssd1 vssd1 vccd1 vccd1 _20160_/A sky130_fd_sc_hd__nand3_1
XANTENNA_input8_A wb_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17978__B1 _17644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22971__A0 _21832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater150 _23433_/CLK vssd1 vssd1 vccd1 vccd1 _23401_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__20489__A _21493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20956_ _21497_/A _12981_/C _20953_/X _20955_/X vssd1 vssd1 vccd1 vccd1 _20978_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20887_ _20887_/A _20887_/B vssd1 vssd1 vccd1 vccd1 _21121_/C sky130_fd_sc_hd__nand2_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22626_ _22626_/A _22818_/A _22818_/B vssd1 vssd1 vccd1 vccd1 _22694_/B sky130_fd_sc_hd__nand3_1
XFILLER_139_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22557_ _22641_/B vssd1 vssd1 vccd1 vccd1 _22756_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12310_ _12310_/A vssd1 vssd1 vccd1 vccd1 _12360_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21508_ _21508_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21559_/C sky130_fd_sc_hd__nand2_1
X_13290_ _13523_/A vssd1 vssd1 vccd1 vccd1 _13712_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22488_ _22362_/B _22486_/Y _22647_/A _22477_/Y _22670_/A vssd1 vssd1 vccd1 vccd1
+ _22489_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_166_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11996__D _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20952__A _21295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12241_ _12241_/A vssd1 vssd1 vccd1 vccd1 _16225_/A sky130_fd_sc_hd__clkbuf_2
X_21439_ _21314_/A _21552_/A _21435_/Y _21433_/Y vssd1 vssd1 vccd1 vccd1 _21442_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19655__B1 _19649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12172_ _16122_/A _16122_/B _12256_/A vssd1 vssd1 vccd1 vccd1 _12177_/A sky130_fd_sc_hd__nand3_1
XFILLER_107_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18141__B _23531_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23109_ _23109_/A vssd1 vssd1 vccd1 vccd1 _23380_/D sky130_fd_sc_hd__clkbuf_1
X_16980_ _16969_/X _16975_/Y _16979_/Y vssd1 vssd1 vccd1 vccd1 _17365_/B sky130_fd_sc_hd__o21a_1
XFILLER_111_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19958__A1 _12237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15931_ _15931_/A vssd1 vssd1 vccd1 vccd1 _15932_/A sky130_fd_sc_hd__buf_4
XANTENNA__15781__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18650_ _18798_/A _11608_/A _23394_/Q vssd1 vssd1 vccd1 vccd1 _18973_/A sky130_fd_sc_hd__a21o_1
XANTENNA__18630__A1 _16194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15862_ _15862_/A _15862_/B vssd1 vssd1 vccd1 vccd1 _15863_/A sky130_fd_sc_hd__nor2_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18630__B2 _12103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17601_ _17761_/A vssd1 vssd1 vccd1 vccd1 _19709_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12258__A1 _12308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14813_ _14814_/A _14814_/B _14814_/C vssd1 vssd1 vccd1 vccd1 _14816_/B sky130_fd_sc_hd__a21o_1
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _12563_/Y _19090_/A _18749_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _18588_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_76_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12258__B2 _19503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15793_ _15792_/X _15640_/Y _15772_/X vssd1 vssd1 vccd1 vccd1 _15793_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17532_ _23524_/Q _17531_/X _17382_/B _17382_/D vssd1 vssd1 vccd1 vccd1 _17533_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _23256_/A _12036_/B _14738_/A vssd1 vssd1 vccd1 vccd1 _23267_/D sky130_fd_sc_hd__a21o_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _17626_/A vssd1 vssd1 vccd1 vccd1 _17642_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13732__C _13732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22190__A1 _21902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12629__B _21035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17463_ _17473_/C _17469_/A _17462_/Y vssd1 vssd1 vccd1 vccd1 _17463_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__19700__B _19700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14675_ _23369_/Q _14667_/X _14674_/X vssd1 vssd1 vccd1 vccd1 _14675_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11887_ _11887_/A _18445_/B _11887_/C vssd1 vssd1 vccd1 vccd1 _12022_/A sky130_fd_sc_hd__nand3_2
X_19202_ _19013_/X _19192_/Y _19197_/Y _19201_/Y vssd1 vssd1 vccd1 vccd1 _19202_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_189_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12348__C _12348_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16414_ _16066_/A _16408_/X _15852_/X _16469_/B vssd1 vssd1 vccd1 vccd1 _16415_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_60_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13626_ _13364_/A _13434_/B _13433_/B vssd1 vssd1 vccd1 vccd1 _13626_/Y sky130_fd_sc_hd__a21boi_4
X_17394_ _17140_/B _17305_/Y _17318_/B _17307_/Y vssd1 vssd1 vccd1 vccd1 _17810_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_620 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ _19133_/A _19133_/B vssd1 vssd1 vccd1 vccd1 _19354_/A sky130_fd_sc_hd__nor2_1
XANTENNA__21023__A _23563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16345_ _16347_/A _16347_/B _16347_/C vssd1 vssd1 vccd1 vccd1 _16348_/A sky130_fd_sc_hd__a21o_1
XFILLER_157_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13557_ _13494_/Y _13511_/Y _13507_/Y vssd1 vssd1 vccd1 vccd1 _13557_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19064_ _19058_/A _19057_/D _19060_/B vssd1 vssd1 vccd1 vccd1 _19069_/A sky130_fd_sc_hd__a21o_2
X_12508_ _12508_/A _19543_/B _19811_/A _12508_/D vssd1 vssd1 vccd1 vccd1 _18540_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_185_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13488_ _13479_/X _13482_/Y _13487_/Y _13313_/X vssd1 vssd1 vccd1 vccd1 _13555_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_16276_ _16276_/A vssd1 vssd1 vccd1 vccd1 _16581_/C sky130_fd_sc_hd__inv_2
XFILLER_9_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18015_ _18001_/X _18330_/A _17889_/Y _17896_/C _18014_/Y vssd1 vssd1 vccd1 vccd1
+ _18015_/X sky130_fd_sc_hd__o311a_1
X_15227_ _15120_/D _15164_/B _15154_/X _15156_/X vssd1 vssd1 vccd1 vccd1 _15227_/Y
+ sky130_fd_sc_hd__a211oi_1
X_12439_ _12119_/Y _12122_/Y _12131_/Y vssd1 vssd1 vccd1 vccd1 _12443_/A sky130_fd_sc_hd__a21oi_1
XFILLER_172_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22245__A2 _21981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18332__A _19425_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13391__C1 _13379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15158_ _15154_/X _15156_/X _15120_/D _15164_/B vssd1 vssd1 vccd1 vccd1 _15228_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14109_ _14029_/A _14086_/A _14029_/C _14015_/B vssd1 vssd1 vccd1 vccd1 _15085_/B
+ sky130_fd_sc_hd__a31oi_2
X_19966_ _19966_/A _20062_/C _20133_/B _20061_/A vssd1 vssd1 vccd1 vccd1 _19967_/D
+ sky130_fd_sc_hd__nand4_1
X_15089_ _14097_/X _14976_/A _15488_/C _14987_/Y vssd1 vssd1 vccd1 vccd1 _15089_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_114_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21205__B1 _21207_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18917_ _18726_/Y _18727_/X _18728_/Y _19091_/B _19091_/C vssd1 vssd1 vccd1 vccd1
+ _18918_/B sky130_fd_sc_hd__o311a_1
XANTENNA__16880__B1 _16592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19897_ _19897_/A _19897_/B _19897_/C vssd1 vssd1 vccd1 vccd1 _20017_/B sky130_fd_sc_hd__nand3_1
XFILLER_110_941 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21756__A1 _13430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19163__A _19163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15691__A _15691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18848_ _11935_/A _11846_/A _11669_/A _11936_/A vssd1 vssd1 vccd1 vccd1 _18958_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_95_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12249__A1 _12246_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18779_ _19087_/C _18615_/Y _18620_/Y vssd1 vssd1 vccd1 vccd1 _18882_/A sky130_fd_sc_hd__a21oi_4
XFILLER_83_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20810_ _20817_/A _20810_/B vssd1 vssd1 vccd1 vccd1 _20812_/B sky130_fd_sc_hd__nand2_1
XANTENNA__19177__A2 _18992_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21790_ _13471_/A _13765_/X _13768_/Y vssd1 vssd1 vccd1 vccd1 _21801_/A sky130_fd_sc_hd__o21ai_1
XFILLER_169_1090 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20741_ _20868_/A _20867_/A vssd1 vssd1 vccd1 vccd1 _20743_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15199__B1 _15298_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23460_ _23462_/CLK _23472_/Q vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
X_20672_ _21431_/A _21431_/B _20681_/C _20801_/C _12695_/A vssd1 vssd1 vccd1 vccd1
+ _20672_/X sky130_fd_sc_hd__a32o_1
XANTENNA__18451__A2_N _12441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23130__A0 _12113_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16143__B1_N _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22411_ _22509_/A _22504_/A _22410_/A vssd1 vssd1 vccd1 vccd1 _22411_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23391_ _23391_/CLK _23391_/D vssd1 vssd1 vccd1 vccd1 _23391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16027__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22342_ _22342_/A _22342_/B vssd1 vssd1 vccd1 vccd1 _22439_/A sky130_fd_sc_hd__nor2_1
XFILLER_164_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15866__A _15985_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22273_ _22182_/X _22151_/Y _22192_/Y _22272_/Y vssd1 vssd1 vccd1 vccd1 _22289_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_3_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21224_ _21232_/A _21232_/B _21232_/C _21223_/Y vssd1 vssd1 vccd1 vccd1 _21333_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18860__A1 _18952_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21155_ _20597_/C _20614_/Y _20615_/Y _20616_/Y vssd1 vssd1 vccd1 vccd1 _21158_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_120_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14477__A2 _13985_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20106_ _20106_/A _20106_/B _20106_/C vssd1 vssd1 vccd1 vccd1 _20111_/C sky130_fd_sc_hd__nand3_2
XANTENNA__16871__B1 _16058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21086_ _21057_/A _21057_/B _20941_/Y _20940_/X vssd1 vssd1 vccd1 vccd1 _21097_/A
+ sky130_fd_sc_hd__o2bb2ai_2
X_20037_ _19923_/Y _19789_/Y _19920_/A vssd1 vssd1 vccd1 vccd1 _20039_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__18612__A1 _12167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15977__A2 _16123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20970__A2 _12648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11916_/A _11711_/C _11708_/Y _11809_/Y vssd1 vssd1 vccd1 vccd1 _15707_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _23454_/Q vssd1 vssd1 vccd1 vccd1 _20669_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21988_ _21988_/A _21988_/B _21992_/A _22663_/D vssd1 vssd1 vccd1 vccd1 _21989_/C
+ sky130_fd_sc_hd__nand4_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11741_ _11741_/A _11860_/A vssd1 vssd1 vccd1 vccd1 _11741_/Y sky130_fd_sc_hd__nand2_8
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ _20810_/B _20819_/B _20819_/A vssd1 vssd1 vccd1 vccd1 _20945_/B sky130_fd_sc_hd__a21bo_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14460_ _14456_/B _14456_/C _14181_/X _13964_/Y vssd1 vssd1 vccd1 vccd1 _14461_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11745_/A vssd1 vssd1 vccd1 vccd1 _11672_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_144_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23121__A0 _11743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13411_ _13804_/B vssd1 vssd1 vccd1 vccd1 _22270_/C sky130_fd_sc_hd__buf_2
XFILLER_23_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18679__A1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14391_ _14442_/A vssd1 vssd1 vccd1 vccd1 _14439_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_22609_ _22609_/A _22609_/B vssd1 vssd1 vccd1 vccd1 _22611_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12412__A1 _12410_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23589_ _23598_/CLK _23589_/D vssd1 vssd1 vccd1 vccd1 _23589_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16130_ _16119_/Y _16120_/Y _16125_/Y _16129_/X vssd1 vssd1 vccd1 vccd1 _16174_/C
+ sky130_fd_sc_hd__o22ai_4
X_13342_ _22276_/A _21987_/C _21987_/A _13341_/X _13320_/X vssd1 vssd1 vccd1 vccd1
+ _13474_/B sky130_fd_sc_hd__a32o_1
XFILLER_128_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21778__A _22487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16154__A2 _15884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16061_ _16094_/A _16052_/X _16326_/A vssd1 vssd1 vccd1 vccd1 _16061_/Y sky130_fd_sc_hd__o21ai_1
X_13273_ _13339_/A vssd1 vssd1 vccd1 vccd1 _13366_/B sky130_fd_sc_hd__buf_2
XFILLER_182_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_667 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12224_ _12222_/X _12223_/X _12090_/A vssd1 vssd1 vccd1 vccd1 _12227_/C sky130_fd_sc_hd__a21o_2
X_15012_ _15013_/A _15013_/B _15013_/C _15013_/D vssd1 vssd1 vccd1 vccd1 _15015_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17103__A1 _14599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21986__A1 _22508_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19820_ _19820_/A _19820_/B vssd1 vssd1 vccd1 vccd1 _19992_/C sky130_fd_sc_hd__nand2_1
X_12155_ _12399_/A _12399_/B _12399_/C vssd1 vssd1 vccd1 vccd1 _12217_/C sky130_fd_sc_hd__nand3_1
XFILLER_150_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18851__B2 _17642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19751_ _19747_/Y _19587_/X _19749_/Y _19750_/Y _19743_/X vssd1 vssd1 vccd1 vccd1
+ _19751_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_123_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12086_ _12086_/A vssd1 vssd1 vccd1 vccd1 _17610_/A sky130_fd_sc_hd__buf_2
X_16963_ _16964_/A _16964_/B _16964_/C vssd1 vssd1 vccd1 vccd1 _17202_/A sky130_fd_sc_hd__a21o_1
XFILLER_96_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18702_ _18667_/Y _18672_/Y _18696_/Y _18697_/X vssd1 vssd1 vccd1 vccd1 _18702_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15914_ _11868_/A _15797_/A _15907_/A vssd1 vssd1 vccd1 vccd1 _15916_/B sky130_fd_sc_hd__o21ai_1
X_19682_ _19682_/A _19682_/B _19682_/C vssd1 vssd1 vccd1 vccd1 _19685_/B sky130_fd_sc_hd__nand3_1
X_16894_ _16894_/A _16894_/B _16894_/C _16894_/D vssd1 vssd1 vccd1 vccd1 _16895_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18633_ _18645_/A _18453_/A _18632_/Y vssd1 vssd1 vccd1 vccd1 _18634_/B sky130_fd_sc_hd__o21ai_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _16634_/C vssd1 vssd1 vccd1 vccd1 _16443_/C sky130_fd_sc_hd__buf_2
XFILLER_76_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18564_ _18584_/B _18564_/B _18584_/A vssd1 vssd1 vccd1 vccd1 _18912_/B sky130_fd_sc_hd__nand3_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15776_ _15686_/A _15686_/B _15920_/B _15716_/C vssd1 vssd1 vccd1 vccd1 _15821_/A
+ sky130_fd_sc_hd__a31oi_4
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _12988_/A _12988_/B vssd1 vssd1 vccd1 vccd1 _12991_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _17700_/A _17700_/B vssd1 vssd1 vccd1 vccd1 _17515_/X sky130_fd_sc_hd__and2_1
XFILLER_18_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14727_ _23595_/Q vssd1 vssd1 vccd1 vccd1 _16815_/C sky130_fd_sc_hd__clkbuf_2
X_18495_ _18495_/A _18495_/B _18495_/C vssd1 vssd1 vccd1 vccd1 _18523_/A sky130_fd_sc_hd__nand3_1
X_11939_ _12207_/A vssd1 vssd1 vccd1 vccd1 _15882_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_178_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17446_ _17446_/A _17446_/B vssd1 vssd1 vccd1 vccd1 _17446_/Y sky130_fd_sc_hd__nand2_1
X_14658_ _21852_/A _14636_/X _14642_/X _20902_/B _14657_/X vssd1 vssd1 vccd1 vccd1
+ _14658_/X sky130_fd_sc_hd__a221o_1
XFILLER_162_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13609_ _13793_/A vssd1 vssd1 vccd1 vccd1 _13609_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17377_ _17698_/B _18059_/B _17698_/A vssd1 vssd1 vccd1 vccd1 _17379_/B sky130_fd_sc_hd__a21o_1
X_14589_ _23269_/Q _14551_/X _14587_/X _14588_/X vssd1 vssd1 vccd1 vccd1 _14589_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19331__A2 _19482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19116_ _19116_/A _19116_/B _19116_/C vssd1 vssd1 vccd1 vccd1 _19133_/B sky130_fd_sc_hd__and3_1
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16328_ _16093_/Y _16096_/A _16325_/X _16327_/Y vssd1 vssd1 vccd1 vccd1 _16475_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_185_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_955 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19047_ _19047_/A _19047_/B _19047_/C vssd1 vssd1 vccd1 vccd1 _19047_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__17893__A2 _17763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16259_ _15949_/X _16004_/X _16268_/C _16268_/D vssd1 vssd1 vccd1 vccd1 _16266_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_173_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18997__A _18997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11719__A _11969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18842__A1 _18803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19949_ _19949_/A _20217_/B _20142_/B _19949_/D vssd1 vssd1 vccd1 vccd1 _19951_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12260__D _12260_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13934__A _23495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17406__A _17406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22960_ _23314_/Q input27/X _22962_/S vssd1 vssd1 vccd1 vccd1 _22961_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16605__B1 _16058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21911_ _21911_/A _21911_/B _21911_/C vssd1 vssd1 vccd1 vccd1 _21912_/A sky130_fd_sc_hd__nand3_1
XANTENNA__13419__B1 _13486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22891_ _22891_/A _22891_/B _22891_/C vssd1 vssd1 vccd1 vccd1 _22892_/B sky130_fd_sc_hd__and3_1
XFILLER_56_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21842_ _21842_/A vssd1 vssd1 vccd1 vccd1 _21981_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22154__A1 _13415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21773_ _21771_/X _21772_/X _21755_/X _21760_/X vssd1 vssd1 vccd1 vccd1 _21782_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17030__B1 _17029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20724_ _20724_/A _20724_/B _20724_/C vssd1 vssd1 vccd1 vccd1 _20868_/A sky130_fd_sc_hd__nand3_2
X_23512_ _23518_/CLK input48/X vssd1 vssd1 vccd1 vccd1 _23512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19307__C1 _19163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23443_ _23443_/CLK _23443_/D vssd1 vssd1 vccd1 vccd1 _23443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20655_ _20634_/B _20487_/X _20488_/Y _20490_/Y vssd1 vssd1 vccd1 vccd1 _20655_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23374_ _23377_/CLK _23374_/D vssd1 vssd1 vccd1 vccd1 _23374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20586_ _20583_/Y _20585_/Y _20585_/A vssd1 vssd1 vccd1 vccd1 _21008_/C sky130_fd_sc_hd__o21a_1
XFILLER_109_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18530__B1 _18526_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22325_ _22332_/C _22332_/A _22332_/B vssd1 vssd1 vccd1 vccd1 _22325_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_87_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19086__A1 _12167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22256_ _22451_/A _22451_/B _22452_/A vssd1 vssd1 vccd1 vccd1 _22256_/X sky130_fd_sc_hd__and3_1
XFILLER_151_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21207_ _21267_/C _21270_/A _21207_/C vssd1 vssd1 vccd1 vccd1 _21208_/B sky130_fd_sc_hd__nand3_1
XANTENNA__17097__B1 _15991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17636__A2 _18002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11629__A _12207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22187_ _22187_/A _22187_/B vssd1 vssd1 vccd1 vccd1 _22553_/A sky130_fd_sc_hd__nand2_1
XFILLER_105_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21138_ _20885_/A _20851_/Y _20998_/Y _20996_/X vssd1 vssd1 vccd1 vccd1 _21241_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19515__B _19525_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13844__A _23480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13960_ _14911_/C _15254_/B vssd1 vssd1 vccd1 vccd1 _13960_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21069_ _21064_/X _21069_/B _21069_/C vssd1 vssd1 vccd1 vccd1 _21082_/A sky130_fd_sc_hd__nand3b_2
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12911_ _12911_/A _12911_/B vssd1 vssd1 vccd1 vccd1 _12911_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17035__B _18277_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13563__B _22035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13891_ _14386_/B vssd1 vssd1 vccd1 vccd1 _14149_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15630_ _15712_/A _16187_/B vssd1 vssd1 vccd1 vccd1 _15630_/Y sky130_fd_sc_hd__nand2_2
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16072__B2 _16071_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ _13131_/A _13157_/B _12833_/B _12805_/Y _12809_/B vssd1 vssd1 vccd1 vccd1
+ _12988_/B sky130_fd_sc_hd__a32o_1
XFILLER_73_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19888__D _19888_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23053__A _23110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15561_/A _15561_/B vssd1 vssd1 vccd1 vccd1 _23284_/D sky130_fd_sc_hd__xor2_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12845_/B _12845_/C vssd1 vssd1 vccd1 vccd1 _12777_/A sky130_fd_sc_hd__nand2_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17337_/A _17337_/B vssd1 vssd1 vccd1 vccd1 _17332_/A sky130_fd_sc_hd__nand2_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16593__C _16840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14512_ input2/X vssd1 vssd1 vccd1 vccd1 _14538_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _18275_/X _18277_/X _18279_/D _18279_/Y vssd1 vssd1 vccd1 vccd1 _18324_/C
+ sky130_fd_sc_hd__o211ai_2
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11724_/A vssd1 vssd1 vccd1 vccd1 _11838_/A sky130_fd_sc_hd__inv_2
X_15492_ _15493_/A _15493_/B _15493_/C _15508_/C vssd1 vssd1 vccd1 vccd1 _15497_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_30_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22892__A _22895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17752_/A _12237_/A _17236_/C _17236_/B vssd1 vssd1 vccd1 vccd1 _17232_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17986__A _18172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11655_ _11844_/B vssd1 vssd1 vccd1 vccd1 _12323_/A sky130_fd_sc_hd__buf_2
X_14443_ _14443_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14446_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19313__A2 _19307_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17162_ _17156_/A _17156_/B _17154_/X _17155_/X _17152_/B vssd1 vssd1 vccd1 vccd1
+ _17163_/C sky130_fd_sc_hd__o221ai_1
XFILLER_80_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11586_ _19017_/A vssd1 vssd1 vccd1 vccd1 _19662_/C sky130_fd_sc_hd__clkbuf_4
X_14374_ _15195_/C _15195_/A _14374_/C _14374_/D vssd1 vssd1 vccd1 vccd1 _14393_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18521__B1 _12463_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16113_ _16113_/A vssd1 vssd1 vccd1 vccd1 _17420_/B sky130_fd_sc_hd__clkbuf_4
X_13325_ _13325_/A _13325_/B vssd1 vssd1 vccd1 vccd1 _13663_/A sky130_fd_sc_hd__nand2_1
X_17093_ _15621_/X _15618_/X _17712_/B _17712_/A _16866_/A vssd1 vssd1 vccd1 vccd1
+ _17093_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_116_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ _16044_/A vssd1 vssd1 vccd1 vccd1 _16194_/A sky130_fd_sc_hd__buf_4
X_13256_ _13256_/A vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12207_ _12207_/A vssd1 vssd1 vccd1 vccd1 _12208_/A sky130_fd_sc_hd__clkbuf_2
X_13187_ _13186_/C _13115_/A _13115_/B _13168_/B _13180_/X vssd1 vssd1 vccd1 vccd1
+ _13191_/C sky130_fd_sc_hd__a32o_1
XFILLER_97_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18610__A _18620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19803_ _19803_/A vssd1 vssd1 vccd1 vccd1 _19803_/X sky130_fd_sc_hd__clkbuf_2
X_12138_ _12138_/A _12138_/B _12138_/C vssd1 vssd1 vccd1 vccd1 _12153_/A sky130_fd_sc_hd__nand3_1
XFILLER_97_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19425__B _19900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17995_ _17990_/Y _17991_/X _18085_/A _17994_/Y vssd1 vssd1 vccd1 vccd1 _18085_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__22369__D1 _22548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19734_ _19734_/A _19734_/B vssd1 vssd1 vccd1 vccd1 _19734_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17226__A _19840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ _23592_/Q vssd1 vssd1 vccd1 vccd1 _23258_/B sky130_fd_sc_hd__buf_2
X_16946_ _16934_/X _16936_/Y _16937_/Y _16924_/Y vssd1 vssd1 vccd1 vccd1 _16946_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11885__A1_N _11882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19665_ _19665_/A vssd1 vssd1 vccd1 vccd1 _19667_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16877_ _16849_/X _16850_/X _16836_/A vssd1 vssd1 vccd1 vccd1 _16877_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16063__A1 _16062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18616_ _12090_/A _17980_/A _18931_/A _18615_/Y vssd1 vssd1 vccd1 vccd1 _18619_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _16315_/A vssd1 vssd1 vccd1 vccd1 _16377_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19596_ _19587_/A _19588_/B _19570_/X vssd1 vssd1 vccd1 vccd1 _19596_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18547_ _18554_/A _18554_/B _18547_/C vssd1 vssd1 vccd1 vccd1 _18562_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19001__A1 _16032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15759_ _12174_/A _12173_/A _12175_/A _16160_/A vssd1 vssd1 vccd1 vccd1 _15759_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_79_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21895__B1 _21906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11832__C1 _11743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18478_ _18478_/A vssd1 vssd1 vccd1 vccd1 _18479_/A sky130_fd_sc_hd__buf_2
XFILLER_100_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17429_ _17429_/A _17485_/B _17485_/C vssd1 vssd1 vccd1 vccd1 _17430_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20440_ _20393_/A _20393_/B _20418_/Y _20420_/Y vssd1 vssd1 vccd1 vccd1 _20440_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_158_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17315__A1 _16464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18512__B1 _12460_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20371_ _20371_/A _20371_/B _20371_/C _20371_/D vssd1 vssd1 vccd1 vccd1 _20373_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_107_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22110_ _22617_/A _22108_/X _22109_/Y vssd1 vssd1 vccd1 vccd1 _22112_/A sky130_fd_sc_hd__a21oi_2
XFILLER_161_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23090_ _23090_/A vssd1 vssd1 vccd1 vccd1 _23371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22041_ _22037_/X _22153_/A _22040_/Y vssd1 vssd1 vccd1 vccd1 _22041_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12271__C _19675_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20622__A1 _14615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21881__A _22521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22943_ _23306_/Q input19/X _22951_/S vssd1 vssd1 vccd1 vccd1 _22944_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12863__A1 _12709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17251__B1 _16308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22874_ _22874_/A _22874_/B _22874_/C vssd1 vssd1 vccd1 vccd1 _22875_/B sky130_fd_sc_hd__nand3_1
XFILLER_43_316 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15801__A1 _11738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21825_ _13839_/B _13839_/C _13839_/A _13853_/B _13853_/C vssd1 vssd1 vccd1 vccd1
+ _21844_/C sky130_fd_sc_hd__a32oi_4
XFILLER_197_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22678__A2 _22548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21756_ _13430_/A _22484_/A _21753_/A vssd1 vssd1 vccd1 vccd1 _21759_/A sky130_fd_sc_hd__o21ai_1
XFILLER_145_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16357__A2 _15800_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20707_ _20775_/A _20773_/D _20701_/X _20553_/A vssd1 vssd1 vccd1 vccd1 _20707_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21687_ _21688_/A _21688_/B _21688_/C _21688_/D vssd1 vssd1 vccd1 vccd1 _21689_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_156_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20638_ _23296_/Q _23297_/Q vssd1 vssd1 vccd1 vccd1 _20639_/B sky130_fd_sc_hd__nor2_1
X_23426_ _23427_/CLK _23426_/D vssd1 vssd1 vccd1 vccd1 _23426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17306__A1 _16032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21121__A _21121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16860__D _17066_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23357_ _23359_/CLK _23357_/D vssd1 vssd1 vccd1 vccd1 _23357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20569_ _20579_/A vssd1 vssd1 vccd1 vccd1 _20589_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22308_ _22403_/A _22405_/B _22405_/C vssd1 vssd1 vccd1 vccd1 _22314_/B sky130_fd_sc_hd__and3_1
X_13110_ _21050_/D vssd1 vssd1 vccd1 vccd1 _21177_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_192_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14090_ _14203_/A _14203_/B _14089_/Y vssd1 vssd1 vccd1 vccd1 _14090_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23288_ _23297_/CLK _23288_/D vssd1 vssd1 vccd1 vccd1 _23288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ _13041_/A _13041_/B _20955_/C vssd1 vssd1 vccd1 vccd1 _13041_/X sky130_fd_sc_hd__and3_1
XANTENNA__14540__A1 _14298_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22239_ _22228_/Y _22234_/Y _22238_/X vssd1 vssd1 vccd1 vccd1 _22242_/C sky130_fd_sc_hd__a21bo_1
XFILLER_79_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19464__D1 _19116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14540__B2 _19261_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12181__C _12181_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input46_A x[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16800_ _16800_/A _23258_/B _23593_/Q _16800_/D vssd1 vssd1 vccd1 vccd1 _16816_/B
+ sky130_fd_sc_hd__nor4_2
XANTENNA__16293__A1 _14735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17780_ _17616_/A _17616_/B _17616_/C _17657_/B _17657_/C vssd1 vssd1 vccd1 vccd1
+ _17780_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_8_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14992_ _15000_/A _15000_/B vssd1 vssd1 vccd1 vccd1 _14992_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16731_ _16735_/C _16735_/B _16735_/A vssd1 vssd1 vccd1 vccd1 _16732_/C sky130_fd_sc_hd__nand3b_1
X_13943_ _13994_/A _13994_/B _13942_/X vssd1 vssd1 vccd1 vccd1 _13943_/X sky130_fd_sc_hd__a21o_1
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19231__B2 _19046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16045__A1 _11799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19261__A _19261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19450_ _19447_/A _19447_/B _19295_/X _19293_/A _23545_/Q vssd1 vssd1 vccd1 vccd1
+ _19450_/X sky130_fd_sc_hd__a41o_1
X_16662_ _16662_/A _16662_/B vssd1 vssd1 vccd1 vccd1 _16662_/Y sky130_fd_sc_hd__nor2_1
X_13874_ _23270_/Q _21971_/B vssd1 vssd1 vccd1 vccd1 _13875_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18401_ _18399_/Y _18400_/X _23536_/Q vssd1 vssd1 vccd1 vccd1 _18407_/C sky130_fd_sc_hd__o21ai_2
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15613_ _23414_/Q _23415_/Q _23416_/Q vssd1 vssd1 vccd1 vccd1 _15622_/A sky130_fd_sc_hd__nor3_1
XFILLER_74_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19381_ _19799_/C _19381_/B _19530_/A _19381_/D vssd1 vssd1 vccd1 vccd1 _19381_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_62_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12825_ _12835_/D vssd1 vssd1 vccd1 vccd1 _13157_/B sky130_fd_sc_hd__clkbuf_2
X_16593_ _16593_/A _16860_/C _16840_/A _16593_/D vssd1 vssd1 vccd1 vccd1 _16601_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA__22669__A2 _22476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18332_ _19425_/C vssd1 vssd1 vccd1 vccd1 _20369_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11822__A _11822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15544_ _15545_/B _15544_/B vssd1 vssd1 vccd1 vccd1 _15558_/A sky130_fd_sc_hd__and2b_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_844 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12756_/A _12756_/B vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__nand2_2
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _18263_/A _18263_/B vssd1 vssd1 vccd1 vccd1 _18264_/C sky130_fd_sc_hd__nand2_1
X_11707_ _23588_/Q vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__buf_2
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15475_ _15475_/A _15475_/B vssd1 vssd1 vccd1 vccd1 _15476_/B sky130_fd_sc_hd__nand2_2
XFILLER_147_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12687_ _12687_/A _12687_/B vssd1 vssd1 vccd1 vccd1 _20670_/C sky130_fd_sc_hd__nand2_1
X_17214_ _17381_/C _17382_/A vssd1 vssd1 vccd1 vccd1 _17216_/A sky130_fd_sc_hd__nand2_2
XFILLER_147_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14426_ _14886_/B vssd1 vssd1 vccd1 vccd1 _15094_/C sky130_fd_sc_hd__clkbuf_2
X_18194_ _18194_/A vssd1 vssd1 vccd1 vccd1 _18195_/B sky130_fd_sc_hd__inv_2
X_11638_ _16591_/A _16591_/B vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__nand2_4
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22127__A _22365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18324__B _18335_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17145_ _17151_/A _17145_/B _17145_/C vssd1 vssd1 vccd1 vccd1 _17152_/A sky130_fd_sc_hd__nand3b_1
XFILLER_196_1020 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17848__A2 _20133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16505__C1 _19653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14357_ _14354_/Y _14355_/X _14403_/B vssd1 vssd1 vccd1 vccd1 _14357_/X sky130_fd_sc_hd__o21a_1
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11569_ _23584_/Q _23583_/Q vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__nor2_1
XFILLER_143_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13308_ _13377_/A _13377_/B _13377_/D vssd1 vssd1 vccd1 vccd1 _13308_/Y sky130_fd_sc_hd__nand3_2
XFILLER_143_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17076_ _17073_/Y _16843_/Y _17075_/Y vssd1 vssd1 vccd1 vccd1 _17221_/B sky130_fd_sc_hd__o21ai_1
XFILLER_157_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14288_ _14284_/A _14284_/B _14285_/B _14285_/C vssd1 vssd1 vccd1 vccd1 _14292_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16027_ _16027_/A _16027_/B _16308_/C _16027_/D vssd1 vssd1 vccd1 vccd1 _16028_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_171_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13239_ _13299_/A _13563_/C _13563_/A _21878_/A vssd1 vssd1 vccd1 vccd1 _13247_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20604__A1 _13202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15087__A2 _15231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11750__D1 _11749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17978_ _16638_/X _16639_/X _17644_/X vssd1 vssd1 vccd1 vccd1 _17978_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19717_ _19717_/A _19717_/B vssd1 vssd1 vccd1 vccd1 _19723_/C sky130_fd_sc_hd__nor2_2
X_16929_ _17304_/A _16662_/B _16917_/X _16923_/A vssd1 vssd1 vccd1 vccd1 _16936_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_66_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16036__A1 _16447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19648_ _19648_/A _19651_/A _19652_/A vssd1 vssd1 vccd1 vccd1 _19656_/B sky130_fd_sc_hd__nand3_2
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_619 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19579_ _19576_/Y _19577_/X _19578_/Y vssd1 vssd1 vccd1 vccd1 _19734_/B sky130_fd_sc_hd__o21ai_2
XFILLER_168_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21610_ _21521_/B _21521_/A _21568_/B vssd1 vssd1 vccd1 vccd1 _21611_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14062__A3 _14061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22590_ _22589_/B _22589_/C _22589_/A vssd1 vssd1 vccd1 vccd1 _22591_/A sky130_fd_sc_hd__a21o_1
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21541_ _21541_/A _23569_/Q _21541_/C vssd1 vssd1 vccd1 vccd1 _21627_/B sky130_fd_sc_hd__nand3_1
XFILLER_139_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21472_ _21472_/A _21472_/B vssd1 vssd1 vccd1 vccd1 _21474_/B sky130_fd_sc_hd__or2_1
XFILLER_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15858__B _15858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23211_ _15921_/C input9/X _23217_/S vssd1 vssd1 vccd1 vccd1 _23212_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20423_ _20423_/A _20423_/B vssd1 vssd1 vccd1 vccd1 _23536_/D sky130_fd_sc_hd__nand2_1
XFILLER_105_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13659__A _13659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1074 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23142_ _23142_/A vssd1 vssd1 vccd1 vccd1 _23394_/D sky130_fd_sc_hd__clkbuf_1
X_20354_ _20354_/A _20354_/B vssd1 vssd1 vccd1 vccd1 _20354_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16511__A2 _18017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_906 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23073_ _23364_/Q input12/X _23073_/S vssd1 vssd1 vccd1 vccd1 _23074_/A sky130_fd_sc_hd__mux2_1
X_20285_ _20285_/A vssd1 vssd1 vccd1 vccd1 _20327_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17792__C _17792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22024_ _22026_/A _22039_/B _22024_/C vssd1 vssd1 vccd1 vccd1 _22038_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15078__A2 _14068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11907__A _11969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22926_ _22926_/A vssd1 vssd1 vccd1 vccd1 _23298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19512__C _19512_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14589__A1 _23269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14589__B2 _14588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22857_ _22850_/Y _22847_/Y _22856_/C _22852_/Y vssd1 vssd1 vccd1 vccd1 _22874_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11642__A _23583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ _20528_/A vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__clkbuf_2
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21808_ _21807_/Y _13829_/Y _13834_/B vssd1 vssd1 vccd1 vccd1 _21808_/Y sky130_fd_sc_hd__a21boi_1
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13590_ _13577_/Y _13590_/B _13590_/C vssd1 vssd1 vccd1 vccd1 _13590_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22788_ _22710_/A _22709_/A _22800_/C _22718_/X _22766_/Y vssd1 vssd1 vccd1 vccd1
+ _22788_/X sky130_fd_sc_hd__o311a_2
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _18437_/D vssd1 vssd1 vccd1 vccd1 _12541_/Y sky130_fd_sc_hd__inv_2
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21739_ _21739_/A _21745_/B vssd1 vssd1 vccd1 vccd1 _21740_/B sky130_fd_sc_hd__and2_1
XFILLER_197_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15260_ _14212_/X _15166_/Y _15259_/C _15259_/A vssd1 vssd1 vccd1 vccd1 _15260_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12472_ _12104_/X _12107_/A _12151_/Y _12093_/X vssd1 vssd1 vccd1 vccd1 _12473_/C
+ sky130_fd_sc_hd__o2bb2ai_4
X_14211_ _14879_/A _14878_/A vssd1 vssd1 vccd1 vccd1 _14764_/B sky130_fd_sc_hd__nand2_1
X_23409_ _23409_/CLK _23409_/D vssd1 vssd1 vccd1 vccd1 _23409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15191_ _15191_/A _15191_/B vssd1 vssd1 vccd1 vccd1 _15192_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14142_ _14056_/A _14056_/B _14056_/C _14284_/B _14284_/A vssd1 vssd1 vccd1 vccd1
+ _14143_/B sky130_fd_sc_hd__a32o_1
XFILLER_153_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16502__A2 _15974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18950_ _18950_/A _18950_/B vssd1 vssd1 vccd1 vccd1 _18950_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14073_ _14752_/C vssd1 vssd1 vccd1 vccd1 _14178_/A sky130_fd_sc_hd__buf_2
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17901_ _17901_/A _17901_/B vssd1 vssd1 vccd1 vccd1 _17902_/B sky130_fd_sc_hd__nor2_1
XFILLER_152_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13024_ _13041_/A _20805_/C _20669_/A vssd1 vssd1 vccd1 vccd1 _13027_/A sky130_fd_sc_hd__nand3_1
X_18881_ _18773_/C _18773_/D _18880_/Y vssd1 vssd1 vccd1 vccd1 _18882_/B sky130_fd_sc_hd__a21oi_4
XFILLER_79_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17832_ _17832_/A _17832_/B _17832_/C _17832_/D vssd1 vssd1 vccd1 vccd1 _17928_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_39_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14277__B1 _15225_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17763_ _17763_/A vssd1 vssd1 vccd1 vccd1 _17763_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18007__A2 _17029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19204__A1 _19196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19204__B2 _19803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19703__B _19703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14975_ _15316_/A _15317_/A _14975_/C vssd1 vssd1 vccd1 vccd1 _14983_/A sky130_fd_sc_hd__nand3_1
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19502_ _19502_/A vssd1 vssd1 vccd1 vccd1 _20369_/B sky130_fd_sc_hd__clkbuf_2
X_16714_ _16957_/A _16956_/A _16956_/B vssd1 vssd1 vccd1 vccd1 _16714_/X sky130_fd_sc_hd__and3_1
XANTENNA__18412__C1 _18376_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13926_ _14172_/A vssd1 vssd1 vccd1 vccd1 _15353_/A sky130_fd_sc_hd__clkbuf_2
X_17694_ _17684_/X _17689_/X _17693_/Y vssd1 vssd1 vccd1 vccd1 _17951_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15232__A2_N _15054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19433_ _19428_/Y _19616_/B _19430_/Y _19432_/Y vssd1 vssd1 vccd1 vccd1 _19433_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16645_ _16645_/A _16655_/D _16655_/A vssd1 vssd1 vccd1 vccd1 _16645_/Y sky130_fd_sc_hd__nand3_1
X_13857_ _13857_/A _13857_/B vssd1 vssd1 vccd1 vccd1 _13857_/X sky130_fd_sc_hd__or2_1
XANTENNA__15777__B1 _15664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19364_ _19364_/A _19364_/B _19364_/C vssd1 vssd1 vccd1 vccd1 _19540_/A sky130_fd_sc_hd__nand3_2
X_12808_ _13166_/A _20969_/A vssd1 vssd1 vccd1 vccd1 _12809_/B sky130_fd_sc_hd__nor2_1
X_16576_ _16576_/A _16576_/B vssd1 vssd1 vccd1 vccd1 _16755_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13788_ _23328_/Q vssd1 vssd1 vccd1 vccd1 _21744_/B sky130_fd_sc_hd__clkbuf_4
X_18315_ _18315_/A _23534_/Q _18315_/C vssd1 vssd1 vccd1 vccd1 _18319_/D sky130_fd_sc_hd__nand3_1
XFILLER_163_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1044 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23241__A _23241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15529__B1 _15528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15527_ _15527_/A _15527_/B _15478_/C vssd1 vssd1 vccd1 vccd1 _15528_/C sky130_fd_sc_hd__nor3b_1
X_19295_ _19295_/A vssd1 vssd1 vccd1 vccd1 _19295_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15959__A _23594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12739_ _12846_/A vssd1 vssd1 vccd1 vccd1 _12901_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14863__A _14863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18246_ _18241_/Y _18243_/Y _18293_/A _18267_/A vssd1 vssd1 vccd1 vccd1 _18246_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_124_1047 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ _15458_/A _15458_/B vssd1 vssd1 vccd1 vccd1 _15460_/A sky130_fd_sc_hd__nand2_1
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14409_ _14354_/Y _14355_/X _14403_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14410_/D
+ sky130_fd_sc_hd__o211ai_1
X_18177_ _18165_/A _18165_/B _18176_/B _18227_/A vssd1 vssd1 vccd1 vccd1 _18179_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_163_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15389_ _15385_/Y _15403_/A _15299_/B _15388_/X vssd1 vssd1 vccd1 vccd1 _15435_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_156_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17128_ _17125_/A _17298_/A _17117_/Y _17118_/X vssd1 vssd1 vccd1 vccd1 _17128_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_117_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17059_ _17048_/Y _17052_/X _17053_/Y _17058_/Y vssd1 vssd1 vccd1 vccd1 _17089_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_144_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22578__A1 _13547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_831 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20070_ _19955_/X _20043_/Y _20068_/Y _20069_/X vssd1 vssd1 vccd1 vccd1 _20070_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11869__A2 _11740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20053__A2 _18211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1056 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14807__A2 _15019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17414__A _17414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20972_ _20959_/X _20960_/Y _21431_/C _20963_/Y _12980_/A vssd1 vssd1 vccd1 vccd1
+ _20974_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__15860__C _15860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21553__A2 _21358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22711_ _22656_/B _22700_/A _22656_/A _22656_/D _22709_/Y vssd1 vssd1 vccd1 vccd1
+ _22717_/B sky130_fd_sc_hd__a41o_1
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18757__A2_N _18755_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22642_ _22649_/C _22642_/B _22642_/C vssd1 vssd1 vccd1 vccd1 _22643_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__17509__A1 _16480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20775__A _20775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15869__A _19703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22573_ _22573_/A vssd1 vssd1 vccd1 vccd1 _22573_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21524_ _21524_/A _21524_/B _21524_/C vssd1 vssd1 vccd1 vccd1 _21611_/A sky130_fd_sc_hd__nand3_2
XFILLER_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23301__D _23301_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23446__CLK _23492_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13389__A _22145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21455_ _21455_/A _21455_/B vssd1 vssd1 vccd1 vccd1 _21455_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19131__B1 _19391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20406_ _20379_/A _20379_/B _20401_/B _20376_/B vssd1 vssd1 vccd1 vccd1 _20407_/B
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12724__C _20781_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21386_ _21386_/A _21386_/B _21386_/C _21490_/B vssd1 vssd1 vccd1 vccd1 _21387_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16496__A1 _12149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20337_ _20337_/A _20343_/A _20337_/C vssd1 vssd1 vccd1 vccd1 _20337_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__16496__B2 _16549_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23125_ _23182_/S vssd1 vssd1 vccd1 vccd1 _23134_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_162_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23596__CLK _23598_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput57 _14629_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[12] sky130_fd_sc_hd__buf_2
X_23056_ _14031_/X input35/X _23062_/S vssd1 vssd1 vccd1 vccd1 _23057_/A sky130_fd_sc_hd__mux2_1
X_20268_ _20268_/A _20268_/B _20268_/C _20268_/D vssd1 vssd1 vccd1 vccd1 _20274_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_103_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput68 _14687_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput79 _14567_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_89_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22007_ _21997_/X _21892_/X _21881_/Y _22006_/X vssd1 vssd1 vccd1 vccd1 _22218_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_89_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19804__A _19804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20199_ _23551_/Q _20199_/B _20199_/C vssd1 vssd1 vccd1 vccd1 _20200_/B sky130_fd_sc_hd__nor3_1
XFILLER_193_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20669__B _21124_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17324__A _17391_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14760_ _15254_/A _14760_/B _15254_/C vssd1 vssd1 vccd1 vccd1 _14760_/X sky130_fd_sc_hd__and3_1
XFILLER_57_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ _11972_/A vssd1 vssd1 vccd1 vccd1 _11972_/X sky130_fd_sc_hd__buf_2
XANTENNA__12285__A2 _12238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13711_ _13711_/A _13711_/B _13711_/C vssd1 vssd1 vccd1 vccd1 _13748_/C sky130_fd_sc_hd__nand3_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22909_ _22966_/S vssd1 vssd1 vccd1 vccd1 _22918_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14691_ _23373_/Q _14688_/X _14690_/X vssd1 vssd1 vccd1 vccd1 _14691_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16430_ _16472_/A _16472_/B _16472_/C vssd1 vssd1 vccd1 vccd1 _16432_/B sky130_fd_sc_hd__and3_1
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ _13642_/A vssd1 vssd1 vccd1 vccd1 _13642_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16389_/A _16300_/A _16306_/A vssd1 vssd1 vccd1 vccd1 _16402_/A sky130_fd_sc_hd__o21ai_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13573_ _13573_/A _22553_/C _13712_/A _13573_/D vssd1 vssd1 vccd1 vccd1 _13756_/B
+ sky130_fd_sc_hd__and4_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18173__A1 _18219_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18100_ _18100_/A vssd1 vssd1 vccd1 vccd1 _18217_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11796__A1 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15312_ _15311_/A _15311_/B _15366_/A _15166_/Y vssd1 vssd1 vccd1 vccd1 _15312_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19080_ _18901_/X _19077_/Y _19078_/Y _19079_/Y vssd1 vssd1 vccd1 vccd1 _19080_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12524_ _12536_/A _12528_/B _12527_/A vssd1 vssd1 vccd1 vccd1 _12529_/A sky130_fd_sc_hd__a21o_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _17035_/C _17974_/D _18172_/D _17326_/D vssd1 vssd1 vccd1 vccd1 _16292_/X
+ sky130_fd_sc_hd__and4_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16184__B1 _15937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18031_ _18033_/A _18033_/B _18032_/B _18032_/A vssd1 vssd1 vccd1 vccd1 _18037_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15243_ _14773_/Y _15241_/Y _15242_/X vssd1 vssd1 vccd1 vccd1 _15245_/C sky130_fd_sc_hd__o21a_1
X_12455_ _19648_/A _19530_/D _12455_/C _12455_/D vssd1 vssd1 vccd1 vccd1 _12455_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19673__A1 _19675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15174_ _14181_/X _15375_/A _15173_/Y vssd1 vssd1 vccd1 vccd1 _15179_/B sky130_fd_sc_hd__o21ai_1
XFILLER_67_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12386_ _12059_/A _12200_/B _12205_/A _12059_/D vssd1 vssd1 vccd1 vccd1 _12388_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_158_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14125_ _13965_/X _14086_/A _14029_/C _13922_/D _14124_/Y vssd1 vssd1 vccd1 vccd1
+ _14125_/Y sky130_fd_sc_hd__a41oi_2
XFILLER_193_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19982_ _20073_/A _20073_/B _20073_/C vssd1 vssd1 vccd1 vccd1 _19982_/Y sky130_fd_sc_hd__nand3_1
XFILLER_181_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12931__A _20773_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18933_ _18765_/B _18932_/Y _18759_/Y vssd1 vssd1 vccd1 vccd1 _18944_/C sky130_fd_sc_hd__o21ai_4
XFILLER_141_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output77_A _14717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14056_ _14056_/A _14056_/B _14056_/C vssd1 vssd1 vccd1 vccd1 _14285_/B sky130_fd_sc_hd__nand3_2
XFILLER_97_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12650__B _13121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16122__B _16122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17436__B1 _15682_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ _13005_/Y _13001_/X _13029_/B vssd1 vssd1 vccd1 vccd1 _13007_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__19976__A2 _17763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_983 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15019__A _15019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18864_ _18828_/Y _18840_/Y _18875_/C _18875_/B vssd1 vssd1 vccd1 vccd1 _18864_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_94_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17987__B2 _20210_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17815_ _17817_/A _17817_/B vssd1 vssd1 vccd1 vccd1 _17832_/D sky130_fd_sc_hd__nand2_4
X_18795_ _18639_/B _18804_/A _18443_/A _18453_/A vssd1 vssd1 vccd1 vccd1 _18802_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14858__A _14858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23319__CLK input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17746_ _17840_/A _17840_/B _17750_/B _17745_/Y vssd1 vssd1 vccd1 vccd1 _17759_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12276__A2 _11760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14958_ _15065_/A _15065_/B _14959_/C _15065_/C vssd1 vssd1 vccd1 vccd1 _14960_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17739__A1 _17285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18936__B1 _18938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ _14011_/B vssd1 vssd1 vccd1 vccd1 _13946_/A sky130_fd_sc_hd__clkbuf_2
X_17677_ _17705_/A _17705_/B _17677_/C vssd1 vssd1 vccd1 vccd1 _17680_/C sky130_fd_sc_hd__nand3_4
XFILLER_39_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12378__A _12378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14889_ _14889_/A _14889_/B vssd1 vssd1 vccd1 vccd1 _14890_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19416_ _19242_/Y _19415_/Y _19244_/B vssd1 vssd1 vccd1 vccd1 _19416_/Y sky130_fd_sc_hd__a21oi_1
X_16628_ _15863_/A _16146_/A _16627_/X vssd1 vssd1 vccd1 vccd1 _16628_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17888__B _18016_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19347_ _19345_/X _19346_/Y _19350_/A _19325_/Y vssd1 vssd1 vccd1 vccd1 _19470_/A
+ sky130_fd_sc_hd__o211ai_2
X_16559_ _16500_/Y _16503_/Y _16545_/Y _16555_/Y vssd1 vssd1 vccd1 vccd1 _16559_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__18164__A1 _18163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19278_ _19284_/C _19293_/A _19278_/C vssd1 vssd1 vccd1 vccd1 _19278_/X sky130_fd_sc_hd__and3_1
XFILLER_148_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18229_ _20269_/D _18157_/C _18212_/X _18165_/A vssd1 vssd1 vccd1 vccd1 _18231_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12736__B1 _21271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21240_ _21240_/A _21240_/B vssd1 vssd1 vccd1 vccd1 _21240_/Y sky130_fd_sc_hd__nor2_1
XFILLER_191_658 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17409__A _17409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21171_ _20662_/A _20662_/B _20957_/A vssd1 vssd1 vccd1 vccd1 _21453_/D sky130_fd_sc_hd__a21oi_2
XFILLER_85_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19327__C _19804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20122_ _20118_/X _20113_/B _20025_/B _20117_/X _20121_/X vssd1 vssd1 vccd1 vccd1
+ _20122_/X sky130_fd_sc_hd__a311o_1
XFILLER_172_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20053_ _20210_/C _18211_/B _20056_/A vssd1 vssd1 vccd1 vccd1 _20054_/C sky130_fd_sc_hd__o21ai_1
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17978__A1 _16638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22971__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater140 _23435_/CLK vssd1 vssd1 vccd1 vccd1 _23434_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater151 _23432_/CLK vssd1 vssd1 vccd1 vccd1 _23433_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20489__B _21493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_444 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ _20955_/A _21302_/A _20955_/C vssd1 vssd1 vccd1 vccd1 _20955_/X sky130_fd_sc_hd__and3_1
XANTENNA__16983__A _16988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20886_/A _21124_/B vssd1 vssd1 vccd1 vccd1 _20890_/A sky130_fd_sc_hd__nand2_1
XFILLER_42_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22625_ _22818_/A _22818_/B _22626_/A vssd1 vssd1 vccd1 vccd1 _22627_/A sky130_fd_sc_hd__a21o_1
XFILLER_179_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1020 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11920__A _23591_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22556_ _22649_/C _22556_/B vssd1 vssd1 vccd1 vccd1 _22556_/X sky130_fd_sc_hd__or2_1
XFILLER_50_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21507_ _21510_/C _21507_/B vssd1 vssd1 vccd1 vccd1 _21508_/B sky130_fd_sc_hd__nand2_1
XFILLER_181_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14008__A _23496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22487_ _22487_/A vssd1 vssd1 vccd1 vccd1 _22670_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12240_ _12240_/A vssd1 vssd1 vccd1 vccd1 _16523_/B sky130_fd_sc_hd__buf_4
XANTENNA__19655__A1 _16437_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21438_ _21438_/A vssd1 vssd1 vccd1 vccd1 _21552_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12171_ _11851_/A _11852_/A _18600_/C _16122_/B _16122_/A vssd1 vssd1 vccd1 vccd1
+ _12171_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_162_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21369_ _21369_/A vssd1 vssd1 vccd1 vccd1 _21371_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23108_ _23380_/Q input30/X _23110_/S vssd1 vssd1 vccd1 vccd1 _23109_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21214__A1 _21218_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15930_ _16251_/A _16237_/A _15926_/X _15929_/Y vssd1 vssd1 vccd1 vccd1 _15948_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_122_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23039_ _23039_/A vssd1 vssd1 vccd1 vccd1 _23349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22962__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _15861_/A vssd1 vssd1 vccd1 vccd1 _15861_/X sky130_fd_sc_hd__buf_2
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _17600_/A vssd1 vssd1 vccd1 vccd1 _17613_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _14809_/Y _14810_/X _14811_/X vssd1 vssd1 vccd1 vccd1 _14825_/A sky130_fd_sc_hd__o21ai_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _12564_/Y _18749_/A _12565_/X _18574_/X _18579_/Y vssd1 vssd1 vccd1 vccd1
+ _18589_/A sky130_fd_sc_hd__o32ai_2
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12258__A2 _16364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15792_ _11792_/A _11792_/B _15644_/X _15791_/X _15647_/B vssd1 vssd1 vccd1 vccd1
+ _15792_/X sky130_fd_sc_hd__a221o_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22895__A _22895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22714__A1 _22713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _17943_/A _17530_/Y _17212_/A vssd1 vssd1 vccd1 vccd1 _17531_/X sky130_fd_sc_hd__o21a_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14743_ _14734_/X _11647_/B _14738_/X vssd1 vssd1 vccd1 vccd1 _23266_/D sky130_fd_sc_hd__a21o_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _11856_/X _11850_/Y _11844_/Y vssd1 vssd1 vccd1 vccd1 _11967_/A sky130_fd_sc_hd__a21o_1
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12629__C _13052_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17462_ _17473_/A _17473_/B vssd1 vssd1 vccd1 vccd1 _17462_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14674_ _23337_/Q _14668_/X _14673_/X _23305_/Q _14657_/X vssd1 vssd1 vccd1 vccd1
+ _14674_/X sky130_fd_sc_hd__a221o_1
XANTENNA__19700__C _19700_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11886_ _11886_/A vssd1 vssd1 vccd1 vccd1 _18445_/B sky130_fd_sc_hd__clkbuf_2
X_19201_ _19201_/A _19709_/A _19201_/C _19847_/C vssd1 vssd1 vccd1 vccd1 _19201_/Y
+ sky130_fd_sc_hd__nand4_4
X_16413_ _16167_/C _17406_/A _17406_/B _17723_/C _16549_/C vssd1 vssd1 vccd1 vccd1
+ _16469_/B sky130_fd_sc_hd__a32o_1
XFILLER_177_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13625_ _13486_/B _13613_/A _22484_/A _13486_/A vssd1 vssd1 vccd1 vccd1 _13625_/X
+ sky130_fd_sc_hd__o22a_2
X_17393_ _17393_/A vssd1 vssd1 vccd1 vccd1 _17810_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12926__A _21036_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19132_ _19391_/A _19354_/B vssd1 vssd1 vccd1 vccd1 _19134_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11830__A _11830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16344_ _16576_/B _16339_/X _16575_/A vssd1 vssd1 vccd1 vccd1 _16582_/C sky130_fd_sc_hd__o21ai_4
X_13556_ _13554_/X _13555_/Y _13507_/Y _13494_/Y vssd1 vssd1 vccd1 vccd1 _13556_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_964 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater98 hold23/A vssd1 vssd1 vccd1 vccd1 _15574_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_40_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19063_ _19063_/A _19063_/B _19063_/C vssd1 vssd1 vccd1 vccd1 _19071_/A sky130_fd_sc_hd__nand3_2
X_12507_ _15868_/A vssd1 vssd1 vccd1 vccd1 _19543_/B sky130_fd_sc_hd__buf_2
XFILLER_160_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19709__A _19709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16275_ _16275_/A _16281_/C _16281_/D vssd1 vssd1 vccd1 vccd1 _16275_/X sky130_fd_sc_hd__and3_1
XFILLER_173_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13487_ _21793_/A _13566_/D vssd1 vssd1 vccd1 vccd1 _13487_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18014_ _18114_/A _18014_/B vssd1 vssd1 vccd1 vccd1 _18014_/Y sky130_fd_sc_hd__nand2_1
X_15226_ _15538_/C _15201_/B _15075_/A _15225_/X vssd1 vssd1 vccd1 vccd1 _15292_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12438_ _12438_/A _12438_/B _12438_/C vssd1 vssd1 vccd1 vccd1 _18497_/A sky130_fd_sc_hd__nand3_2
XANTENNA__22245__A3 _21981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15157_ _15120_/D _15121_/A _15154_/X _15156_/X vssd1 vssd1 vccd1 vccd1 _15159_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12369_ _12366_/A _12372_/A _12368_/Y vssd1 vssd1 vccd1 vccd1 _12369_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14108_ _23497_/Q vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__inv_2
X_19965_ _19218_/X _17976_/A _19803_/X _17565_/X vssd1 vssd1 vccd1 vccd1 _19967_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15088_ _14981_/X _14976_/Y _14985_/X _15090_/A _15090_/B vssd1 vssd1 vccd1 vccd1
+ _15092_/A sky130_fd_sc_hd__o2111ai_1
XANTENNA__16880__A1 _16319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15683__A2 _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18916_ _18911_/X _18912_/Y _18915_/Y vssd1 vssd1 vccd1 vccd1 _18918_/A sky130_fd_sc_hd__o21ai_1
X_14039_ _14039_/A _14116_/A vssd1 vssd1 vccd1 vccd1 _14039_/Y sky130_fd_sc_hd__nand2_1
X_19896_ _19896_/A _19896_/B vssd1 vssd1 vccd1 vccd1 _20017_/A sky130_fd_sc_hd__nand2_1
XANTENNA__21756__A2 _22484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18847_ _11822_/A _12053_/A _12007_/Y _18657_/Y vssd1 vssd1 vccd1 vccd1 _18959_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16632__A1 _15731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12249__A2 _12247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18778_ _18778_/A _18778_/B _18778_/C vssd1 vssd1 vccd1 vccd1 _19087_/C sky130_fd_sc_hd__and3_1
XFILLER_67_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17729_ _17629_/Y _18161_/B _18017_/D _17728_/X vssd1 vssd1 vccd1 vccd1 _17729_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22181__A2 _21853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15199__A1 _14029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20740_ _20868_/A _20867_/A _20867_/B vssd1 vssd1 vccd1 vccd1 _20740_/Y sky130_fd_sc_hd__nand3_1
XFILLER_51_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20671_ _20782_/A vssd1 vssd1 vccd1 vccd1 _21431_/A sky130_fd_sc_hd__buf_2
XFILLER_51_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16308__A _16674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23130__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22410_ _22410_/A _22509_/A _22504_/A vssd1 vssd1 vccd1 vccd1 _22410_/Y sky130_fd_sc_hd__nand3_1
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23390_ _23396_/CLK _23390_/D vssd1 vssd1 vccd1 vccd1 _23390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_986 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22341_ _22341_/A _22341_/B _22341_/C vssd1 vssd1 vccd1 vccd1 _22342_/B sky130_fd_sc_hd__and3_1
XFILLER_192_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22272_ _22474_/C _22269_/Y _22271_/Y vssd1 vssd1 vccd1 vccd1 _22272_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15866__B _15866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22045__A _22045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21223_ _21115_/A _21106_/A _21106_/B vssd1 vssd1 vccd1 vccd1 _21223_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_105_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16043__A _17098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21154_ _21150_/Y _21152_/Y _21153_/Y _21132_/Y vssd1 vssd1 vccd1 vccd1 _21154_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__16320__B1 _16458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13386__B _13804_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18860__A2 _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20105_ _20106_/B _20106_/C _20106_/A vssd1 vssd1 vccd1 vccd1 _20111_/B sky130_fd_sc_hd__a21o_1
XFILLER_59_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16871__A1 _16604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15882__A _15882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14477__A3 _13972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16871__B2 _11926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21085_ _21097_/C vssd1 vssd1 vccd1 vccd1 _21212_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14882__B1 _14883_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20036_ _19923_/Y _19789_/Y _19920_/A _20035_/Y vssd1 vssd1 vccd1 vccd1 _20201_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_112_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18612__A2 _12168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11915__A _11915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11634__B _11634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21987_ _21987_/A _21987_/B _21987_/C vssd1 vssd1 vccd1 vccd1 _21989_/B sky130_fd_sc_hd__and3_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11860_/B vssd1 vssd1 vccd1 vccd1 _11740_/X sky130_fd_sc_hd__buf_4
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _20943_/A _20943_/B _20947_/A _20947_/B vssd1 vssd1 vccd1 vccd1 _20945_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_148_1164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15016__A2_N _15366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _23384_/Q vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__buf_2
XFILLER_169_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20869_ _20885_/A _20869_/B _20885_/B vssd1 vssd1 vccd1 vccd1 _20872_/C sky130_fd_sc_hd__nand3_1
XFILLER_168_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23121__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13410_ _13410_/A vssd1 vssd1 vccd1 vccd1 _13410_/X sky130_fd_sc_hd__buf_2
X_22608_ _22610_/A _22606_/Y _22609_/A _22609_/B vssd1 vssd1 vccd1 vccd1 _22631_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18679__A2 _19334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14390_ _14390_/A _14390_/B _14390_/C vssd1 vssd1 vccd1 vccd1 _14442_/A sky130_fd_sc_hd__nand3_1
X_23588_ _23588_/CLK _23588_/D vssd1 vssd1 vccd1 vccd1 _23588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17887__B1 _17960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ _13456_/A _13456_/B _13269_/A vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__a21o_1
XFILLER_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22539_ _22729_/A _22729_/B vssd1 vssd1 vccd1 vccd1 _22540_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21778__B _22364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16060_ _16060_/A _16060_/B _16060_/C vssd1 vssd1 vccd1 vccd1 _16326_/A sky130_fd_sc_hd__nand3_4
XFILLER_154_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13272_ _13498_/A vssd1 vssd1 vccd1 vccd1 _13741_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_850 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15362__B2 _15415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15011_ _14976_/A _14983_/A _15371_/B _14985_/X _15262_/A vssd1 vssd1 vccd1 vccd1
+ _15013_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_68_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12223_ _12223_/A vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__buf_2
XFILLER_120_1072 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11923__A1 _11916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21986__A2 _21988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20643__C1 _20894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ _12131_/Y _12134_/Y _12122_/Y vssd1 vssd1 vccd1 vccd1 _12399_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11809__B _16796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19750_ _19734_/Y _19735_/Y _19736_/Y _19733_/C vssd1 vssd1 vccd1 vccd1 _19750_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12085_ _12509_/A vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16962_ _16735_/C _16721_/Y _16735_/B vssd1 vssd1 vccd1 vccd1 _16964_/C sky130_fd_sc_hd__o21ai_2
XFILLER_89_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18701_ _18689_/X _18692_/X _18667_/Y _18672_/Y vssd1 vssd1 vccd1 vccd1 _18701_/Y
+ sky130_fd_sc_hd__o211ai_1
X_15913_ _15719_/B _15908_/Y _15721_/X vssd1 vssd1 vccd1 vccd1 _15916_/A sky130_fd_sc_hd__o21a_1
X_19681_ _19669_/X _19680_/X _19673_/Y _19676_/X vssd1 vssd1 vccd1 vccd1 _19685_/A
+ sky130_fd_sc_hd__o22ai_2
X_16893_ _16893_/A _16893_/B _16893_/C vssd1 vssd1 vccd1 vccd1 _16894_/C sky130_fd_sc_hd__nand3_1
XANTENNA__15417__A2 _15446_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15844_ _15844_/A vssd1 vssd1 vccd1 vccd1 _15993_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18632_ _11864_/X _11865_/X _18439_/X _18440_/X _19805_/A vssd1 vssd1 vccd1 vccd1
+ _18632_/Y sky130_fd_sc_hd__o221ai_2
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18563_ _12522_/C _18559_/X _18728_/A _18562_/Y vssd1 vssd1 vccd1 vccd1 _18584_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15775_ _16480_/A _15802_/B _17409_/A _15772_/X _15641_/Y vssd1 vssd1 vccd1 vccd1
+ _15775_/X sky130_fd_sc_hd__o311a_1
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18367__A1 _23534_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _12985_/A _13088_/B _20464_/D vssd1 vssd1 vccd1 vccd1 _12987_/Y sky130_fd_sc_hd__o21ai_4
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _23596_/Q vssd1 vssd1 vccd1 vccd1 _16815_/D sky130_fd_sc_hd__buf_2
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ _17514_/A _17514_/B _17514_/C _17514_/D vssd1 vssd1 vccd1 vccd1 _17700_/B
+ sky130_fd_sc_hd__nand4_1
X_11938_ _11856_/X _11850_/Y _11844_/Y vssd1 vssd1 vccd1 vccd1 _11938_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16378__B1 _16377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18494_ _12445_/C _12423_/A _12423_/B _12451_/Y vssd1 vssd1 vccd1 vccd1 _18495_/C
+ sky130_fd_sc_hd__a31oi_2
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _17445_/A _17581_/A _18778_/B vssd1 vssd1 vccd1 vccd1 _17446_/B sky130_fd_sc_hd__and3_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14657_ _14657_/A vssd1 vssd1 vccd1 vccd1 _14657_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11869_ _11738_/X _11740_/X _11741_/Y vssd1 vssd1 vccd1 vccd1 _16044_/A sky130_fd_sc_hd__o21ai_4
XFILLER_14_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13608_ _21752_/A _21752_/B _22024_/C vssd1 vssd1 vccd1 vccd1 _13793_/A sky130_fd_sc_hd__nand3_1
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17376_ _17376_/A vssd1 vssd1 vccd1 vccd1 _18059_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_159_964 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14588_ _14588_/A vssd1 vssd1 vccd1 vccd1 _14588_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19115_ _19116_/A _19116_/B _19116_/C vssd1 vssd1 vccd1 vccd1 _19133_/A sky130_fd_sc_hd__a21oi_1
X_16327_ _16094_/A _16052_/X _16331_/A vssd1 vssd1 vccd1 vccd1 _16327_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__20477__A2 _20471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15967__A _15998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13539_ _13477_/X _13598_/A _13538_/X vssd1 vssd1 vccd1 vccd1 _13540_/C sky130_fd_sc_hd__a21o_1
XFILLER_71_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19046_ _19047_/A _19047_/C _19047_/B vssd1 vssd1 vccd1 vccd1 _19046_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_174_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16258_ _16258_/A _16258_/B _16258_/C vssd1 vssd1 vccd1 vccd1 _16268_/D sky130_fd_sc_hd__nand3_2
XFILLER_145_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15209_ _15208_/Y _15077_/X _15076_/Y vssd1 vssd1 vccd1 vccd1 _15282_/B sky130_fd_sc_hd__o21bai_2
XFILLER_160_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ _15604_/X _16658_/C _16667_/D _16668_/C vssd1 vssd1 vccd1 vccd1 _16671_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_126_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18997__B _18997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11719__B _11907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19948_ _19948_/A _19948_/B vssd1 vssd1 vccd1 vccd1 _20217_/B sky130_fd_sc_hd__nand2_4
XFILLER_101_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11678__B1 _11677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19879_ _19879_/A _19879_/B _19879_/C vssd1 vssd1 vccd1 vccd1 _19897_/A sky130_fd_sc_hd__nand3_1
XANTENNA__17406__B _17406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16605__A1 _15698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16605__B2 _11936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21910_ _21913_/A _21910_/B vssd1 vssd1 vccd1 vccd1 _21911_/C sky130_fd_sc_hd__nand2_1
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11735__A _16364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13419__A1 _13415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14111__A _23496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22890_ _22891_/A _22891_/C _22891_/B vssd1 vssd1 vccd1 vccd1 _22895_/B sky130_fd_sc_hd__a21oi_4
X_21841_ _21835_/Y _21838_/X _21847_/C vssd1 vssd1 vccd1 vccd1 _21842_/A sky130_fd_sc_hd__o21bai_4
XFILLER_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19555__B1 _19554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22154__A2 _22164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17422__A _17625_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_572 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21772_ _13410_/X _21762_/Y _22276_/A _22264_/B _21984_/A vssd1 vssd1 vccd1 vccd1
+ _21772_/X sky130_fd_sc_hd__o2111a_1
XANTENNA__17030__A1 _16781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23511_ _23518_/CLK input47/X vssd1 vssd1 vccd1 vccd1 _23511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20723_ _20589_/A _20589_/C _20578_/X vssd1 vssd1 vccd1 vccd1 _20724_/C sky130_fd_sc_hd__a21oi_1
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19307__B1 _19308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23442_ _23442_/CLK _23442_/D vssd1 vssd1 vccd1 vccd1 _23442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20654_ _20624_/X _20631_/X _20636_/X _20653_/Y vssd1 vssd1 vccd1 vccd1 _20654_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15877__A _19363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20585_ _20585_/A _20585_/B vssd1 vssd1 vccd1 vccd1 _20585_/Y sky130_fd_sc_hd__nand2_1
X_23373_ _23377_/CLK _23373_/D vssd1 vssd1 vccd1 vccd1 _23373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_720 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22324_ _22324_/A _22324_/B _22324_/C vssd1 vssd1 vccd1 vccd1 _22332_/B sky130_fd_sc_hd__nand3_2
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16541__B1 _16531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22255_ _22451_/A _22451_/B _22451_/C _22452_/A vssd1 vssd1 vccd1 vccd1 _22355_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_191_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19086__A2 _12168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21206_ _21206_/A vssd1 vssd1 vccd1 vccd1 _21270_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_544 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22186_ _22142_/B _22186_/B _22186_/C vssd1 vssd1 vccd1 vccd1 _22187_/B sky130_fd_sc_hd__nand3b_2
XANTENNA__15536__D_N _15225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21137_ _21003_/X _21020_/Y _21241_/C vssd1 vssd1 vccd1 vccd1 _21344_/A sky130_fd_sc_hd__o21ai_1
XFILLER_28_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21068_ _20900_/Y _20909_/X _20905_/Y vssd1 vssd1 vccd1 vccd1 _21069_/C sky130_fd_sc_hd__a21boi_2
XFILLER_120_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12866__C1 _21174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12330__A1 _12323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20019_ _20015_/X _20016_/Y _20018_/X vssd1 vssd1 vccd1 vccd1 _20021_/A sky130_fd_sc_hd__a21oi_2
X_12910_ _12975_/C _12975_/B _12975_/A vssd1 vssd1 vccd1 vccd1 _12910_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_4_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13890_ _13890_/A _13890_/B vssd1 vssd1 vccd1 vccd1 _14386_/B sky130_fd_sc_hd__nand2_1
XFILLER_73_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_bq_clk_i clkbuf_2_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12841_ _21193_/C vssd1 vssd1 vccd1 vccd1 _13131_/A sky130_fd_sc_hd__buf_2
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18428__A _23538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15528_/A _15552_/A _15552_/B vssd1 vssd1 vccd1 vccd1 _15561_/B sky130_fd_sc_hd__o21ai_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12845_/A _12901_/A vssd1 vssd1 vccd1 vccd1 _12774_/A sky130_fd_sc_hd__nand2_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ input1/X vssd1 vssd1 vccd1 vccd1 _14633_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11723_/A vssd1 vssd1 vccd1 vccd1 _11916_/A sky130_fd_sc_hd__buf_2
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _15446_/X _15447_/Y _15488_/X _15489_/X vssd1 vssd1 vccd1 vccd1 _15508_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17230_/A vssd1 vssd1 vccd1 vccd1 _17752_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14442_/A _14442_/B vssd1 vssd1 vccd1 vccd1 _14443_/A sky130_fd_sc_hd__nand2_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11654_ _11654_/A vssd1 vssd1 vccd1 vccd1 _11844_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_156_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17161_ _17161_/A _17161_/B vssd1 vssd1 vccd1 vccd1 _17163_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14373_ _13890_/A _13890_/B _14097_/A vssd1 vssd1 vccd1 vccd1 _14374_/C sky130_fd_sc_hd__a21oi_1
XFILLER_122_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11585_ _16593_/A vssd1 vssd1 vccd1 vccd1 _19017_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__18163__A _18163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16112_ _18093_/A vssd1 vssd1 vccd1 vccd1 _18172_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_155_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13324_ _13366_/B _13323_/X _13253_/A vssd1 vssd1 vccd1 vccd1 _13325_/B sky130_fd_sc_hd__o21ai_1
XFILLER_196_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17092_ _17092_/A vssd1 vssd1 vccd1 vccd1 _17712_/B sky130_fd_sc_hd__buf_4
XFILLER_171_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16043_ _17098_/B vssd1 vssd1 vccd1 vccd1 _17226_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_7_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13255_ _13660_/C _13660_/A vssd1 vssd1 vccd1 vccd1 _13256_/A sky130_fd_sc_hd__nand2_1
XFILLER_170_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ _12206_/A vssd1 vssd1 vccd1 vccd1 _18559_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13186_ _13186_/A _20726_/D _13186_/C vssd1 vssd1 vccd1 vccd1 _13188_/B sky130_fd_sc_hd__and3_1
X_19802_ _19802_/A _19802_/B vssd1 vssd1 vccd1 vccd1 _19822_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17507__A _18211_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ _12010_/B _12125_/Y _12122_/Y _12119_/Y vssd1 vssd1 vccd1 vccd1 _12138_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_151_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19425__C _19425_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17994_ _17994_/A _17994_/B _17994_/C vssd1 vssd1 vccd1 vccd1 _17994_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__16411__A _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19733_ _19733_/A _19733_/B _19733_/C vssd1 vssd1 vccd1 vccd1 _19733_/Y sky130_fd_sc_hd__nand3_1
XFILLER_78_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17226__B _17860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16945_ _16924_/Y _17166_/B _16937_/Y vssd1 vssd1 vccd1 vccd1 _16945_/Y sky130_fd_sc_hd__a21oi_1
X_12068_ _11969_/A _11969_/B _12227_/A vssd1 vssd1 vccd1 vccd1 _12080_/B sky130_fd_sc_hd__a21boi_2
XANTENNA__16048__C1 _16451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19664_ _19674_/A _19664_/B _19674_/C _19969_/A vssd1 vssd1 vccd1 vccd1 _19665_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__21971__B _21971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16876_ _16885_/A _16894_/B _16873_/X _16875_/Y vssd1 vssd1 vccd1 vccd1 _16888_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_93_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16063__A2 _16073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18615_ _18615_/A _18615_/B _18615_/C vssd1 vssd1 vccd1 vccd1 _18615_/Y sky130_fd_sc_hd__nand3_4
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _15827_/A _15827_/B vssd1 vssd1 vccd1 vccd1 _15836_/A sky130_fd_sc_hd__nand2_1
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19595_ _19572_/X _19376_/A _19573_/C _19587_/A _19747_/A vssd1 vssd1 vccd1 vccd1
+ _19595_/Y sky130_fd_sc_hd__o2111ai_2
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17242__A _19334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20147__A1 _20146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18546_ _12528_/A _12537_/B _12528_/B vssd1 vssd1 vccd1 vccd1 _18562_/A sky130_fd_sc_hd__a21boi_1
X_15758_ _16612_/A vssd1 vssd1 vccd1 vccd1 _16160_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__19001__A2 _16033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13821__A1 _13552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14709_ _23346_/Q _14531_/A _14694_/X _23314_/Q _14699_/X vssd1 vssd1 vccd1 vccd1
+ _14709_/X sky130_fd_sc_hd__a221o_1
X_18477_ _12410_/Y _18434_/A _18476_/X vssd1 vssd1 vccd1 vccd1 _20320_/B sky130_fd_sc_hd__a21o_2
X_15689_ _15656_/X _15727_/B _15664_/A vssd1 vssd1 vccd1 vccd1 _16591_/D sky130_fd_sc_hd__a21o_2
X_17428_ _17485_/A _17485_/B _17485_/C vssd1 vssd1 vccd1 vccd1 _17487_/A sky130_fd_sc_hd__a21o_1
XFILLER_127_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17359_ _17359_/A _17359_/B vssd1 vssd1 vccd1 vccd1 _17362_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17315__A2 _17635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18512__B2 _18503_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20370_ _18335_/B _19862_/B _19862_/C _20369_/X vssd1 vssd1 vccd1 vccd1 _20371_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_147_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19029_ _19029_/A _19029_/B _19029_/C _19029_/D vssd1 vssd1 vccd1 vccd1 _19139_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_173_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_959 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22040_ _22040_/A _22040_/B vssd1 vssd1 vccd1 vccd1 _22040_/Y sky130_fd_sc_hd__nand2_2
XFILLER_47_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1035 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22942_ _22953_/A vssd1 vssd1 vccd1 vccd1 _22951_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_141_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12863__A2 _12862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22873_ _22874_/B _22874_/C _22874_/A vssd1 vssd1 vccd1 vccd1 _22873_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__19528__B1 _19332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15801__A2 _11740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21824_ _21824_/A _21824_/B _21824_/C vssd1 vssd1 vccd1 vccd1 _21844_/B sky130_fd_sc_hd__nand3_2
XFILLER_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18200__B1 _18154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__B _11912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21755_ _21755_/A vssd1 vssd1 vccd1 vccd1 _21755_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_197_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1014 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16991__A _17217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20706_ _20553_/B _20547_/C _20702_/Y _20534_/X vssd1 vssd1 vccd1 vccd1 _20725_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21686_ _21704_/B _21684_/Y _23573_/Q _21685_/X vssd1 vssd1 vccd1 vccd1 _21688_/D
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__17378__A_N _23525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23425_ _23425_/CLK _23425_/D vssd1 vssd1 vccd1 vccd1 _23425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20637_ _23298_/Q vssd1 vssd1 vccd1 vccd1 _20641_/A sky130_fd_sc_hd__inv_2
XFILLER_138_945 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17306__A2 _16033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_764 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16514__B1 _12379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23356_ _23359_/CLK _23356_/D vssd1 vssd1 vccd1 vccd1 _23356_/Q sky130_fd_sc_hd__dfxtp_1
X_20568_ _20579_/A _20570_/A _20566_/X _20567_/Y vssd1 vssd1 vccd1 vccd1 _20568_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_192_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22307_ _22403_/A _22405_/B _22405_/C vssd1 vssd1 vccd1 vccd1 _22314_/A sky130_fd_sc_hd__a21oi_1
XFILLER_125_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23287_ _23297_/CLK _23287_/D vssd1 vssd1 vccd1 vccd1 _23287_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_180_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20499_ _20782_/B vssd1 vssd1 vccd1 vccd1 _21431_/B sky130_fd_sc_hd__buf_2
XFILLER_106_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13040_ _13028_/Y _13032_/X _20557_/A _20557_/B vssd1 vssd1 vccd1 vccd1 _13078_/A
+ sky130_fd_sc_hd__o211ai_4
X_22238_ _22237_/X _22096_/B _22090_/D _21989_/C vssd1 vssd1 vccd1 vccd1 _22238_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_65_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22169_ _22057_/X _22168_/X _22280_/B _22391_/A vssd1 vssd1 vccd1 vccd1 _22169_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16293__A2 _18172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12839__C1 _12845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ _14991_/A vssd1 vssd1 vccd1 vccd1 _15000_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_input39_A wb_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13942_ _14096_/A vssd1 vssd1 vccd1 vccd1 _13942_/X sky130_fd_sc_hd__clkbuf_2
X_16730_ _16715_/Y _16718_/Y _16720_/Y vssd1 vssd1 vccd1 vccd1 _16735_/A sky130_fd_sc_hd__a21o_1
XFILLER_93_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_634 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16045__A2 _11801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23064__A _23110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16661_ _16661_/A _19308_/B _16661_/C _17148_/A vssd1 vssd1 vccd1 vccd1 _16662_/B
+ sky130_fd_sc_hd__nand4_4
X_13873_ _21971_/B _23270_/Q vssd1 vssd1 vccd1 vccd1 _13875_/A sky130_fd_sc_hd__and2_1
XFILLER_75_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18400_ _18400_/A _18414_/C _18400_/C vssd1 vssd1 vccd1 vccd1 _18400_/X sky130_fd_sc_hd__and3_1
X_15612_ _15612_/A _15612_/B vssd1 vssd1 vccd1 vccd1 _16113_/A sky130_fd_sc_hd__nand2_4
XANTENNA__17062__A _17761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ _12824_/A _12824_/B vssd1 vssd1 vccd1 vccd1 _12835_/D sky130_fd_sc_hd__and2_1
X_19380_ _18673_/A _17846_/X _17431_/A _12324_/X vssd1 vssd1 vccd1 vccd1 _19380_/X
+ sky130_fd_sc_hd__o22a_2
X_16592_ _16592_/A _16592_/B vssd1 vssd1 vccd1 vccd1 _16601_/C sky130_fd_sc_hd__nand2_1
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22669__A3 _22476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18331_ _19900_/A vssd1 vssd1 vccd1 vccd1 _18335_/B sky130_fd_sc_hd__buf_2
X_15543_ _15543_/A _15543_/B vssd1 vssd1 vccd1 vccd1 _15544_/B sky130_fd_sc_hd__and2_1
XFILLER_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _23294_/Q vssd1 vssd1 vccd1 vccd1 _12756_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_884 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18262_/A _18262_/B _18262_/C vssd1 vssd1 vccd1 vccd1 _18264_/B sky130_fd_sc_hd__nand3_2
X_11706_ _11820_/A _11844_/B _11705_/Y vssd1 vssd1 vccd1 vccd1 _11717_/C sky130_fd_sc_hd__o21ai_4
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15474_ _15474_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15475_/B sky130_fd_sc_hd__nand2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12674_/X _12766_/A _20509_/A vssd1 vssd1 vccd1 vccd1 _12812_/A sky130_fd_sc_hd__o21ai_4
XFILLER_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17213_ _17212_/C _17212_/A _23524_/Q vssd1 vssd1 vccd1 vccd1 _17382_/A sky130_fd_sc_hd__a21o_1
XFILLER_129_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14425_ _14396_/B _14396_/C _14009_/X _13969_/Y vssd1 vssd1 vccd1 vccd1 _14436_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_187_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18193_ _18155_/A _18155_/B _18133_/A _18133_/B vssd1 vssd1 vccd1 vccd1 _18195_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_11637_ _11637_/A vssd1 vssd1 vccd1 vccd1 _16591_/B sky130_fd_sc_hd__buf_4
XFILLER_128_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17144_ _16360_/X _17635_/A _17150_/A vssd1 vssd1 vccd1 vccd1 _17145_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__15310__A _15371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14356_ _14356_/A _14356_/B _14356_/C vssd1 vssd1 vccd1 vccd1 _14403_/B sky130_fd_sc_hd__nand3_2
XFILLER_155_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ _23322_/Q _23321_/Q vssd1 vssd1 vccd1 vccd1 _13377_/B sky130_fd_sc_hd__nor2_2
XFILLER_143_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17075_ _17565_/A _16632_/X _17074_/X _16824_/Y vssd1 vssd1 vccd1 vccd1 _17075_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14287_ _14273_/X _14283_/X _14285_/Y _14286_/X vssd1 vssd1 vccd1 vccd1 _14367_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_170_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16026_ _16160_/A vssd1 vssd1 vccd1 vccd1 _16308_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__18258__B1 _23533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13238_ _21997_/A _13241_/A vssd1 vssd1 vccd1 vccd1 _21878_/A sky130_fd_sc_hd__nor2_1
XFILLER_170_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15964__B _15964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20065__B1 _20066_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13169_ _13174_/A _13169_/B _13169_/C _13169_/D vssd1 vssd1 vccd1 vccd1 _13191_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__16141__A _16141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11750__C1 _11747_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19207__C1 _11849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17977_ _17285_/X _18096_/A _20210_/A _17465_/X vssd1 vssd1 vccd1 vccd1 _17986_/B
+ sky130_fd_sc_hd__o22ai_4
X_19716_ _19723_/A _19716_/B vssd1 vssd1 vccd1 vccd1 _19722_/A sky130_fd_sc_hd__nand2_1
X_16928_ _16928_/A vssd1 vssd1 vccd1 vccd1 _17304_/A sky130_fd_sc_hd__buf_2
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16036__A2 _15766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19647_ _19656_/A _19491_/B _19667_/D _19675_/A vssd1 vssd1 vccd1 vccd1 _19647_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16859_ _15882_/A _17465_/A _16592_/B _17095_/A _17107_/A vssd1 vssd1 vccd1 vccd1
+ _16879_/B sky130_fd_sc_hd__o221ai_4
XFILLER_1_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15231__D_N _15054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19578_ _19578_/A _19578_/B vssd1 vssd1 vccd1 vccd1 _19578_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12828__B _20532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18529_ _18529_/A _18529_/B vssd1 vssd1 vccd1 vccd1 _18529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21540_ _21540_/A _21540_/B _21540_/C vssd1 vssd1 vccd1 vccd1 _21540_/X sky130_fd_sc_hd__or3_1
XFILLER_194_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_2_0_bq_clk_i_A clkbuf_2_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21471_ _21474_/A vssd1 vssd1 vccd1 vccd1 _21524_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23210_ _23210_/A vssd1 vssd1 vccd1 vccd1 _23424_/D sky130_fd_sc_hd__clkbuf_1
X_20422_ _20393_/A _20393_/B _20418_/Y _20419_/X _20420_/Y vssd1 vssd1 vccd1 vccd1
+ _20423_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_101_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13659__B _13659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23141_ _18799_/B input10/X _23145_/S vssd1 vssd1 vccd1 vccd1 _23142_/A sky130_fd_sc_hd__mux2_1
X_20353_ _20307_/B _20307_/C _20307_/A _20118_/X vssd1 vssd1 vccd1 vccd1 _20354_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18531__A _18531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20284_ _20285_/A _20282_/Y _20283_/Y _20235_/X vssd1 vssd1 vccd1 vccd1 _20284_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23072_ _23072_/A vssd1 vssd1 vccd1 vccd1 _23363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22023_ _21902_/B _22028_/A _22022_/Y vssd1 vssd1 vccd1 vccd1 _22039_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21892__A _21892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15078__A3 _14069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11907__B _11907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15890__A _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14002__C _14433_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22925_ _20894_/B input10/X _22929_/S vssd1 vssd1 vccd1 vccd1 _22926_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19512__D _19512_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22856_ _22856_/A _22856_/B _22856_/C _22856_/D vssd1 vssd1 vccd1 vccd1 _22874_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__17313__C _17313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21807_ _13799_/X _13813_/X _13819_/A _13819_/B vssd1 vssd1 vccd1 vccd1 _21807_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_197_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22787_ _22750_/A _22750_/B _22774_/B vssd1 vssd1 vccd1 vccd1 _22810_/A sky130_fd_sc_hd__a21o_1
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17610__A _17610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12540_ _12540_/A _12540_/B _12540_/C vssd1 vssd1 vccd1 vccd1 _18571_/B sky130_fd_sc_hd__nand3_2
XFILLER_52_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21738_ _13602_/C _21901_/B _21738_/C _21901_/D vssd1 vssd1 vccd1 vccd1 _22047_/B
+ sky130_fd_sc_hd__nand4b_4
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _12177_/B _18675_/C _18506_/A _12461_/Y _12260_/D vssd1 vssd1 vccd1 vccd1
+ _12473_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_185_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21669_ _21637_/A _21668_/B _21637_/C _21635_/X _21668_/Y vssd1 vssd1 vccd1 vccd1
+ _21671_/A sky130_fd_sc_hd__a32o_1
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ _15111_/A _14194_/A _14865_/A vssd1 vssd1 vccd1 vccd1 _14879_/A sky130_fd_sc_hd__o21ai_1
XFILLER_32_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23408_ _23442_/CLK _23408_/D vssd1 vssd1 vccd1 vccd1 _23408_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__22284__A1 _13465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_99 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15190_ _15190_/A _15190_/B vssd1 vssd1 vccd1 vccd1 _15192_/A sky130_fd_sc_hd__nand2_1
XFILLER_126_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13564__A3 _21778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14141_ _14141_/A _14141_/B _14141_/C vssd1 vssd1 vccd1 vccd1 _14230_/A sky130_fd_sc_hd__nand3_2
X_23339_ _23339_/CLK _23339_/D vssd1 vssd1 vccd1 vccd1 _23339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16502__A3 _15682_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14072_ _14070_/X _13927_/A _14865_/A _14188_/A vssd1 vssd1 vccd1 vccd1 _14752_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_152_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17900_ _17898_/X _17899_/X _17896_/Y _18030_/A vssd1 vssd1 vccd1 vccd1 _17901_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13023_ _12952_/A _13025_/A _13022_/Y vssd1 vssd1 vccd1 vccd1 _13041_/A sky130_fd_sc_hd__o21ai_1
XFILLER_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17057__A _17057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18880_ _18880_/A _18880_/B vssd1 vssd1 vccd1 vccd1 _18880_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21795__B1 _13465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22898__A _22966_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17831_ _17831_/A _17831_/B vssd1 vssd1 vccd1 vccd1 _23588_/D sky130_fd_sc_hd__xor2_2
XFILLER_121_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17762_ _18604_/A vssd1 vssd1 vccd1 vccd1 _17763_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19204__A2 _19218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14974_ _15171_/B vssd1 vssd1 vccd1 vccd1 _15317_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19703__C _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19501_ _19492_/C _19500_/X _19321_/A vssd1 vssd1 vccd1 vccd1 _19525_/B sky130_fd_sc_hd__o21ai_1
X_16713_ _16957_/A _16956_/A _16956_/B vssd1 vssd1 vccd1 vccd1 _16713_/Y sky130_fd_sc_hd__a21oi_1
X_13925_ _14173_/A vssd1 vssd1 vccd1 vccd1 _14172_/A sky130_fd_sc_hd__buf_2
X_17693_ _17693_/A _17693_/B _17693_/C vssd1 vssd1 vccd1 vccd1 _17693_/Y sky130_fd_sc_hd__nand3_1
XFILLER_48_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19432_ _19434_/A _19434_/B _19434_/C _19431_/Y vssd1 vssd1 vccd1 vccd1 _19432_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16644_ _16644_/A _16853_/A _16649_/B vssd1 vssd1 vccd1 vccd1 _16655_/A sky130_fd_sc_hd__nand3_1
X_13856_ _13856_/A _13856_/B _13856_/C vssd1 vssd1 vccd1 vccd1 _21839_/A sky130_fd_sc_hd__nand3_2
XFILLER_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12807_ _12796_/X _12801_/Y _12805_/Y vssd1 vssd1 vccd1 vccd1 _12809_/A sky130_fd_sc_hd__o21ai_1
X_19363_ _19363_/A _19363_/B _19363_/C _19363_/D vssd1 vssd1 vccd1 vccd1 _19363_/Y
+ sky130_fd_sc_hd__nand4_4
X_16575_ _16575_/A _16575_/B vssd1 vssd1 vccd1 vccd1 _16576_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13787_ _13339_/A _22141_/A _21738_/C vssd1 vssd1 vccd1 vccd1 _22064_/A sky130_fd_sc_hd__o21ai_4
XFILLER_37_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18314_ _18314_/A _18314_/B _18314_/C _18314_/D vssd1 vssd1 vccd1 vccd1 _18315_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_31_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15526_ _15526_/A _15525_/Y vssd1 vssd1 vccd1 vccd1 _15528_/B sky130_fd_sc_hd__or2b_4
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12738_/A _12738_/B _12738_/C vssd1 vssd1 vccd1 vccd1 _12846_/A sky130_fd_sc_hd__nand3_1
X_19294_ _19095_/Y _19294_/B _19294_/C _19294_/D vssd1 vssd1 vccd1 vccd1 _19295_/A
+ sky130_fd_sc_hd__nand4b_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18335__B _18335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21042__A _21174_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18245_ _18245_/A _18298_/C _18245_/C vssd1 vssd1 vccd1 vccd1 _18267_/A sky130_fd_sc_hd__or3_2
X_15457_ _15457_/A _15457_/B vssd1 vssd1 vccd1 vccd1 _15458_/B sky130_fd_sc_hd__or2_1
XFILLER_198_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ _20493_/B vssd1 vssd1 vccd1 vccd1 _12794_/A sky130_fd_sc_hd__inv_2
XFILLER_129_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12664__A _23452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14408_ _14403_/A _14403_/B _14406_/Y _14407_/X vssd1 vssd1 vccd1 vccd1 _14410_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_128_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18176_ _18176_/A _18176_/B _18227_/A vssd1 vssd1 vccd1 vccd1 _18227_/B sky130_fd_sc_hd__nand3_1
X_15388_ _15538_/C _15388_/B _15388_/C vssd1 vssd1 vccd1 vccd1 _15388_/X sky130_fd_sc_hd__and3_1
XANTENNA__13479__B _22035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17127_ _16878_/Y _16877_/X _16894_/A _16884_/Y vssd1 vssd1 vccd1 vccd1 _17127_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__15975__A _15975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14339_ _14108_/Y _13964_/Y _14381_/A _14333_/X _14334_/Y vssd1 vssd1 vccd1 vccd1
+ _14356_/A sky130_fd_sc_hd__o32a_1
XANTENNA__21696__B _21704_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ _17058_/A _17058_/B vssd1 vssd1 vccd1 vccd1 _17058_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16009_ _16009_/A vssd1 vssd1 vccd1 vccd1 _16347_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1068 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19182__A _19332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14807__A3 _14819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18939__D1 _18080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21217__A _21217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17414__B _17414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20971_ _21302_/A vssd1 vssd1 vccd1 vccd1 _21431_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_26_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21553__A3 _21358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22710_ _22710_/A _22709_/Y vssd1 vssd1 vccd1 vccd1 _22717_/A sky130_fd_sc_hd__or2b_1
XFILLER_54_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11743__A _11743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17133__C _17133_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22641_ _22641_/A _22641_/B _22647_/A vssd1 vssd1 vccd1 vccd1 _22642_/C sky130_fd_sc_hd__nand3_1
XANTENNA__17509__A2 _12379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22572_ _22469_/X _22567_/Y _22468_/X _22650_/B vssd1 vssd1 vccd1 vccd1 _22572_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_181_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20494__C _20798_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21523_ _21524_/A _21524_/B _21524_/C vssd1 vssd1 vccd1 vccd1 _21526_/A sky130_fd_sc_hd__a21o_1
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16193__A1 _12373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21454_ _21455_/B _21455_/A _21377_/A _21377_/C _21453_/X vssd1 vssd1 vccd1 vccd1
+ _21513_/A sky130_fd_sc_hd__a221oi_4
XFILLER_31_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20405_ _20405_/A _20405_/B vssd1 vssd1 vccd1 vccd1 _20408_/B sky130_fd_sc_hd__xnor2_2
XFILLER_175_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21385_ _21386_/A _21490_/B _21386_/C _21386_/B vssd1 vssd1 vccd1 vccd1 _21387_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16496__A2 _16167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23215__A0 _14631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23124_ _23124_/A vssd1 vssd1 vccd1 vccd1 _23386_/D sky130_fd_sc_hd__clkbuf_1
X_20336_ _20336_/A _20336_/B vssd1 vssd1 vccd1 vccd1 _20337_/C sky130_fd_sc_hd__nor2_1
XFILLER_123_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput58 _14639_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[13] sky130_fd_sc_hd__buf_2
X_23055_ _23055_/A vssd1 vssd1 vccd1 vccd1 _23355_/D sky130_fd_sc_hd__clkbuf_1
X_20267_ _20055_/A _20055_/B _20268_/D _20268_/A _20268_/B vssd1 vssd1 vccd1 vccd1
+ _20274_/A sky130_fd_sc_hd__a32o_1
Xoutput69 _14692_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_163_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22006_ _13485_/A _13485_/B _21884_/A _21884_/B _22121_/A vssd1 vssd1 vccd1 vccd1
+ _22006_/X sky130_fd_sc_hd__a221o_1
XFILLER_88_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18642__B1 _18479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20198_ _20199_/B _20199_/C _23551_/Q vssd1 vssd1 vccd1 vccd1 _20311_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17605__A _17605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12552__A1_N _12227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _11971_/A vssd1 vssd1 vccd1 vccd1 _11971_/X sky130_fd_sc_hd__buf_2
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13710_ _13707_/X _13582_/B _13705_/D _13709_/X vssd1 vssd1 vccd1 vccd1 _13711_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22908_ _22908_/A vssd1 vssd1 vccd1 vccd1 _23290_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_648 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14690_ _23341_/Q _14689_/X _14673_/X _23309_/Q _14678_/X vssd1 vssd1 vccd1 vccd1
+ _14690_/X sky130_fd_sc_hd__a221o_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20966__A _20966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_61 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13641_ _13630_/A _13630_/B _13634_/X vssd1 vssd1 vccd1 vccd1 _13641_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22839_ _22839_/A _22839_/B vssd1 vssd1 vccd1 vccd1 _22840_/C sky130_fd_sc_hd__nor2_1
XANTENNA__18158__C1 _18001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18436__A _19279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16360_/A vssd1 vssd1 vccd1 vccd1 _16360_/X sky130_fd_sc_hd__buf_2
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _13709_/C _13712_/D _22278_/B _22566_/C vssd1 vssd1 vccd1 vccd1 _13573_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19370__A1 _12246_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15311_ _15311_/A _15311_/B _15311_/C vssd1 vssd1 vccd1 vccd1 _15348_/A sky130_fd_sc_hd__nand3_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12534_/A _12523_/B vssd1 vssd1 vccd1 vccd1 _12527_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11796__A2 _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16291_ _17974_/C vssd1 vssd1 vccd1 vccd1 _18172_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__16184__A1 _15932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18030_ _18030_/A vssd1 vssd1 vccd1 vccd1 _18032_/A sky130_fd_sc_hd__inv_2
X_15242_ _15096_/A _15096_/B _15310_/B _15305_/A _15010_/A vssd1 vssd1 vccd1 vccd1
+ _15242_/X sky130_fd_sc_hd__a32o_1
X_12454_ _19512_/C _19530_/D _18511_/A _12422_/D vssd1 vssd1 vccd1 vccd1 _12454_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_172_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15173_ _15095_/X _15170_/Y _15172_/Y vssd1 vssd1 vccd1 vccd1 _15173_/Y sky130_fd_sc_hd__o21ai_1
X_12385_ _12304_/X _12305_/Y _12370_/Y _12384_/Y vssd1 vssd1 vccd1 vccd1 _12398_/B
+ sky130_fd_sc_hd__o22a_1
X_14124_ _14124_/A vssd1 vssd1 vccd1 vccd1 _14124_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23206__A0 _14599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19981_ _19815_/B _19975_/A _19807_/X _19701_/B vssd1 vssd1 vccd1 vccd1 _20073_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_125_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1019 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18932_ _18932_/A _18932_/B vssd1 vssd1 vccd1 vccd1 _18932_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14055_ _14049_/Y _14911_/A _14760_/B _14054_/Y vssd1 vssd1 vccd1 vccd1 _14056_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_140_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21768__B1 _13816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16122__C _16314_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12650__C _20781_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ _20906_/A _20907_/A _20784_/C _20908_/A vssd1 vssd1 vccd1 vccd1 _13029_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18863_ _18863_/A _18863_/B vssd1 vssd1 vccd1 vccd1 _18875_/B sky130_fd_sc_hd__nor2_2
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17814_ _17705_/B _17814_/B _17814_/C vssd1 vssd1 vccd1 vccd1 _17817_/B sky130_fd_sc_hd__nand3b_1
XFILLER_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17841__D1 _17414_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18794_ _12130_/X _19184_/A _18806_/A vssd1 vssd1 vccd1 vccd1 _18802_/A sky130_fd_sc_hd__o21ai_1
XFILLER_48_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17745_ _16479_/X _18096_/A _17734_/Y vssd1 vssd1 vccd1 vccd1 _17745_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_130_1052 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14957_ _14957_/A _14957_/B vssd1 vssd1 vccd1 vccd1 _15065_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12276__A3 _11885_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17739__A2 _17980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18936__A1 _18755_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13908_ _14191_/A _14191_/B _13908_/C vssd1 vssd1 vccd1 vccd1 _13940_/B sky130_fd_sc_hd__nand3_1
X_17676_ _17705_/A _17705_/B _17677_/C vssd1 vssd1 vccd1 vccd1 _17680_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13481__C _22159_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14888_ _14756_/B _15000_/A _15004_/A vssd1 vssd1 vccd1 vccd1 _14893_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12378__B _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19415_ _19239_/X _19240_/Y _19256_/C vssd1 vssd1 vccd1 vccd1 _19415_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16627_ _16627_/A vssd1 vssd1 vccd1 vccd1 _16627_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ _13839_/A _13839_/B _13839_/C vssd1 vssd1 vccd1 vccd1 _13853_/A sky130_fd_sc_hd__nand3_1
XFILLER_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17888__C _19957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19346_ _19345_/A _19345_/B _19345_/C vssd1 vssd1 vccd1 vccd1 _19346_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_188_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16558_ _16558_/A _16558_/B vssd1 vssd1 vccd1 vccd1 _16558_/X sky130_fd_sc_hd__xor2_1
XANTENNA__12433__B1 _12100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18164__A2 _18163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15509_ _15508_/A _15533_/A _15508_/C vssd1 vssd1 vccd1 vccd1 _15509_/Y sky130_fd_sc_hd__a21oi_1
X_19277_ _19294_/C _19294_/D vssd1 vssd1 vccd1 vccd1 _19278_/C sky130_fd_sc_hd__nand2_1
XFILLER_31_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16489_ _16433_/X _16757_/D _16572_/B vssd1 vssd1 vccd1 vccd1 _16492_/A sky130_fd_sc_hd__a21boi_1
X_18228_ _18268_/A _18268_/B vssd1 vssd1 vccd1 vccd1 _18269_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18159_ _20271_/A vssd1 vssd1 vccd1 vccd1 _18324_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21170_ _21276_/A _21438_/A _20786_/Y _12674_/X vssd1 vssd1 vccd1 vccd1 _21187_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20121_ _19783_/X _19776_/X _20032_/A _20205_/A _20120_/X vssd1 vssd1 vccd1 vccd1
+ _20121_/X sky130_fd_sc_hd__o32a_1
XFILLER_132_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20052_ _20045_/Y _20048_/Y _20050_/Y vssd1 vssd1 vccd1 vccd1 _20056_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__17427__A1 _17228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17978__A2 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20982__A1 _20984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater130 _23343_/CLK vssd1 vssd1 vccd1 vccd1 _23378_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater141 _23441_/CLK vssd1 vssd1 vccd1 vccd1 _23442_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater152 _23432_/CLK vssd1 vssd1 vccd1 vccd1 _23398_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ _20966_/C vssd1 vssd1 vccd1 vccd1 _21302_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ _20885_/A _20885_/B vssd1 vssd1 vccd1 vccd1 _20885_/X sky130_fd_sc_hd__and2_1
XFILLER_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22624_ _22533_/X _22536_/B _22532_/Y _22530_/Y vssd1 vssd1 vccd1 vccd1 _22626_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_53_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1070 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22555_ _22656_/B _22790_/A _22757_/B _13465_/X vssd1 vssd1 vccd1 vccd1 _22556_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_194_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21506_ _21506_/A _21507_/B vssd1 vssd1 vccd1 vccd1 _21508_/A sky130_fd_sc_hd__or2_1
XFILLER_166_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22486_ _22057_/X _22168_/X _22636_/C _22392_/A vssd1 vssd1 vccd1 vccd1 _22486_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12727__A1 _12712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21437_ _20957_/X _21371_/Y _21434_/X _21436_/Y vssd1 vssd1 vccd1 vccd1 _21445_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_182_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19655__A2 _20080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12170_ _16856_/A vssd1 vssd1 vccd1 vccd1 _16122_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_108_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21368_ _21440_/C vssd1 vssd1 vccd1 vccd1 _21546_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_56 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11950__A2 _18434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23107_ _23107_/A vssd1 vssd1 vccd1 vccd1 _23379_/D sky130_fd_sc_hd__clkbuf_1
X_20319_ _20317_/X _20371_/C _20269_/C _20318_/X vssd1 vssd1 vccd1 vccd1 _20321_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_122_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21299_ _21299_/A vssd1 vssd1 vccd1 vccd1 _21455_/A sky130_fd_sc_hd__buf_2
XANTENNA__21214__A2 _21217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23038_ _23349_/Q input31/X _23038_/S vssd1 vssd1 vccd1 vccd1 _23039_/A sky130_fd_sc_hd__mux2_1
XANTENNA__19534__B _19534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_984 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13863__A _21832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15860_ _16821_/A _15868_/A _15860_/C _15860_/D vssd1 vssd1 vccd1 vccd1 _15985_/C
+ sky130_fd_sc_hd__and4_4
XFILLER_103_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15781__C _17066_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input21_A wb_dat_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14811_ _14228_/B _14816_/A _14218_/Y _14215_/Y vssd1 vssd1 vccd1 vccd1 _14811_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12479__A _18524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15791_ _15791_/A vssd1 vssd1 vccd1 vccd1 _15791_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12258__A3 _16364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22895__B _22895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22714__A2 _22392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _16994_/A _17210_/X _17524_/C _17524_/D vssd1 vssd1 vccd1 vccd1 _17530_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_57_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11954_ _11934_/Y _11937_/X _11938_/Y _11953_/X vssd1 vssd1 vccd1 vccd1 _11969_/A
+ sky130_fd_sc_hd__o211ai_4
X_14742_ _14734_/X _11860_/C _14738_/X vssd1 vssd1 vccd1 vccd1 _23265_/D sky130_fd_sc_hd__a21o_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17461_ _17610_/A _17465_/A _17454_/Y _17597_/A _17457_/Y vssd1 vssd1 vccd1 vccd1
+ _17473_/B sky130_fd_sc_hd__o221ai_4
X_14673_ _22896_/D vssd1 vssd1 vccd1 vccd1 _14673_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11885_ _11882_/X _11883_/X _11884_/Y _11784_/C vssd1 vssd1 vccd1 vccd1 _11885_/Y
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_189_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18166__A _19967_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19700__D _19700_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19200_ _11936_/X _19196_/B _19196_/C vssd1 vssd1 vccd1 vccd1 _19201_/C sky130_fd_sc_hd__o21ai_2
X_16412_ _19494_/D vssd1 vssd1 vccd1 vccd1 _17723_/C sky130_fd_sc_hd__clkbuf_2
X_13624_ _22292_/A _22293_/A vssd1 vssd1 vccd1 vccd1 _22484_/A sky130_fd_sc_hd__nand2_2
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22478__A1 _13547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17392_ _17392_/A _17392_/B _17549_/A vssd1 vssd1 vccd1 vccd1 _17393_/A sky130_fd_sc_hd__nand3_1
XFILLER_34_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19131_ _19133_/A _19133_/B _19391_/A _19354_/B vssd1 vssd1 vccd1 vccd1 _19409_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_186_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16343_ _16343_/A vssd1 vssd1 vccd1 vccd1 _16575_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13555_ _13555_/A _13555_/B vssd1 vssd1 vccd1 vccd1 _13555_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ _12506_/A _12506_/B vssd1 vssd1 vccd1 vccd1 _15868_/A sky130_fd_sc_hd__nand2_1
X_19062_ _19062_/A _19062_/B vssd1 vssd1 vccd1 vccd1 _19063_/C sky130_fd_sc_hd__nand2_1
Xrepeater99 _23507_/Q vssd1 vssd1 vccd1 vccd1 _15577_/A sky130_fd_sc_hd__clkbuf_1
X_16274_ _16106_/Y _16276_/A _16581_/A _16272_/Y _16273_/X vssd1 vssd1 vccd1 vccd1
+ _16988_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_145_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13486_ _13486_/A _13486_/B vssd1 vssd1 vccd1 vccd1 _13566_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18013_ _18013_/A _18013_/B _18013_/C _18013_/D vssd1 vssd1 vccd1 vccd1 _18014_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_139_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15225_ _15225_/A _15225_/B _15225_/C vssd1 vssd1 vccd1 vccd1 _15225_/X sky130_fd_sc_hd__and3_1
XFILLER_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12437_ _12119_/Y _12122_/Y _12131_/Y vssd1 vssd1 vccd1 vccd1 _12438_/C sky130_fd_sc_hd__a21o_1
XFILLER_148_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15156_ _15388_/C _15267_/B _15267_/C _15265_/A vssd1 vssd1 vccd1 vccd1 _15156_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_153_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12368_ _12368_/A _12368_/B vssd1 vssd1 vccd1 vccd1 _12368_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18854__B1 _12464_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _14107_/A vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__buf_2
X_19964_ _19674_/A _19667_/B _19943_/B _19850_/Y vssd1 vssd1 vccd1 vccd1 _19987_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15087_ _15488_/A _15231_/A _15082_/Y _15083_/X vssd1 vssd1 vccd1 vccd1 _15090_/B
+ sky130_fd_sc_hd__o211ai_1
X_12299_ _12364_/B _12364_/C _12364_/A vssd1 vssd1 vccd1 vccd1 _12300_/C sky130_fd_sc_hd__a21boi_1
XFILLER_80_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18915_ _18913_/X _18914_/Y _18728_/Y _18584_/Y _18568_/A vssd1 vssd1 vccd1 vccd1
+ _18915_/Y sky130_fd_sc_hd__a32oi_2
XFILLER_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14038_ _14312_/B _14262_/A _14777_/C vssd1 vssd1 vccd1 vccd1 _14116_/A sky130_fd_sc_hd__nand3_1
XFILLER_68_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19895_ _19725_/C _19725_/A _19725_/B _19730_/B vssd1 vssd1 vccd1 vccd1 _19896_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_122_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18846_ _18846_/A vssd1 vssd1 vccd1 vccd1 _18875_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__20964__A1 _20969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16632__A2 _15731_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21990__A _22236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18777_ _18773_/A _18773_/B _18775_/Y _18776_/X vssd1 vssd1 vccd1 vccd1 _18781_/B
+ sky130_fd_sc_hd__o2bb2ai_2
X_15989_ _15995_/A _15986_/A _16181_/B vssd1 vssd1 vccd1 vccd1 _15999_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__14643__A1 _22142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14643__B2 _23300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17728_ _19951_/D _17885_/A _17969_/D _19957_/A vssd1 vssd1 vccd1 vccd1 _17728_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13851__C1 _21987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1070 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17659_ _17667_/A _17666_/A _17666_/B vssd1 vssd1 vccd1 vccd1 _17661_/B sky130_fd_sc_hd__nand3_1
XANTENNA__15199__A2 _14015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23586__CLK _23588_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20670_ _20670_/A _20673_/A _20670_/C vssd1 vssd1 vccd1 vccd1 _20670_/X sky130_fd_sc_hd__and3_1
XFILLER_91_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16308__B _18481_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19329_ _19196_/C _19482_/A _19328_/Y vssd1 vssd1 vccd1 vccd1 _19335_/A sky130_fd_sc_hd__o21ai_1
XFILLER_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_902 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16027__C _16308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22340_ _22341_/C _22341_/B _22341_/A vssd1 vssd1 vccd1 vccd1 _22342_/A sky130_fd_sc_hd__a21oi_2
XFILLER_148_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_bq_clk_i clkbuf_3_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_192_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22271_ _22271_/A _22271_/B vssd1 vssd1 vccd1 vccd1 _22271_/Y sky130_fd_sc_hd__nand2_1
XFILLER_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22045__B _22045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21222_ _21221_/B _21221_/C _21221_/A vssd1 vssd1 vccd1 vccd1 _21232_/C sky130_fd_sc_hd__a21o_1
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21153_ _21153_/A _21153_/B vssd1 vssd1 vccd1 vccd1 _21153_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13386__C _22521_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16320__B2 _16382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20104_ _19966_/A _20151_/A _18335_/B _20369_/A _19985_/A vssd1 vssd1 vccd1 vccd1
+ _20106_/A sky130_fd_sc_hd__a41o_1
XANTENNA__13134__B2 _12785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16871__A2 _16315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21084_ _21084_/A _21212_/A _21084_/C vssd1 vssd1 vccd1 vccd1 _21097_/C sky130_fd_sc_hd__nand3_1
X_20035_ _20042_/B _20042_/A _20034_/Y vssd1 vssd1 vccd1 vccd1 _20035_/Y sky130_fd_sc_hd__a21oi_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12893__B1 _12899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19022__B1 _19021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20707__A1 _20775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ _22508_/C _21988_/A _21988_/B _21992_/A vssd1 vssd1 vccd1 vccd1 _21989_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16387__A1 _16462_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20937_ _20937_/A _20937_/B _20937_/C vssd1 vssd1 vccd1 vccd1 _20947_/B sky130_fd_sc_hd__nand3_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_595 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__A _11931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _19203_/A vssd1 vssd1 vccd1 vccd1 _11670_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__21124__B _21124_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20868_ _20868_/A _20868_/B vssd1 vssd1 vccd1 vccd1 _20872_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22607_ _22607_/A _22607_/B vssd1 vssd1 vccd1 vccd1 _22609_/B sky130_fd_sc_hd__nand2_1
XFILLER_169_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_954 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23587_ _23588_/CLK _23587_/D vssd1 vssd1 vccd1 vccd1 _23587_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18533__C1 _18755_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20799_ _20799_/A _21047_/C vssd1 vssd1 vccd1 vccd1 _20800_/B sky130_fd_sc_hd__nor2_1
XFILLER_139_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13340_ _13377_/A _13338_/X _13377_/D _13339_/X _13304_/X vssd1 vssd1 vccd1 vccd1
+ _13456_/B sky130_fd_sc_hd__a311o_2
XFILLER_194_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17887__A1 _11948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22538_ _22538_/A _22538_/B vssd1 vssd1 vccd1 vccd1 _22729_/A sky130_fd_sc_hd__nand2_1
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21778__C _21778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22236__A _22236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_957 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ _13226_/X _13224_/B _13355_/A _13233_/Y vssd1 vssd1 vccd1 vccd1 _13498_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22469_ _22569_/A _22553_/C _22569_/C vssd1 vssd1 vccd1 vccd1 _22469_/X sky130_fd_sc_hd__and3_2
XANTENNA__12762__A _23452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15010_ _15010_/A vssd1 vssd1 vccd1 vccd1 _15371_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__17639__A1 _16408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12222_ _12222_/A vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__buf_2
XANTENNA__13373__A1 _23325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14570__B1 _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11923__A2 _11921_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20643__B1 _12601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21986__A3 _21988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ _12153_/A vssd1 vssd1 vccd1 vccd1 _12217_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12084_ _15861_/A vssd1 vssd1 vccd1 vccd1 _12509_/A sky130_fd_sc_hd__buf_2
X_16961_ _16961_/A _16961_/B _16961_/C vssd1 vssd1 vccd1 vccd1 _16964_/B sky130_fd_sc_hd__nand3_2
XANTENNA__23459__CLK _23492_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21199__A1 _20509_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18700_ _18499_/A _18499_/C _18499_/B _18529_/B vssd1 vssd1 vccd1 vccd1 _18700_/Y
+ sky130_fd_sc_hd__a31oi_1
X_15912_ _16236_/A _16236_/B _16236_/C vssd1 vssd1 vccd1 vccd1 _16251_/A sky130_fd_sc_hd__nand3_2
X_19680_ _19668_/X _18000_/A _19482_/B _19482_/A vssd1 vssd1 vccd1 vccd1 _19680_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_1_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16892_ _16894_/A _16894_/B _16890_/X _16891_/X vssd1 vssd1 vccd1 vccd1 _16895_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_49_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_816 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18631_ _18788_/A vssd1 vssd1 vccd1 vccd1 _19805_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _15843_/A _15843_/B vssd1 vssd1 vccd1 vccd1 _15844_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14625__A1 _21902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14625__B2 _20894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19280__A _19280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18562_ _18562_/A _18562_/B _18562_/C vssd1 vssd1 vccd1 vccd1 _18562_/Y sky130_fd_sc_hd__nand3_1
XFILLER_18_743 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _12978_/Y _13106_/A _12985_/Y vssd1 vssd1 vccd1 vccd1 _20464_/D sky130_fd_sc_hd__o21a_4
X_15774_ _15774_/A vssd1 vssd1 vccd1 vccd1 _17409_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17513_ _17513_/A _17513_/B _17513_/C vssd1 vssd1 vccd1 vccd1 _17514_/C sky130_fd_sc_hd__nand3_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _16800_/D _16807_/B vssd1 vssd1 vccd1 vccd1 _14725_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _18670_/A _18670_/B _18458_/Y _18465_/X vssd1 vssd1 vccd1 vccd1 _18495_/B
+ sky130_fd_sc_hd__o211ai_1
X_11937_ _11766_/A _11935_/X _11815_/A _11936_/X vssd1 vssd1 vccd1 vccd1 _11937_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16378__B2 _16225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16409__A _18503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _17444_/A vssd1 vssd1 vccd1 vccd1 _18778_/B sky130_fd_sc_hd__buf_2
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14656_ _21047_/B vssd1 vssd1 vccd1 vccd1 _20902_/B sky130_fd_sc_hd__buf_6
X_11868_ _11868_/A vssd1 vssd1 vccd1 vccd1 _16464_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19316__A1 _19320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13607_ _23472_/Q vssd1 vssd1 vccd1 vccd1 _22024_/C sky130_fd_sc_hd__buf_2
X_17375_ _17535_/A _17536_/A _17698_/A _17698_/B vssd1 vssd1 vccd1 vccd1 _17379_/A
+ sky130_fd_sc_hd__o211ai_1
X_14587_ _23040_/D vssd1 vssd1 vccd1 vccd1 _14587_/X sky130_fd_sc_hd__clkbuf_2
X_11799_ _11896_/A vssd1 vssd1 vccd1 vccd1 _11799_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_186_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_976 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19114_ _12167_/X _12168_/X _17435_/X _17434_/X _17567_/X vssd1 vssd1 vccd1 vccd1
+ _19116_/C sky130_fd_sc_hd__o221a_2
XFILLER_192_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16326_ _16326_/A _16326_/B vssd1 vssd1 vccd1 vccd1 _16331_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15967__B _15998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13538_ _13538_/A _13538_/B vssd1 vssd1 vccd1 vccd1 _13538_/X sky130_fd_sc_hd__or2_1
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15889__B1 _15864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19045_ _19045_/A _19045_/B vssd1 vssd1 vccd1 vccd1 _19047_/B sky130_fd_sc_hd__nand2_2
X_13469_ _13469_/A vssd1 vssd1 vccd1 vccd1 _13470_/A sky130_fd_sc_hd__clkbuf_2
X_16257_ _16254_/A _16254_/B _16255_/X _16256_/Y vssd1 vssd1 vccd1 vccd1 _16258_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15208_ _15208_/A _15408_/A vssd1 vssd1 vccd1 vccd1 _15208_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16188_ _16191_/A vssd1 vssd1 vccd1 vccd1 _16667_/D sky130_fd_sc_hd__clkinv_2
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ _15140_/C _15140_/B _15138_/X vssd1 vssd1 vccd1 vccd1 _15141_/A sky130_fd_sc_hd__a21bo_1
XFILLER_82_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16798__B _16798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19947_ _19156_/B _19156_/A _18996_/C _18434_/A vssd1 vssd1 vccd1 vccd1 _19948_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22387__B1 _13527_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19878_ _19875_/Y _19876_/X _19877_/Y vssd1 vssd1 vccd1 vccd1 _19879_/C sky130_fd_sc_hd__o21ai_1
XFILLER_114_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17406__C _17753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16605__A2 _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11735__B _16364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18829_ _18455_/A _18461_/C _18453_/X _18639_/B _18804_/A vssd1 vssd1 vccd1 vccd1
+ _18830_/A sky130_fd_sc_hd__o311a_1
XFILLER_56_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19190__A _19190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21840_ _21840_/A _21840_/B vssd1 vssd1 vccd1 vccd1 _21847_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12627__B1 _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19555__A1 _19534_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21771_ _13642_/X _13431_/A _21783_/B vssd1 vssd1 vccd1 vccd1 _21771_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16319__A _16319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23510_ _23510_/CLK input46/X vssd1 vssd1 vccd1 vccd1 _23510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17030__A2 _16665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20722_ _20722_/A _20853_/B vssd1 vssd1 vccd1 vccd1 _20724_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15223__A _15298_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19307__A1 _12018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23441_ _23441_/CLK _23441_/D vssd1 vssd1 vccd1 vccd1 _23441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20653_ _20653_/A _20653_/B vssd1 vssd1 vccd1 vccd1 _20653_/Y sky130_fd_sc_hd__nand2_2
XFILLER_23_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23372_ _23372_/CLK _23372_/D vssd1 vssd1 vccd1 vccd1 _23372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15877__B _19363_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20584_ _20584_/A vssd1 vssd1 vccd1 vccd1 _20585_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22323_ _22323_/A _22323_/B _22323_/C vssd1 vssd1 vccd1 vccd1 _22324_/C sky130_fd_sc_hd__nand3_1
XFILLER_118_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16541__B2 _16558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16054__A _16054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22254_ _22252_/C _22252_/A _23274_/Q vssd1 vssd1 vccd1 vccd1 _22452_/A sky130_fd_sc_hd__a21oi_1
XFILLER_145_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21205_ _21267_/C _21206_/A _21207_/C vssd1 vssd1 vccd1 vccd1 _21208_/A sky130_fd_sc_hd__a21o_1
XFILLER_155_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22185_ _13339_/X _22141_/D _22142_/B _22144_/C _22028_/Y vssd1 vssd1 vccd1 vccd1
+ _22187_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21136_ _21123_/X _21129_/Y _21135_/Y vssd1 vssd1 vccd1 vccd1 _21241_/C sky130_fd_sc_hd__o21a_1
XFILLER_120_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1000 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11926__A _11926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21067_ _21063_/Y _21066_/Y _21062_/X vssd1 vssd1 vccd1 vccd1 _21069_/B sky130_fd_sc_hd__a21o_1
XFILLER_115_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12866__B1 _21065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16057__B1 _16056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12330__A2 _12324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20018_ _19894_/Y _19901_/X _20017_/X vssd1 vssd1 vccd1 vccd1 _20018_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14607__A1 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17035__D _18157_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14607__B2 _20481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17613__A _17613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12840_ _20962_/B vssd1 vssd1 vccd1 vccd1 _21193_/C sky130_fd_sc_hd__clkbuf_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_55 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12845_/A _12901_/A _12845_/B _12845_/C vssd1 vssd1 vccd1 vccd1 _12775_/C
+ sky130_fd_sc_hd__nand4_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21969_ _21981_/A _21981_/C _22117_/D vssd1 vssd1 vccd1 vccd1 _21970_/A sky130_fd_sc_hd__a21boi_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _16549_/A vssd1 vssd1 vccd1 vccd1 _16510_/C sky130_fd_sc_hd__clkbuf_4
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11798_/A _11798_/B vssd1 vssd1 vccd1 vccd1 _11726_/A sky130_fd_sc_hd__or2_1
X_15490_ _15488_/X _15489_/X _15446_/X _15447_/Y vssd1 vssd1 vccd1 vccd1 _15493_/C
+ sky130_fd_sc_hd__a211oi_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14441_ _14446_/A _14441_/B _14441_/C vssd1 vssd1 vccd1 vccd1 _14441_/Y sky130_fd_sc_hd__nand3b_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11848_/A vssd1 vssd1 vccd1 vccd1 _11654_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_187_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21105__A1 _21268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17160_ _16879_/A _16879_/B _16879_/C _16893_/B _16873_/C vssd1 vssd1 vccd1 vccd1
+ _17163_/A sky130_fd_sc_hd__a32o_1
X_14372_ _14790_/C vssd1 vssd1 vccd1 vccd1 _15195_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_70_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11584_ _11577_/Y _12173_/A _16856_/B vssd1 vssd1 vccd1 vccd1 _16593_/A sky130_fd_sc_hd__a21boi_4
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18163__B _18163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16111_ _17860_/A vssd1 vssd1 vccd1 vccd1 _18093_/A sky130_fd_sc_hd__buf_2
XFILLER_122_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13323_ _13344_/A vssd1 vssd1 vccd1 vccd1 _13323_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17091_ _16617_/X _17068_/A _16830_/X vssd1 vssd1 vccd1 vccd1 _17091_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13254_ _22022_/A _13344_/A _13260_/C vssd1 vssd1 vccd1 vccd1 _13660_/A sky130_fd_sc_hd__o21ai_4
X_16042_ _16089_/A _16089_/B _16089_/C vssd1 vssd1 vccd1 vccd1 _16326_/B sky130_fd_sc_hd__nand3_2
XFILLER_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12205_ _12205_/A _12205_/B vssd1 vssd1 vccd1 vccd1 _12531_/A sky130_fd_sc_hd__nand2_1
XANTENNA__20616__B1 _13202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185_ _20704_/B vssd1 vssd1 vccd1 vccd1 _20726_/D sky130_fd_sc_hd__clkbuf_2
X_19801_ _20013_/A _20013_/B _19040_/X _18097_/A vssd1 vssd1 vccd1 vccd1 _19802_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12136_ _12029_/B _12011_/X _12025_/X _12022_/X vssd1 vssd1 vccd1 vccd1 _12138_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_111_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17993_ _17982_/B _17982_/A _17988_/A vssd1 vssd1 vccd1 vccd1 _17994_/C sky130_fd_sc_hd__a21boi_1
XFILLER_151_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22369__B1 _22647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_80 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19732_ _19730_/A _19730_/B _19740_/A _19880_/A vssd1 vssd1 vccd1 vccd1 _19733_/C
+ sky130_fd_sc_hd__o211ai_2
X_12067_ _12327_/A vssd1 vssd1 vccd1 vccd1 _18778_/C sky130_fd_sc_hd__buf_2
X_16944_ _16944_/A vssd1 vssd1 vccd1 vccd1 _16944_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23030__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20919__A1 _21358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17226__C _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20919__B2 _21431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19663_ _19674_/C _19674_/A _17643_/A _19859_/A vssd1 vssd1 vccd1 vccd1 _19667_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16875_ _16893_/A _16893_/B _16873_/C vssd1 vssd1 vccd1 vccd1 _16875_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16599__A1 _16153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18993__C1 _19805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18614_ _12374_/A _18604_/X _18599_/A _18599_/B _18763_/A vssd1 vssd1 vccd1 vccd1
+ _18615_/C sky130_fd_sc_hd__o221ai_4
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12609__B1 _12608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15826_ _15716_/C _15686_/X _12020_/X _12018_/X _16591_/D vssd1 vssd1 vccd1 vccd1
+ _15827_/B sky130_fd_sc_hd__o221a_1
XFILLER_92_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19594_ _19571_/Y _19574_/X _19590_/Y vssd1 vssd1 vccd1 vccd1 _19598_/B sky130_fd_sc_hd__o21ai_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18545_ _18554_/A _18554_/B _18547_/C vssd1 vssd1 vccd1 vccd1 _18545_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_882 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _15757_/A _15757_/B vssd1 vssd1 vccd1 vccd1 _16612_/A sky130_fd_sc_hd__nand2_8
XANTENNA__20147__A2 _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12969_ _13151_/A _12785_/X _12815_/C _12968_/X vssd1 vssd1 vccd1 vccd1 _12972_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_61_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11571__A _23587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14708_ _23409_/Q _14693_/X _14698_/X _23441_/Q _14707_/X vssd1 vssd1 vccd1 vccd1
+ _14708_/X sky130_fd_sc_hd__a221o_2
X_18476_ _18476_/A vssd1 vssd1 vccd1 vccd1 _18476_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15688_ _15688_/A vssd1 vssd1 vccd1 vccd1 _15716_/C sky130_fd_sc_hd__buf_2
XFILLER_166_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17427_ _17228_/X _17236_/B _17406_/Y _17093_/Y vssd1 vssd1 vccd1 vccd1 _17485_/C
+ sky130_fd_sc_hd__a22oi_4
XANTENNA__23260__A _23260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15978__A _19017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14639_ _19156_/B _14544_/X _14575_/X _14631_/X _14638_/X vssd1 vssd1 vccd1 vccd1
+ _14639_/X sky130_fd_sc_hd__a221o_1
XFILLER_14_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17358_ _17361_/B _17358_/B vssd1 vssd1 vccd1 vccd1 _17359_/A sky130_fd_sc_hd__nand2_1
XFILLER_158_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18512__A2 _17627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12793__C1 _12667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16309_ _16309_/A _16309_/B vssd1 vssd1 vccd1 vccd1 _16310_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13498__A _13498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ _17291_/A _17291_/B _17290_/A _17297_/D vssd1 vssd1 vccd1 vccd1 _17289_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19028_ _11948_/X _11951_/X _19018_/X _19020_/Y _19548_/A vssd1 vssd1 vccd1 vccd1
+ _19029_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_118_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19301__A2_N _19179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11899__A1 _11670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1069 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23021__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22941_ _22941_/A vssd1 vssd1 vccd1 vccd1 _23305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21881__C _22521_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22872_ _23284_/Q _22872_/B vssd1 vssd1 vccd1 vccd1 _22874_/A sky130_fd_sc_hd__xor2_1
XFILLER_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21823_ _21811_/X _21812_/Y _21803_/Y _21806_/X vssd1 vssd1 vccd1 vccd1 _21824_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__17152__B _17152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21754_ _21754_/A _21754_/B _21754_/C vssd1 vssd1 vccd1 vccd1 _21755_/A sky130_fd_sc_hd__nand3_1
XFILLER_184_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11912__C _11912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16991__B _17218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20705_ _20553_/A _20702_/Y _20701_/X _20704_/Y vssd1 vssd1 vccd1 vccd1 _20705_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21685_ _21694_/A _21698_/B _21542_/X _21704_/A vssd1 vssd1 vccd1 vccd1 _21685_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23424_ _23424_/CLK _23424_/D vssd1 vssd1 vccd1 vccd1 _23424_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21638__A2 _21432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20636_ _20636_/A vssd1 vssd1 vccd1 vccd1 _20636_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_957 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23355_ _23358_/CLK _23355_/D vssd1 vssd1 vccd1 vccd1 _23355_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16514__A1 _16480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20567_ _20566_/C _20566_/A _20566_/B vssd1 vssd1 vccd1 vccd1 _20567_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16514__B2 _16479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22306_ _22135_/B _22128_/Y _22123_/Y _22126_/X vssd1 vssd1 vccd1 vccd1 _22405_/C
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_166_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23286_ _23297_/CLK _23286_/D vssd1 vssd1 vccd1 vccd1 _23286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20498_ _20498_/A _20498_/B vssd1 vssd1 vccd1 vccd1 _20782_/B sky130_fd_sc_hd__nand2_1
XFILLER_124_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22237_ _22237_/A vssd1 vssd1 vccd1 vccd1 _22237_/X sky130_fd_sc_hd__buf_2
XANTENNA__21453__A_N _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22168_ _22168_/A vssd1 vssd1 vccd1 vccd1 _22168_/X sky130_fd_sc_hd__buf_2
XFILLER_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21119_ _21119_/A _21119_/B _21119_/C vssd1 vssd1 vccd1 vccd1 _21134_/B sky130_fd_sc_hd__nand3_1
XANTENNA__23012__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12839__B1 _12770_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14990_ _14990_/A _14990_/B _15094_/C vssd1 vssd1 vccd1 vccd1 _14991_/A sky130_fd_sc_hd__nand3_1
XFILLER_8_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22099_ _22099_/A _22240_/A _22099_/C vssd1 vssd1 vccd1 vccd1 _22240_/B sky130_fd_sc_hd__nand3_2
XANTENNA__20969__A _20969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13941_ _23499_/Q vssd1 vssd1 vccd1 vccd1 _14096_/A sky130_fd_sc_hd__inv_2
XFILLER_86_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16660_ _17029_/A _16665_/A _17722_/A vssd1 vssd1 vccd1 vccd1 _16928_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__19261__C _19261_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13872_ _21732_/A vssd1 vssd1 vccd1 vccd1 _21971_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15611_ _15931_/A _15610_/X _15605_/A vssd1 vssd1 vccd1 vccd1 _15612_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__17062__B _17062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12823_ _20673_/A vssd1 vssd1 vccd1 vccd1 _20966_/C sky130_fd_sc_hd__clkbuf_2
X_16591_ _16591_/A _16591_/B _16591_/C _16591_/D vssd1 vssd1 vccd1 vccd1 _16592_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18330_ _18330_/A _18373_/A _20368_/B _18376_/B vssd1 vssd1 vccd1 vccd1 _18378_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15542_ _15508_/X _15513_/D _15540_/Y vssd1 vssd1 vccd1 vccd1 _15543_/B sky130_fd_sc_hd__o21ai_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12754_/A _13151_/C vssd1 vssd1 vccd1 vccd1 _12770_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18261_ _18204_/B _18204_/C _23532_/Q vssd1 vssd1 vccd1 vccd1 _18264_/A sky130_fd_sc_hd__a21bo_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _19363_/A _12024_/B _12105_/C vssd1 vssd1 vccd1 vccd1 _11705_/Y sky130_fd_sc_hd__nand3_2
X_15473_ _15474_/B _15474_/A vssd1 vssd1 vccd1 vccd1 _15475_/A sky130_fd_sc_hd__or2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12685_ _12677_/X _12704_/A _12696_/A _12851_/C vssd1 vssd1 vccd1 vccd1 _20509_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_187_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _17212_/A _23524_/Q _17212_/C vssd1 vssd1 vccd1 vccd1 _17381_/C sky130_fd_sc_hd__nand3_1
X_11636_ _16856_/A vssd1 vssd1 vccd1 vccd1 _16591_/A sky130_fd_sc_hd__buf_4
X_14424_ _14311_/X _14369_/X _14310_/Y _14423_/Y vssd1 vssd1 vccd1 vccd1 _14498_/A
+ sky130_fd_sc_hd__a31oi_1
X_18192_ _18192_/A _18194_/A vssd1 vssd1 vccd1 vccd1 _18192_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20209__A _20209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17143_ _16908_/A _17138_/A _17140_/Y vssd1 vssd1 vccd1 vccd1 _17150_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__16505__A1 _12238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15310__B _15310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14355_ _14355_/A _14407_/B _14355_/C vssd1 vssd1 vccd1 vccd1 _14355_/X sky130_fd_sc_hd__and3_1
XANTENNA__12653__C _20782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13306_ _13318_/C vssd1 vssd1 vccd1 vccd1 _21882_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_157_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17074_ _16814_/X _16821_/Y _16822_/X vssd1 vssd1 vccd1 vccd1 _17074_/X sky130_fd_sc_hd__a21o_1
XFILLER_116_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14286_ _14285_/B _14285_/C _14285_/A vssd1 vssd1 vccd1 vccd1 _14286_/X sky130_fd_sc_hd__a21o_1
XFILLER_170_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13237_ _23478_/Q vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__inv_2
X_16025_ _16021_/Y _16022_/Y _15895_/C _16347_/A _16347_/B vssd1 vssd1 vccd1 vccd1
+ _16108_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_171_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13168_ _13168_/A _13168_/B _13168_/C _13168_/D vssd1 vssd1 vccd1 vccd1 _13169_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_152_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11750__B1 _11741_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _12131_/A _12425_/A vssd1 vssd1 vccd1 vccd1 _12119_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__19207__B1 _11948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17976_ _17976_/A vssd1 vssd1 vccd1 vccd1 _20210_/A sky130_fd_sc_hd__buf_2
X_13099_ _13205_/C _13205_/A _13205_/B vssd1 vssd1 vccd1 vccd1 _13099_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19758__A1 _19554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19715_ _19717_/A _19717_/B _19723_/A _19723_/B vssd1 vssd1 vccd1 vccd1 _19719_/B
+ sky130_fd_sc_hd__o211ai_1
X_16927_ _16318_/C _17391_/B _17391_/C _16923_/C _16923_/B vssd1 vssd1 vccd1 vccd1
+ _16936_/B sky130_fd_sc_hd__a32o_1
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19646_ _16032_/X _16033_/X _18800_/A _18800_/B vssd1 vssd1 vccd1 vccd1 _19675_/A
+ sky130_fd_sc_hd__a2bb2oi_4
X_16858_ _16858_/A vssd1 vssd1 vccd1 vccd1 _17107_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15809_ _16225_/A _17409_/A _17465_/A _15800_/Y _15802_/Y vssd1 vssd1 vccd1 vccd1
+ _16019_/B sky130_fd_sc_hd__o221ai_4
X_19577_ _19577_/A _19577_/B _19577_/C vssd1 vssd1 vccd1 vccd1 _19577_/X sky130_fd_sc_hd__and3_1
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16789_ _17369_/B vssd1 vssd1 vccd1 vccd1 _17025_/A sky130_fd_sc_hd__buf_2
XFILLER_46_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18528_ _18499_/A _18499_/C _18499_/B vssd1 vssd1 vccd1 vccd1 _18528_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18459_ _12425_/X _12427_/X _12429_/Y _12441_/B vssd1 vssd1 vccd1 vccd1 _18464_/A
+ sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__15547__A2 _15525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21470_ _21472_/B _21472_/A vssd1 vssd1 vccd1 vccd1 _21474_/A sky130_fd_sc_hd__nand2_1
XFILLER_105_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20421_ _20418_/Y _20419_/X _20420_/Y _20394_/B vssd1 vssd1 vccd1 vccd1 _20423_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23140_ _23140_/A vssd1 vssd1 vccd1 vccd1 _23393_/D sky130_fd_sc_hd__clkbuf_1
X_20352_ _20352_/A _20352_/B vssd1 vssd1 vccd1 vccd1 _23534_/D sky130_fd_sc_hd__xor2_1
XFILLER_174_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23242__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23071_ _14632_/X input11/X _23073_/S vssd1 vssd1 vccd1 vccd1 _23072_/A sky130_fd_sc_hd__mux2_1
X_20283_ _20283_/A _20283_/B _20283_/C vssd1 vssd1 vccd1 vccd1 _20283_/Y sky130_fd_sc_hd__nor3_1
XFILLER_161_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22022_ _22022_/A _22141_/D vssd1 vssd1 vccd1 vccd1 _22022_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15890__B _15890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22924_ _22924_/A vssd1 vssd1 vccd1 vccd1 _23297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22855_ _22856_/B _22855_/B vssd1 vssd1 vccd1 vccd1 _23572_/D sky130_fd_sc_hd__xor2_4
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14994__B1 _14621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21806_ _21806_/A vssd1 vssd1 vccd1 vccd1 _21806_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22786_ _22786_/A _22786_/B vssd1 vssd1 vccd1 vccd1 _23570_/D sky130_fd_sc_hd__xor2_4
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_643 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18724__A2 _18723_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21737_ _23327_/Q _23326_/Q _23325_/Q vssd1 vssd1 vccd1 vccd1 _21901_/B sky130_fd_sc_hd__nor3_2
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12470_ _18531_/A _18506_/A _12461_/Y _12463_/Y vssd1 vssd1 vccd1 vccd1 _12473_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14746__B1 _14738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21668_ _21668_/A _21668_/B vssd1 vssd1 vccd1 vccd1 _21668_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23407_ _23409_/CLK _23407_/D vssd1 vssd1 vccd1 vccd1 _23407_/Q sky130_fd_sc_hd__dfxtp_1
X_20619_ _21070_/A _21054_/D _21035_/C _21036_/C vssd1 vssd1 vccd1 vccd1 _20619_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__22284__A2 _22059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21599_ _21556_/A _21556_/B _21555_/B vssd1 vssd1 vccd1 vccd1 _21599_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14140_ _14139_/A _14139_/B _14131_/A _14138_/A vssd1 vssd1 vccd1 vccd1 _14141_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23338_ _23339_/CLK _23338_/D vssd1 vssd1 vccd1 vccd1 _23338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14071_ _23359_/Q vssd1 vssd1 vccd1 vccd1 _14188_/A sky130_fd_sc_hd__buf_4
XANTENNA__23233__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23269_ _23584_/CLK _23269_/D vssd1 vssd1 vccd1 vccd1 _23269_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_153_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13022_ _12957_/Y _12674_/A _12714_/X _13018_/Y _13021_/Y vssd1 vssd1 vccd1 vccd1
+ _13022_/Y sky130_fd_sc_hd__o32ai_4
XFILLER_180_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input51_A x[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17057__B _17443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17830_ _17684_/X _17689_/X _17951_/D _17951_/A vssd1 vssd1 vccd1 vccd1 _17831_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18660__A1 _12245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17761_ _17761_/A _17761_/B vssd1 vssd1 vccd1 vccd1 _18604_/A sky130_fd_sc_hd__nand2_1
X_14973_ _23362_/Q _14868_/Y _15114_/B _23363_/Q vssd1 vssd1 vccd1 vccd1 _15171_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_47_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19500_ _16523_/A _16523_/B _19858_/A _20209_/A _12279_/A vssd1 vssd1 vccd1 vccd1
+ _19500_/X sky130_fd_sc_hd__o32a_1
XANTENNA__19703__D _19703_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16712_ _16712_/A _16712_/B vssd1 vssd1 vccd1 vccd1 _16956_/B sky130_fd_sc_hd__nor2_1
XANTENNA__18412__A1 _18277_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ _13927_/A _13946_/A _14124_/A vssd1 vssd1 vccd1 vccd1 _14173_/A sky130_fd_sc_hd__a21o_1
XFILLER_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17692_ _18058_/A _17945_/A vssd1 vssd1 vccd1 vccd1 _17693_/C sky130_fd_sc_hd__nand2_1
XANTENNA__15226__A1 _15538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19431_ _19431_/A vssd1 vssd1 vccd1 vccd1 _19431_/Y sky130_fd_sc_hd__inv_2
X_16643_ _16154_/Y _16157_/Y _16640_/X vssd1 vssd1 vccd1 vccd1 _16644_/A sky130_fd_sc_hd__a21oi_1
XFILLER_90_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13855_ _13676_/A _13676_/B _13676_/C _13692_/B _13692_/C vssd1 vssd1 vccd1 vccd1
+ _13856_/C sky130_fd_sc_hd__a32oi_1
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19362_ _19118_/Y _19119_/Y _19126_/X _19121_/A vssd1 vssd1 vccd1 vccd1 _19369_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_12806_ _13166_/A _20969_/A _12796_/X _12801_/Y _12805_/Y vssd1 vssd1 vccd1 vccd1
+ _12810_/A sky130_fd_sc_hd__o221ai_2
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16574_ _16294_/A _16575_/A _16575_/B vssd1 vssd1 vccd1 vccd1 _16755_/A sky130_fd_sc_hd__nand3b_2
XFILLER_34_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13786_ _23328_/Q vssd1 vssd1 vccd1 vccd1 _21738_/C sky130_fd_sc_hd__inv_2
XFILLER_76_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18313_ _18207_/X _18208_/X _18251_/A _18251_/B vssd1 vssd1 vccd1 vccd1 _18314_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_128_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15525_ _15525_/A _15525_/B vssd1 vssd1 vccd1 vccd1 _15525_/Y sky130_fd_sc_hd__nand2_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19293_ _19293_/A vssd1 vssd1 vccd1 vccd1 _19793_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12460__A1 _12184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12654_/Y _12661_/B _12652_/X _12651_/X vssd1 vssd1 vccd1 vccd1 _12738_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_128_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18244_/A _18245_/C vssd1 vssd1 vccd1 vccd1 _18293_/A sky130_fd_sc_hd__or2_2
XANTENNA__18335__C _18335_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14737__B1 _18435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1087 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15456_ _15457_/B _15457_/A vssd1 vssd1 vccd1 vccd1 _15458_/A sky130_fd_sc_hd__nand2_1
XANTENNA__21042__B _21174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12668_ _20495_/C vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__buf_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14407_ _14407_/A _14407_/B _14407_/C _14407_/D vssd1 vssd1 vccd1 vccd1 _14407_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_191_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18175_ _18172_/X _18094_/X _18170_/Y _18171_/X vssd1 vssd1 vccd1 vccd1 _18227_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_156_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11619_ _12167_/A _12168_/A vssd1 vssd1 vccd1 vccd1 _11815_/A sky130_fd_sc_hd__nor2_2
X_15387_ _15383_/X _15384_/Y _15386_/X vssd1 vssd1 vccd1 vccd1 _15403_/A sky130_fd_sc_hd__a21o_1
XFILLER_156_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12599_ _23449_/Q vssd1 vssd1 vccd1 vccd1 _20782_/C sky130_fd_sc_hd__buf_2
X_17126_ _17126_/A _17126_/B _17126_/C vssd1 vssd1 vccd1 vccd1 _17126_/X sky130_fd_sc_hd__and3_1
XFILLER_117_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14338_ _14353_/A _14353_/B _14353_/C vssd1 vssd1 vccd1 vccd1 _14403_/A sky130_fd_sc_hd__nand3_2
XFILLER_144_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15975__B _15975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17057_ _17057_/A _17443_/A _17444_/A vssd1 vssd1 vccd1 vccd1 _17058_/B sky130_fd_sc_hd__and3_1
XFILLER_116_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23224__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14269_ _14068_/X _14069_/X _14876_/B _14267_/Y _15195_/A vssd1 vssd1 vccd1 vccd1
+ _14269_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_125_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16008_ _16008_/A _16008_/B _16008_/C vssd1 vssd1 vccd1 vccd1 _16009_/A sky130_fd_sc_hd__nand3_1
XFILLER_135_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_855 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15991__A _15991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _17959_/A _17959_/B _20138_/A _20138_/B vssd1 vssd1 vccd1 vccd1 _17959_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20970_ _21356_/A _12648_/X _20967_/A vssd1 vssd1 vccd1 vccd1 _20974_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__17414__C _17414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_616 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16414__B1 _16469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19629_ _20031_/A _19916_/A _19916_/B _19916_/C vssd1 vssd1 vccd1 vccd1 _19633_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_38_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22640_ _22577_/B _22637_/Y _22646_/A _22703_/A vssd1 vssd1 vccd1 vccd1 _22641_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_198_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12436__D1 _16497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17509__A3 _18376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22571_ _22573_/A vssd1 vssd1 vccd1 vccd1 _22650_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21522_ _21570_/A _21522_/B vssd1 vssd1 vccd1 vccd1 _21524_/C sky130_fd_sc_hd__nor2_1
XFILLER_139_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15231__A _15231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17390__A1 _16529_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21453_ _21278_/A _21453_/B _21453_/C _21453_/D vssd1 vssd1 vccd1 vccd1 _21453_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20404_ _20366_/A _20314_/X _20368_/C _20368_/D _20373_/A vssd1 vssd1 vccd1 vccd1
+ _20405_/B sky130_fd_sc_hd__o41a_1
XFILLER_119_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1050 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21384_ _21191_/Y _21192_/Y _21307_/B _21307_/D vssd1 vssd1 vccd1 vccd1 _21386_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22064__A _22064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__B1 _11961_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23123_ _11784_/C input33/X _23123_/S vssd1 vssd1 vccd1 vccd1 _23124_/A sky130_fd_sc_hd__mux2_1
X_20335_ _20335_/A _20363_/B vssd1 vssd1 vccd1 vccd1 _20336_/B sky130_fd_sc_hd__nor2_1
XANTENNA__23215__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16496__A3 _15704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23054_ _14863_/A input34/X _23062_/S vssd1 vssd1 vccd1 vccd1 _23055_/A sky130_fd_sc_hd__mux2_1
X_20266_ _20317_/A _20215_/B _20215_/C _19425_/C _20146_/B vssd1 vssd1 vccd1 vccd1
+ _20268_/B sky130_fd_sc_hd__a32o_1
XFILLER_1_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput59 _14645_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[14] sky130_fd_sc_hd__buf_2
X_22005_ _22076_/B vssd1 vssd1 vccd1 vccd1 _22220_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18642__A1 _18476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20197_ _20206_/A _20252_/B _20196_/Y _20306_/A vssd1 vssd1 vccd1 vccd1 _20199_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23492__CLK _23492_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17605__B _17605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _12227_/B vssd1 vssd1 vccd1 vccd1 _12059_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22907_ _12601_/B input33/X _22907_/S vssd1 vssd1 vccd1 vccd1 _22908_/A sky130_fd_sc_hd__mux2_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20966__B _20966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13640_ _13639_/Y _13432_/Y _13460_/D _13474_/Y vssd1 vssd1 vccd1 vccd1 _13646_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_112_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22838_ _22800_/A _22861_/B _22792_/C _22797_/C _22836_/Y vssd1 vssd1 vccd1 vccd1
+ _22839_/B sky130_fd_sc_hd__a311oi_1
XANTENNA__18158__B1 _18376_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18436__B _19280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13571_ _22280_/B vssd1 vssd1 vccd1 vccd1 _22566_/C sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12442__A1 _12130_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22769_ _22718_/X _22767_/X _22789_/C vssd1 vssd1 vccd1 vccd1 _22770_/C sky130_fd_sc_hd__a21bo_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19370__A2 _12247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15310_ _15371_/B _15310_/B _15416_/A _15511_/D vssd1 vssd1 vccd1 vccd1 _15311_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_13_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12522_ _18559_/A _18559_/B _12522_/C vssd1 vssd1 vccd1 vccd1 _12523_/B sky130_fd_sc_hd__and3_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16290_ _17243_/B vssd1 vssd1 vccd1 vccd1 _17974_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16184__A2 _15933_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15241_ _15319_/C _15419_/B vssd1 vssd1 vccd1 vccd1 _15241_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19548__A _19548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12453_ _12123_/Y _12129_/Y _12217_/B _12217_/A vssd1 vssd1 vccd1 vccd1 _12484_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__14980__A _14980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12384_ _12384_/A _12384_/B _12383_/Y vssd1 vssd1 vccd1 vccd1 _12384_/Y sky130_fd_sc_hd__nor3b_2
X_15172_ _15001_/X _14999_/Y _15171_/Y vssd1 vssd1 vccd1 vccd1 _15172_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_181_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14123_ _14114_/X _14115_/Y _14133_/A vssd1 vssd1 vccd1 vccd1 _14130_/B sky130_fd_sc_hd__o21ai_1
X_19980_ _20212_/A _20146_/A _19980_/C _20058_/A vssd1 vssd1 vccd1 vccd1 _20073_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17684__A2 _18208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23206__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_874 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12931__C _20773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18931_ _18931_/A _18931_/B _19073_/A vssd1 vssd1 vccd1 vccd1 _18931_/X sky130_fd_sc_hd__and3_1
XFILLER_153_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14054_ _14054_/A _14054_/B vssd1 vssd1 vccd1 vccd1 _14054_/Y sky130_fd_sc_hd__nor2_1
XFILLER_180_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21768__B2 _22381_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14204__B _14246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13005_ _20473_/A _20782_/C _20473_/C _12695_/A _20781_/C vssd1 vssd1 vccd1 vccd1
+ _13005_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18862_ _18862_/A _18862_/B _18862_/C vssd1 vssd1 vccd1 vccd1 _18863_/B sky130_fd_sc_hd__and3_1
XANTENNA__16122__D _16314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17813_ _17673_/A _17673_/B _17814_/B _17814_/C vssd1 vssd1 vccd1 vccd1 _17817_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17841__C1 _18778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18793_ _18796_/A _18790_/X _18792_/Y vssd1 vssd1 vccd1 vccd1 _18806_/A sky130_fd_sc_hd__o21ai_1
XFILLER_95_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_bq_clk_i clkbuf_4_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _23462_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_48_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17744_ _17744_/A vssd1 vssd1 vccd1 vccd1 _18096_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14956_ _14956_/A vssd1 vssd1 vccd1 vccd1 _14959_/C sky130_fd_sc_hd__inv_2
XFILLER_78_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13907_ _23353_/Q vssd1 vssd1 vccd1 vccd1 _13908_/C sky130_fd_sc_hd__clkinv_2
XFILLER_35_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17675_ _17662_/Y _17669_/X _17671_/X _17674_/X vssd1 vssd1 vccd1 vccd1 _17705_/B
+ sky130_fd_sc_hd__o211ai_4
X_14887_ _14887_/A _14887_/B vssd1 vssd1 vccd1 vccd1 _15004_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19414_ _19437_/A vssd1 vssd1 vccd1 vccd1 _19428_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_51_906 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16626_ _17249_/A _17250_/A _16798_/B _16799_/A vssd1 vssd1 vccd1 vccd1 _16627_/A
+ sky130_fd_sc_hd__o211ai_4
X_13838_ _13820_/Y _13830_/Y _13834_/Y _13842_/B vssd1 vssd1 vccd1 vccd1 _13839_/C
+ sky130_fd_sc_hd__o211ai_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17888__D _18016_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19345_ _19345_/A _19345_/B _19345_/C vssd1 vssd1 vccd1 vccd1 _19345_/X sky130_fd_sc_hd__and3_1
XFILLER_16_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16557_ _16530_/A _16552_/Y _16530_/B vssd1 vssd1 vccd1 vccd1 _16558_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__12433__A1 _18435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13769_ _13769_/A vssd1 vssd1 vccd1 vccd1 _21880_/A sky130_fd_sc_hd__inv_2
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15508_ _15508_/A _15533_/A _15508_/C vssd1 vssd1 vccd1 vccd1 _15508_/X sky130_fd_sc_hd__and3_1
X_19276_ _18919_/X _19443_/B _19442_/A _19275_/Y _19442_/B vssd1 vssd1 vccd1 vccd1
+ _19294_/D sky130_fd_sc_hd__o2111ai_4
XANTENNA__21988__A _21988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16488_ _16488_/A vssd1 vssd1 vccd1 vccd1 _16757_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18227_ _18227_/A _18227_/B vssd1 vssd1 vccd1 vccd1 _18268_/B sky130_fd_sc_hd__nand2_1
XFILLER_148_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15439_ _15439_/A _15439_/B _15439_/C vssd1 vssd1 vccd1 vccd1 _15441_/A sky130_fd_sc_hd__and3_1
XFILLER_50_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18158_ _17889_/Y _18157_/B _18157_/Y _18376_/D _18001_/X vssd1 vssd1 vccd1 vccd1
+ _18187_/A sky130_fd_sc_hd__a311o_1
XANTENNA__21500__B _21548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17109_ _17118_/A _17118_/B _17112_/B _17112_/A vssd1 vssd1 vccd1 vccd1 _17109_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_18089_ _18088_/B _18088_/C _12088_/X _18211_/C vssd1 vssd1 vccd1 vccd1 _18090_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20120_ _20120_/A vssd1 vssd1 vccd1 vccd1 _20120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20051_ _20045_/Y _20048_/Y _20050_/Y _20268_/C _20215_/A vssd1 vssd1 vccd1 vccd1
+ _20054_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__19193__A _19327_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13953__B _14777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater120 _23391_/CLK vssd1 vssd1 vccd1 vccd1 _23396_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__20982__A2 _20984_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14110__A1 _14108_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater131 _23309_/CLK vssd1 vssd1 vccd1 vccd1 _23343_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater142 _23437_/CLK vssd1 vssd1 vccd1 vccd1 _23441_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater153 _23431_/CLK vssd1 vssd1 vccd1 vccd1 _23432_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_27_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20953_ _12675_/X _12704_/X _12711_/Y _12705_/X _21358_/C vssd1 vssd1 vccd1 vccd1
+ _20953_/X sky130_fd_sc_hd__o311a_1
XANTENNA__16938__A1 _16934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17596__D1 _17605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _20733_/Y _20717_/A _20846_/Y _20849_/Y vssd1 vssd1 vccd1 vccd1 _20884_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_939 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22623_ _22623_/A _22623_/B _22623_/C vssd1 vssd1 vccd1 vccd1 _22818_/B sky130_fd_sc_hd__nand3_1
XFILLER_107_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12585__A _23301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22554_ _22554_/A vssd1 vssd1 vccd1 vccd1 _22790_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18496__A1_N _18458_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21505_ _21554_/C _21554_/B vssd1 vssd1 vccd1 vccd1 _21507_/B sky130_fd_sc_hd__xnor2_2
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22485_ _22477_/Y _22479_/Y _22644_/A _22484_/X vssd1 vssd1 vccd1 vccd1 _22489_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_158_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21436_ _21435_/Y _21433_/Y _21431_/X vssd1 vssd1 vccd1 vccd1 _21436_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21998__A1 _21997_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21367_ _21377_/A _21377_/B _21377_/C vssd1 vssd1 vccd1 vccd1 _21378_/A sky130_fd_sc_hd__a21o_1
XFILLER_163_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20318_ _20265_/A _20366_/C _20365_/A _20265_/C vssd1 vssd1 vccd1 vccd1 _20318_/X
+ sky130_fd_sc_hd__o22a_1
X_23106_ _23379_/Q input28/X _23106_/S vssd1 vssd1 vccd1 vccd1 _23107_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_68 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21298_ _21173_/X _21298_/B _21298_/C vssd1 vssd1 vccd1 vccd1 _21306_/A sky130_fd_sc_hd__nand3b_1
XFILLER_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18076__C1 _18211_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23037_ _23037_/A vssd1 vssd1 vccd1 vccd1 _23348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13152__A2 _12709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20249_ _20246_/A _20248_/Y _20252_/C vssd1 vssd1 vccd1 vccd1 _20307_/C sky130_fd_sc_hd__o21ai_2
XFILLER_153_1031 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19534__C _19534_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16626__B1 _16798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_996 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15781__D _17062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _14814_/A _14814_/B _14814_/C vssd1 vssd1 vccd1 vccd1 _14810_/X sky130_fd_sc_hd__and3_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _15890_/A vssd1 vssd1 vccd1 vccd1 _15796_/B sky130_fd_sc_hd__inv_2
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A wb_dat_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22714__A3 _22392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ _14734_/X _11694_/X _14738_/X vssd1 vssd1 vccd1 vccd1 _23264_/D sky130_fd_sc_hd__a21o_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _11966_/A _11966_/B _11952_/Y vssd1 vssd1 vccd1 vccd1 _11953_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _17460_/A _17460_/B vssd1 vssd1 vccd1 vccd1 _17473_/A sky130_fd_sc_hd__nand2_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _14693_/A vssd1 vssd1 vccd1 vccd1 _14672_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_76 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11884_ _11676_/X _11980_/B _11840_/X vssd1 vssd1 vccd1 vccd1 _11884_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16411_ _19199_/D vssd1 vssd1 vccd1 vccd1 _19494_/D sky130_fd_sc_hd__buf_2
X_13623_ _21752_/B vssd1 vssd1 vccd1 vccd1 _22293_/A sky130_fd_sc_hd__clkbuf_2
X_17391_ _19653_/A _17391_/B _17391_/C vssd1 vssd1 vccd1 vccd1 _17392_/B sky130_fd_sc_hd__and3_1
XFILLER_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12495__A _12536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19130_ _19127_/X _19128_/Y _19129_/X vssd1 vssd1 vccd1 vccd1 _19354_/B sky130_fd_sc_hd__o21ai_2
X_16342_ _16337_/X _16104_/A _16340_/Y _16341_/X vssd1 vssd1 vccd1 vccd1 _16343_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_198_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _22474_/A _13553_/X _13490_/A vssd1 vssd1 vccd1 vccd1 _13554_/X sky130_fd_sc_hd__o21a_1
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19061_ _18879_/Y _18882_/Y _18884_/A _18884_/B vssd1 vssd1 vccd1 vccd1 _19062_/B
+ sky130_fd_sc_hd__o22ai_1
X_12505_ _12514_/B _23260_/B vssd1 vssd1 vccd1 vccd1 _12506_/B sky130_fd_sc_hd__nand2_1
XFILLER_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16273_ _16281_/C _16585_/A _16275_/A vssd1 vssd1 vccd1 vccd1 _16273_/X sky130_fd_sc_hd__a21o_1
X_13485_ _13485_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _21793_/A sky130_fd_sc_hd__nand2_1
X_18012_ _17032_/A _17032_/B _20081_/A _18007_/Y vssd1 vssd1 vccd1 vccd1 _18013_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_145_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15224_ _15455_/A vssd1 vssd1 vccd1 vccd1 _15225_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_157_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12436_ _12425_/X _12427_/X _12429_/Y _19703_/A _16497_/A vssd1 vssd1 vccd1 vccd1
+ _12438_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_138_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18303__B1 _18417_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15155_ _15155_/A vssd1 vssd1 vccd1 vccd1 _15388_/C sky130_fd_sc_hd__clkbuf_2
X_12367_ _12368_/A _12368_/B _12366_/Y vssd1 vssd1 vccd1 vccd1 _12384_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__18854__B2 _11961_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output82_A _14584_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14106_ _14029_/X _14015_/B _14312_/B vssd1 vssd1 vccd1 vccd1 _14107_/A sky130_fd_sc_hd__o21ai_1
X_19963_ _19963_/A _19963_/B vssd1 vssd1 vccd1 vccd1 _19996_/A sky130_fd_sc_hd__nor2_1
XFILLER_153_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12298_ _12298_/A _12298_/B _12298_/C vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__nand3_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15086_ _15082_/Y _15083_/X _15085_/X vssd1 vssd1 vccd1 vccd1 _15090_/A sky130_fd_sc_hd__a21o_1
XFILLER_45_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18914_ _18914_/A _18914_/B _18914_/C vssd1 vssd1 vccd1 vccd1 _18914_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__18606__A1 _11815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14037_ _14189_/A _14191_/C _14078_/A _14012_/A vssd1 vssd1 vccd1 vccd1 _14777_/C
+ sky130_fd_sc_hd__a31o_2
XFILLER_45_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19894_ _19894_/A _19894_/B _19894_/C vssd1 vssd1 vccd1 vccd1 _19894_/Y sky130_fd_sc_hd__nand3_2
XFILLER_68_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18845_ _18845_/A _18845_/B _18845_/C vssd1 vssd1 vccd1 vccd1 _18846_/A sky130_fd_sc_hd__nand3_1
XFILLER_80_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20964__A2 _12648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11574__A _23598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18776_ _18969_/A _18966_/A _18966_/B vssd1 vssd1 vccd1 vccd1 _18776_/X sky130_fd_sc_hd__and3_1
XFILLER_95_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15988_ _15858_/B _15969_/X _15993_/A vssd1 vssd1 vccd1 vccd1 _16181_/B sky130_fd_sc_hd__o21ai_1
X_17727_ _19949_/A vssd1 vssd1 vccd1 vccd1 _19957_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19031__A1 _18675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14939_ _14939_/A _14939_/B vssd1 vssd1 vccd1 vccd1 _14944_/B sky130_fd_sc_hd__nor2_2
XFILLER_82_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19031__B2 _19196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17899__C _18017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17042__B1 _15884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17261__A _18607_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17658_ _17658_/A _17658_/B _17658_/C vssd1 vssd1 vccd1 vccd1 _17666_/B sky130_fd_sc_hd__nand3_2
XFILLER_51_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_788 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23115__A0 _19261_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16609_ _16123_/A _16123_/B _17235_/A _17454_/B vssd1 vssd1 vccd1 vccd1 _16610_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17589_ _17974_/D _20138_/A _20138_/B _18077_/A _17974_/C vssd1 vssd1 vccd1 vccd1
+ _17589_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19328_ _16604_/A _12103_/X _19478_/A vssd1 vssd1 vccd1 vccd1 _19328_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16308__C _16308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18542__B1 _18721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19259_ _19259_/A _19259_/B _19259_/C vssd1 vssd1 vccd1 vccd1 _19297_/B sky130_fd_sc_hd__nand3_2
XANTENNA__16027__D _16027_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22270_ _22381_/A _22381_/B _22270_/C vssd1 vssd1 vccd1 vccd1 _22271_/B sky130_fd_sc_hd__nand3_1
XFILLER_145_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21221_ _21221_/A _21221_/B _21221_/C vssd1 vssd1 vccd1 vccd1 _21232_/B sky130_fd_sc_hd__nand3_1
XFILLER_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21152_ _20859_/Y _21004_/X _21151_/Y _21005_/Y vssd1 vssd1 vccd1 vccd1 _21152_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__22929__A0 _23300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20103_ _20102_/B _20177_/B _20103_/C vssd1 vssd1 vccd1 vccd1 _20106_/C sky130_fd_sc_hd__nand3b_2
XFILLER_132_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13964__A _14331_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21083_ _21083_/A _21083_/B vssd1 vssd1 vccd1 vccd1 _21083_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20034_ _20042_/B _20033_/Y _23549_/Q vssd1 vssd1 vccd1 vccd1 _20034_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A wb_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19270__B2 _19082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19651__A _19651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20797__A _23296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ _21983_/X _21893_/A _21984_/Y vssd1 vssd1 vccd1 vccd1 _21992_/A sky130_fd_sc_hd__o21ai_2
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23530__CLK _23558_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _12709_/A _21592_/A _20940_/C _20940_/A vssd1 vssd1 vccd1 vccd1 _20937_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__17584__A1 _16356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__B _11931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18417__D _18417_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20867_ _20867_/A _20867_/B vssd1 vssd1 vccd1 vccd1 _20868_/B sky130_fd_sc_hd__nand2_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22606_ _22601_/Y _22510_/X _22602_/Y vssd1 vssd1 vccd1 vccd1 _22606_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_179_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23586_ _23588_/CLK _23586_/D vssd1 vssd1 vccd1 vccd1 _23586_/Q sky130_fd_sc_hd__dfxtp_2
X_20798_ _20798_/A _20897_/C _20798_/C _20897_/D vssd1 vssd1 vccd1 vccd1 _21047_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_169_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18533__B1 _18755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_966 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17887__A2 _11951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22537_ _22538_/B _22525_/B _22523_/Y vssd1 vssd1 vccd1 vccd1 _22537_/X sky130_fd_sc_hd__a21o_1
XFILLER_168_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13270_ _21739_/A vssd1 vssd1 vccd1 vccd1 _13355_/A sky130_fd_sc_hd__clkbuf_2
X_22468_ _22468_/A vssd1 vssd1 vccd1 vccd1 _22468_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15362__A3 _15358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12221_ _12231_/A _12231_/B _12203_/Y _12220_/Y vssd1 vssd1 vccd1 vccd1 _18437_/D
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__14570__A1 _13911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17639__A2 _18002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21419_ _21409_/X _21413_/X _21418_/Y vssd1 vssd1 vccd1 vccd1 _21422_/A sky130_fd_sc_hd__o21a_1
XFILLER_151_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14570__B2 _14569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22399_ _22323_/C _22323_/B _22291_/Y vssd1 vssd1 vccd1 vccd1 _22401_/B sky130_fd_sc_hd__a21oi_1
XFILLER_191_980 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ _16437_/A _12324_/A _12093_/X _12151_/Y _12107_/A vssd1 vssd1 vccd1 vccd1
+ _12152_/X sky130_fd_sc_hd__o221a_1
XFILLER_68_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12083_ _18600_/A _18600_/B vssd1 vssd1 vccd1 vccd1 _15861_/A sky130_fd_sc_hd__nand2_2
X_16960_ _16954_/Y _17173_/B _16944_/X _17184_/A vssd1 vssd1 vccd1 vccd1 _16961_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_151_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21199__A2 _21190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15911_ _11868_/A _15797_/A _15899_/X _15910_/X _15902_/Y vssd1 vssd1 vccd1 vccd1
+ _16236_/C sky130_fd_sc_hd__o221ai_2
X_16891_ _16893_/A _16893_/B _16880_/X _16871_/X vssd1 vssd1 vccd1 vccd1 _16891_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18630_ _16194_/A _18461_/B _18460_/A _16360_/A _12103_/X vssd1 vssd1 vccd1 vccd1
+ _18630_/X sky130_fd_sc_hd__o32a_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _16591_/A _16591_/B _16612_/A vssd1 vssd1 vccd1 vccd1 _15843_/B sky130_fd_sc_hd__nand3_4
XFILLER_92_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15822__A1 _11882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _18549_/Y _18550_/X _18554_/C vssd1 vssd1 vccd1 vccd1 _18562_/C sky130_fd_sc_hd__o21ai_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15773_ _15650_/Y _15641_/Y _15772_/X vssd1 vssd1 vccd1 vccd1 _15773_/Y sky130_fd_sc_hd__a21oi_1
X_12985_ _12985_/A _13088_/B vssd1 vssd1 vccd1 vccd1 _12985_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__22699__A2 _22566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _17513_/A _17513_/B _17513_/C vssd1 vssd1 vccd1 vccd1 _17514_/B sky130_fd_sc_hd__a21o_1
XFILLER_40_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14724_ _23597_/Q vssd1 vssd1 vccd1 vccd1 _16807_/B sky130_fd_sc_hd__buf_2
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ _12323_/A _18474_/X _19670_/B _18481_/X _18473_/X vssd1 vssd1 vccd1 vccd1
+ _18670_/B sky130_fd_sc_hd__o311a_1
X_11936_ _11936_/A vssd1 vssd1 vccd1 vccd1 _11936_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17443_ _17443_/A vssd1 vssd1 vccd1 vccd1 _17581_/A sky130_fd_sc_hd__buf_2
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ _14655_/A vssd1 vssd1 vccd1 vccd1 _21047_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21034__C _21050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11867_ _12016_/A _12016_/B _11866_/Y vssd1 vssd1 vccd1 vccd1 _12032_/B sky130_fd_sc_hd__o21ai_2
XFILLER_159_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19316__A2 _19321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13606_ _21752_/A _21752_/B _23471_/Q vssd1 vssd1 vccd1 vccd1 _13615_/A sky130_fd_sc_hd__nand3_4
X_17374_ _17524_/C _17374_/B _17374_/C _17524_/D vssd1 vssd1 vccd1 vccd1 _17698_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14586_ _23421_/Q vssd1 vssd1 vccd1 vccd1 _15713_/C sky130_fd_sc_hd__buf_2
X_11798_ _11798_/A _11798_/B vssd1 vssd1 vccd1 vccd1 _11896_/A sky130_fd_sc_hd__nor2_2
X_19113_ _19381_/D _19694_/A _19113_/C _19262_/A vssd1 vssd1 vccd1 vccd1 _19116_/B
+ sky130_fd_sc_hd__nand4_1
X_16325_ _16396_/B _16397_/B _16324_/Y vssd1 vssd1 vccd1 vccd1 _16325_/X sky130_fd_sc_hd__a21o_1
X_13537_ _13537_/A _13755_/C vssd1 vssd1 vccd1 vccd1 _13540_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22871__A2 _22869_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15889__A1 _12222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19044_ _19044_/A vssd1 vssd1 vccd1 vccd1 _19047_/C sky130_fd_sc_hd__buf_2
XFILLER_173_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16256_ _16242_/A _16242_/B _16243_/A vssd1 vssd1 vccd1 vccd1 _16256_/Y sky130_fd_sc_hd__a21oi_2
X_13468_ _13465_/X _13284_/Y _21892_/A _13467_/X _13320_/X vssd1 vssd1 vccd1 vccd1
+ _13468_/X sky130_fd_sc_hd__o311a_1
XFILLER_173_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15207_ _15221_/A _15277_/B _15222_/A vssd1 vssd1 vccd1 vccd1 _15211_/B sky130_fd_sc_hd__nand3_1
XFILLER_173_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14561__A1 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__C1 _18755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ _12419_/A vssd1 vssd1 vccd1 vccd1 _19530_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_173_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_874 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16187_ _16187_/A _16187_/B _16187_/C _16667_/C vssd1 vssd1 vccd1 vccd1 _16658_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13399_ _13417_/A vssd1 vssd1 vccd1 vccd1 _21883_/C sky130_fd_sc_hd__buf_2
XFILLER_57_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23258__A _23260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15138_ _13985_/D _13972_/X _15044_/D _15408_/A _15041_/Y vssd1 vssd1 vccd1 vccd1
+ _15138_/X sky130_fd_sc_hd__a41o_1
XFILLER_114_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15105__A3 _14469_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16302__A2 _16140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18204__A_N _23532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16798__C _18947_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15069_ _15063_/Y _15066_/Y _15068_/X vssd1 vssd1 vccd1 vccd1 _15220_/B sky130_fd_sc_hd__a21oi_2
X_19946_ _18435_/A _18998_/D _23396_/Q _18996_/A vssd1 vssd1 vccd1 vccd1 _19948_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_87_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19877_ _20003_/A _19888_/D vssd1 vssd1 vccd1 vccd1 _19877_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__20398__B1 _20368_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17263__B1 _19543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17406__D _17753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23553__CLK _23558_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16605__A3 _17626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18828_ _18844_/C _18872_/B _18872_/A vssd1 vssd1 vccd1 vccd1 _18828_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_28_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19004__A1 _11822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18759_ _12324_/A _15861_/A _18598_/A vssd1 vssd1 vccd1 vccd1 _18759_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21770_ _21755_/X _21760_/X _21764_/X _21769_/X vssd1 vssd1 vccd1 vccd1 _21782_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20721_ _20853_/A _20854_/A vssd1 vssd1 vccd1 vccd1 _20722_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11850__A2 _11848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19307__A2 _12020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23440_ _23442_/CLK _23440_/D vssd1 vssd1 vccd1 vccd1 _23440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20652_ _20652_/A _20652_/B vssd1 vssd1 vccd1 vccd1 _20653_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1030 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23371_ _23372_/CLK _23371_/D vssd1 vssd1 vccd1 vccd1 _23371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20583_ _20583_/A _21387_/C vssd1 vssd1 vccd1 vccd1 _20583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16335__A _16335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22322_ _22288_/Y _22289_/Y _22290_/Y _22166_/Y vssd1 vssd1 vccd1 vccd1 _22323_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22253_ _22451_/A _22451_/B _22451_/C vssd1 vssd1 vccd1 vccd1 _22253_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16829__B1 _15855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21204_ _12785_/X _12862_/X _21194_/A _21062_/X _21203_/X vssd1 vssd1 vccd1 vccd1
+ _21207_/C sky130_fd_sc_hd__o32a_1
XFILLER_151_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22184_ _22040_/Y _22179_/Y _22151_/Y _22183_/Y vssd1 vssd1 vccd1 vccd1 _22184_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21135_ _21132_/Y _21153_/A _21153_/B vssd1 vssd1 vccd1 vccd1 _21135_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_133_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16070__A _17248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21066_ _21070_/A _21196_/A _21079_/A _21193_/C vssd1 vssd1 vccd1 vccd1 _21066_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_150_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16057__A1 _16054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20017_ _20017_/A _20017_/B _20017_/C vssd1 vssd1 vccd1 vccd1 _20017_/X sky130_fd_sc_hd__and3_1
XANTENNA__19381__A _19799_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17254__B1 _17057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20320__A _20320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _13179_/A _12770_/B _12770_/C _21054_/B vssd1 vssd1 vccd1 vccd1 _12845_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_161_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21968_ _21968_/A _21981_/C vssd1 vssd1 vccd1 vccd1 _22107_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11721_/A _11724_/A vssd1 vssd1 vccd1 vccd1 _11798_/B sky130_fd_sc_hd__nand2_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ _21358_/A _21358_/B _21050_/D _20918_/Y _21431_/B vssd1 vssd1 vccd1 vccd1
+ _20919_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21899_ _21905_/A vssd1 vssd1 vccd1 vccd1 _22562_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14439_/C _14442_/B _14438_/A _14438_/B vssd1 vssd1 vccd1 vccd1 _14441_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_35_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17309__A1 _16464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _16802_/A _12147_/A _15704_/B vssd1 vssd1 vccd1 vccd1 _11848_/A sky130_fd_sc_hd__o21ai_1
XFILLER_74_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21105__A2 _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14371_ _14459_/D _14407_/D vssd1 vssd1 vccd1 vccd1 _14371_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23569_ _23582_/CLK _23569_/D vssd1 vssd1 vccd1 vccd1 _23569_/Q sky130_fd_sc_hd__dfxtp_1
X_11583_ _11637_/A vssd1 vssd1 vccd1 vccd1 _16856_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_11_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16110_ _16549_/B vssd1 vssd1 vccd1 vccd1 _17035_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13322_ _13228_/X _13226_/X _13523_/A _13483_/C _13260_/C vssd1 vssd1 vccd1 vccd1
+ _13325_/A sky130_fd_sc_hd__o311ai_1
XFILLER_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17090_ _17126_/A _17126_/B _17126_/C vssd1 vssd1 vccd1 vccd1 _17298_/A sky130_fd_sc_hd__nand3_1
XFILLER_109_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_852 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16041_ _12040_/X _16035_/X _16309_/A _16310_/B vssd1 vssd1 vccd1 vccd1 _16089_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_171_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13253_ _13253_/A vssd1 vssd1 vccd1 vccd1 _13260_/C sky130_fd_sc_hd__clkinv_2
XFILLER_170_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12204_ _12387_/A _12204_/B vssd1 vssd1 vccd1 vccd1 _12205_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13184_ _13184_/A vssd1 vssd1 vccd1 vccd1 _20704_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19800_ _19900_/D _20013_/B _19800_/C _20013_/A vssd1 vssd1 vccd1 vccd1 _19802_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_124_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ _12130_/X _18645_/A _12131_/Y _12134_/Y vssd1 vssd1 vccd1 vccd1 _12138_/A
+ sky130_fd_sc_hd__o22ai_1
X_17992_ _17992_/A _17992_/B _17992_/C vssd1 vssd1 vccd1 vccd1 _18085_/A sky130_fd_sc_hd__nand3_2
XFILLER_124_888 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19731_ _19731_/A _19731_/B vssd1 vssd1 vccd1 vccd1 _19733_/B sky130_fd_sc_hd__nand2_1
X_16943_ _16953_/A _17173_/A _16941_/Y _16942_/X vssd1 vssd1 vccd1 vccd1 _16944_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_92 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12066_ _12066_/A vssd1 vssd1 vccd1 vccd1 _12327_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17226__D _17226_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16048__A1 _11792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20919__A2 _21358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19662_ _19662_/A _20142_/C _19662_/C vssd1 vssd1 vccd1 vccd1 _19674_/A sky130_fd_sc_hd__nand3_2
X_16874_ _16890_/B vssd1 vssd1 vccd1 vccd1 _16893_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19942__B1_N _19888_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18993__B1 _18439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18613_ _12260_/D _19364_/B _17595_/A _19123_/B _12475_/B vssd1 vssd1 vccd1 vccd1
+ _18763_/A sky130_fd_sc_hd__a32o_1
X_15825_ _15813_/A _15709_/A _15785_/A vssd1 vssd1 vccd1 vccd1 _15827_/A sky130_fd_sc_hd__o21ai_1
XFILLER_93_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19593_ _19402_/Y _19398_/B _19401_/A vssd1 vssd1 vccd1 vccd1 _19598_/A sky130_fd_sc_hd__a21boi_2
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11852__A _11852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18544_ _18902_/B _18553_/B vssd1 vssd1 vccd1 vccd1 _18547_/C sky130_fd_sc_hd__or2_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15756_ _15729_/X _15761_/A _15762_/A vssd1 vssd1 vccd1 vccd1 _15757_/B sky130_fd_sc_hd__o21ai_2
XFILLER_79_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12968_ _20563_/A _20563_/B _21358_/C _21295_/B _13158_/A vssd1 vssd1 vccd1 vccd1
+ _12968_/X sky130_fd_sc_hd__a32o_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12667__B _12667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11571__B _23588_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ _23377_/Q _14688_/X _14706_/X vssd1 vssd1 vccd1 vccd1 _14707_/X sky130_fd_sc_hd__o21a_1
X_11919_ _11959_/A vssd1 vssd1 vccd1 vccd1 _11947_/A sky130_fd_sc_hd__buf_2
X_18475_ _18475_/A vssd1 vssd1 vccd1 vccd1 _18476_/A sky130_fd_sc_hd__buf_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ _23420_/Q _23429_/Q vssd1 vssd1 vccd1 vccd1 _15688_/A sky130_fd_sc_hd__nand2_1
X_12899_ _12899_/A _12899_/B _12899_/C vssd1 vssd1 vccd1 vccd1 _13044_/B sky130_fd_sc_hd__nand3_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _17426_/A _17426_/B _17426_/C vssd1 vssd1 vccd1 vccd1 _17485_/B sky130_fd_sc_hd__nand3_1
X_14638_ _14632_/X _14635_/X _14637_/X vssd1 vssd1 vccd1 vccd1 _14638_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15978__B _16314_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17357_ _17357_/A _17357_/B vssd1 vssd1 vccd1 vccd1 _17357_/Y sky130_fd_sc_hd__nand2_2
XFILLER_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14569_ _23418_/Q vssd1 vssd1 vccd1 vccd1 _14569_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ _16674_/A _18481_/C _16308_/C _16308_/D vssd1 vssd1 vccd1 vccd1 _16309_/B
+ sky130_fd_sc_hd__nand4_4
X_17288_ _17277_/Y _17281_/Y _17282_/Y _17287_/Y vssd1 vssd1 vccd1 vccd1 _17297_/D
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13498__B _13498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17720__A1 _12237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19027_ _19548_/A _19485_/A _19018_/A _19020_/Y vssd1 vssd1 vccd1 vccd1 _19029_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13337__A2 _22028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16239_ _16246_/C _16725_/A _16253_/B vssd1 vssd1 vccd1 vccd1 _16239_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11899__A2 _11898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21280__A1 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19929_ _19929_/A _19929_/B vssd1 vssd1 vccd1 vccd1 _19929_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22940_ _23305_/Q input17/X _22940_/S vssd1 vssd1 vccd1 vccd1 _22941_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17787__A1 _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22871_ _22887_/C _22869_/Y _22878_/A vssd1 vssd1 vccd1 vccd1 _22872_/B sky130_fd_sc_hd__a21boi_1
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21822_ _21803_/Y _21806_/X _21809_/Y vssd1 vssd1 vccd1 vccd1 _21824_/A sky130_fd_sc_hd__a21o_1
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16049__B _17414_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21753_ _21753_/A _21753_/B vssd1 vssd1 vccd1 vccd1 _21754_/C sky130_fd_sc_hd__nand2_1
XFILLER_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16211__A1 _11766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20704_ _23457_/Q _20704_/B vssd1 vssd1 vccd1 vccd1 _20704_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21684_ _21542_/X _21704_/A _21698_/B vssd1 vssd1 vccd1 vccd1 _21684_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__23449__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13689__A _22508_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23423_ _23427_/CLK _23423_/D vssd1 vssd1 vccd1 vccd1 _23423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20635_ _20635_/A _20635_/B _20635_/C vssd1 vssd1 vccd1 vccd1 _20636_/A sky130_fd_sc_hd__nand3_1
XFILLER_138_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15970__B1 _15860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16065__A _19196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21638__A3 _21432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12593__A _23301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20566_ _20566_/A _20566_/B _20566_/C vssd1 vssd1 vccd1 vccd1 _20566_/X sky130_fd_sc_hd__and3_1
X_23354_ _23365_/CLK _23354_/D vssd1 vssd1 vccd1 vccd1 _23354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16514__A2 _15698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21121__D _21554_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22048__B1 _14614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22305_ _22167_/C _22279_/A _22174_/Y _22300_/Y _22301_/Y vssd1 vssd1 vccd1 vccd1
+ _22405_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_166_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20497_ _20495_/C _23296_/Q _23297_/Q vssd1 vssd1 vccd1 vccd1 _20498_/B sky130_fd_sc_hd__a21oi_1
X_23285_ _23571_/CLK _23285_/D vssd1 vssd1 vccd1 vccd1 _23285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19464__A1 _19116_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22236_ _22236_/A vssd1 vssd1 vccd1 vccd1 _22237_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15716__A_N _15713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22167_ _22380_/C _22479_/B _22167_/C vssd1 vssd1 vccd1 vccd1 _22167_/X sky130_fd_sc_hd__and3_1
XFILLER_191_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21118_ _20980_/A _21111_/Y _20981_/Y vssd1 vssd1 vccd1 vccd1 _21119_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__19216__A1 _19021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22098_ _22099_/A _22240_/A _22099_/C vssd1 vssd1 vccd1 vccd1 _22102_/A sky130_fd_sc_hd__a21o_1
XFILLER_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13940_ _13911_/C _13940_/B _14091_/A vssd1 vssd1 vccd1 vccd1 _13994_/B sky130_fd_sc_hd__nand3b_2
X_21049_ _20940_/C _21174_/B _21181_/A _20929_/Y vssd1 vssd1 vccd1 vccd1 _21053_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13871_ _21857_/A _13867_/Y _13870_/Y vssd1 vssd1 vccd1 vccd1 _21732_/A sky130_fd_sc_hd__a21o_1
XFILLER_74_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15610_ _16683_/A vssd1 vssd1 vccd1 vccd1 _15610_/X sky130_fd_sc_hd__clkbuf_4
X_12822_ _23455_/Q vssd1 vssd1 vccd1 vccd1 _20673_/A sky130_fd_sc_hd__clkbuf_2
X_16590_ _16590_/A _16590_/B vssd1 vssd1 vccd1 vccd1 _16597_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17062__C _17761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15541_ _15225_/B _15538_/D _15508_/C _15513_/D _15540_/Y vssd1 vssd1 vccd1 vccd1
+ _15543_/A sky130_fd_sc_hd__a311o_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_83 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12753_ _12929_/A _20663_/C _12930_/A vssd1 vssd1 vccd1 vccd1 _13151_/C sky130_fd_sc_hd__nand3_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18455__A _18455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _18319_/A _18319_/B vssd1 vssd1 vccd1 vccd1 _18265_/A sky130_fd_sc_hd__nand2_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11704_ _11704_/A _11704_/B vssd1 vssd1 vccd1 vccd1 _11820_/A sky130_fd_sc_hd__nand2_2
X_15472_ _15472_/A _15501_/B vssd1 vssd1 vccd1 vccd1 _15474_/A sky130_fd_sc_hd__nand2_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12684_ _12577_/A _12682_/Y _12580_/A _12683_/Y vssd1 vssd1 vccd1 vccd1 _12851_/C
+ sky130_fd_sc_hd__a31o_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _16994_/A _17210_/X _17524_/C _17524_/D _17376_/A vssd1 vssd1 vccd1 vccd1
+ _17212_/C sky130_fd_sc_hd__o2111ai_1
XANTENNA__23511__D input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14495_/A _14495_/B _14495_/C _14495_/D vssd1 vssd1 vccd1 vccd1 _14423_/Y
+ sky130_fd_sc_hd__a22oi_1
X_18191_ _18191_/A _18191_/B vssd1 vssd1 vccd1 vccd1 _18194_/A sky130_fd_sc_hd__nand2_2
X_11635_ _11723_/A _11593_/C _11633_/Y _11634_/Y vssd1 vssd1 vccd1 vccd1 _16856_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_128_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17142_ _17142_/A vssd1 vssd1 vccd1 vccd1 _17635_/A sky130_fd_sc_hd__buf_2
XFILLER_7_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14354_ _14344_/B _14407_/C _14355_/A vssd1 vssd1 vccd1 vccd1 _14354_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13305_ _23322_/Q _13483_/B _21739_/A _13304_/X vssd1 vssd1 vccd1 vccd1 _13318_/C
+ sky130_fd_sc_hd__o211ai_2
X_17073_ _17073_/A _17073_/B vssd1 vssd1 vccd1 vccd1 _17073_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14285_ _14285_/A _14285_/B _14285_/C vssd1 vssd1 vccd1 vccd1 _14285_/Y sky130_fd_sc_hd__nand3_1
XFILLER_155_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_736 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16024_ _16347_/A _16347_/B _16347_/C vssd1 vssd1 vccd1 vccd1 _16108_/B sky130_fd_sc_hd__a21bo_1
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13236_ _23477_/Q vssd1 vssd1 vccd1 vccd1 _21997_/A sky130_fd_sc_hd__inv_2
XFILLER_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11847__A _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18663__C1 _18959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ _20563_/A _13181_/C _20563_/B _21279_/D vssd1 vssd1 vccd1 vccd1 _13168_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11750__A1 _11738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19207__A1 _18435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12118_ _12118_/A _18445_/B _12118_/C vssd1 vssd1 vccd1 vccd1 _12425_/A sky130_fd_sc_hd__nand3_2
XANTENNA__19207__B2 _11951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17975_ _17975_/A vssd1 vssd1 vccd1 vccd1 _17976_/A sky130_fd_sc_hd__clkbuf_2
X_13098_ _13203_/A _21554_/D _20583_/A vssd1 vssd1 vccd1 vccd1 _13205_/B sky130_fd_sc_hd__and3_1
X_19714_ _19716_/B vssd1 vssd1 vccd1 vccd1 _19723_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__19758__A2 _19534_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16926_ _17133_/B vssd1 vssd1 vccd1 vccd1 _17391_/C sky130_fd_sc_hd__clkbuf_2
X_12049_ _12049_/A _12049_/B vssd1 vssd1 vccd1 vccd1 _12057_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15892__A1_N _15889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1084 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19645_ _19504_/X _19505_/X _19648_/A _19502_/A vssd1 vssd1 vccd1 vccd1 _19667_/D
+ sky130_fd_sc_hd__o211a_2
X_16857_ _15691_/A _11924_/A _16856_/Y vssd1 vssd1 vccd1 vccd1 _16858_/A sky130_fd_sc_hd__o21ai_1
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15054__A _15054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15808_ _15808_/A _16318_/C _17860_/A vssd1 vssd1 vccd1 vccd1 _16019_/A sky130_fd_sc_hd__nand3_2
XFILLER_19_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19576_ _19522_/A _19521_/B _19577_/C vssd1 vssd1 vccd1 vccd1 _19576_/Y sky130_fd_sc_hd__a21oi_1
X_16788_ _16988_/A _17026_/B _16778_/A vssd1 vssd1 vccd1 vccd1 _17369_/B sky130_fd_sc_hd__a21oi_2
XFILLER_19_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18527_ _18519_/Y _18523_/Y _18526_/Y vssd1 vssd1 vccd1 vccd1 _18554_/A sky130_fd_sc_hd__a21o_1
X_15739_ _15862_/A _15862_/B _16122_/A _16122_/B vssd1 vssd1 vccd1 vccd1 _15852_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18458_ _18458_/A _18458_/B _18458_/C vssd1 vssd1 vccd1 vccd1 _18458_/Y sky130_fd_sc_hd__nand3_2
XFILLER_33_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17409_ _17409_/A vssd1 vssd1 vccd1 vccd1 _17644_/A sky130_fd_sc_hd__clkbuf_2
X_18389_ _18388_/A _18388_/B _18413_/A _18388_/D vssd1 vssd1 vccd1 vccd1 _18392_/B
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__15952__B1 _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_880 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20420_ _20420_/A _20420_/B vssd1 vssd1 vccd1 vccd1 _20420_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20351_ _20313_/A _20313_/B _20359_/A vssd1 vssd1 vccd1 vccd1 _20352_/B sky130_fd_sc_hd__o21a_1
XANTENNA__19196__A _19196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_991 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23070_ _23070_/A vssd1 vssd1 vccd1 vccd1 _23362_/D sky130_fd_sc_hd__clkbuf_1
X_20282_ _20279_/X _20280_/Y _20264_/X _20231_/C vssd1 vssd1 vccd1 vccd1 _20282_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_134_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22021_ _22021_/A vssd1 vssd1 vccd1 vccd1 _22141_/D sky130_fd_sc_hd__buf_2
XFILLER_1_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17444__A _17444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12151__D1 _19700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22753__A1 _22713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18259__B _23533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21363__B1_N _21285_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22923_ _14615_/X input9/X _22929_/S vssd1 vssd1 vccd1 vccd1 _22924_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22854_ _22856_/C _22854_/B vssd1 vssd1 vccd1 vccd1 _22855_/B sky130_fd_sc_hd__nand2_1
XFILLER_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23271__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21805_ _21805_/A _21805_/B _21805_/C vssd1 vssd1 vccd1 vccd1 _21806_/A sky130_fd_sc_hd__nand3_1
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22785_ _22747_/A _22747_/B _22821_/B vssd1 vssd1 vccd1 vccd1 _22786_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__12100__B _12100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19382__B1 _19361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21736_ _21745_/B _21898_/B _21898_/C vssd1 vssd1 vccd1 vccd1 _22033_/A sky130_fd_sc_hd__nand3b_2
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14746__A1 _11633_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21667_ _21643_/A _21642_/A _21642_/B vssd1 vssd1 vccd1 vccd1 _21671_/B sky130_fd_sc_hd__a21boi_1
XFILLER_8_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23406_ _23409_/CLK _23406_/D vssd1 vssd1 vccd1 vccd1 _23406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20618_ _20728_/A _20713_/B _20714_/A vssd1 vssd1 vccd1 vccd1 _20618_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21598_ _21598_/A _21641_/B vssd1 vssd1 vccd1 vccd1 _21602_/B sky130_fd_sc_hd__xor2_2
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23337_ _23445_/CLK _23337_/D vssd1 vssd1 vccd1 vccd1 _23337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20549_ _20553_/A _20553_/B _20547_/C vssd1 vssd1 vccd1 vccd1 _20549_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16523__A _16523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14070_ _14124_/A vssd1 vssd1 vccd1 vccd1 _14070_/X sky130_fd_sc_hd__buf_4
XFILLER_118_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_630 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23268_ _23584_/CLK _23268_/D vssd1 vssd1 vccd1 vccd1 _23268_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_152_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13021_ _13019_/Y _12668_/X _20481_/B vssd1 vssd1 vccd1 vccd1 _13021_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22219_ _22508_/C _22263_/B _22220_/D _22220_/A vssd1 vssd1 vccd1 vccd1 _22221_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_161_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17057__C _17444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23199_ _23199_/A vssd1 vssd1 vccd1 vccd1 _23419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input44_A x[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16120__B1 _15998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18660__A2 _11784_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17760_ _17760_/A _17760_/B vssd1 vssd1 vccd1 vccd1 _17760_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14972_ _15171_/A vssd1 vssd1 vccd1 vccd1 _15316_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18169__B _20151_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13923_ _23358_/Q vssd1 vssd1 vccd1 vccd1 _14124_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16711_ _16183_/X _16193_/Y _16199_/Y _16233_/B vssd1 vssd1 vccd1 vccd1 _16712_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18412__A2 _20317_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17691_ _17935_/D vssd1 vssd1 vccd1 vccd1 _18058_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12498__A _23591_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19430_ _19434_/C _19434_/A _19434_/B vssd1 vssd1 vccd1 vccd1 _19430_/Y sky130_fd_sc_hd__a21oi_1
X_16642_ _16853_/A _16649_/B _16640_/X _16641_/Y vssd1 vssd1 vccd1 vccd1 _16655_/D
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13854_ _13853_/A _13853_/B _13857_/A _13857_/B vssd1 vssd1 vccd1 vccd1 _13856_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__14434__B1 _14867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22076__A_N _22218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ _12815_/C _12805_/B vssd1 vssd1 vccd1 vccd1 _12805_/Y sky130_fd_sc_hd__nand2_1
X_19361_ _19361_/A _19361_/B vssd1 vssd1 vccd1 vccd1 _19376_/A sky130_fd_sc_hd__xor2_2
X_16573_ _16573_/A vssd1 vssd1 vccd1 vccd1 _16573_/Y sky130_fd_sc_hd__inv_2
X_13785_ _21744_/A _23324_/Q _13785_/C vssd1 vssd1 vccd1 vccd1 _22141_/A sky130_fd_sc_hd__nor3_2
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18312_ _18296_/X _18295_/X _18267_/Y _18301_/B vssd1 vssd1 vccd1 vccd1 _18314_/B
+ sky130_fd_sc_hd__a211o_1
X_15524_ _15525_/B _15525_/A vssd1 vssd1 vccd1 vccd1 _15526_/A sky130_fd_sc_hd__nor2_1
XFILLER_76_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19292_ _19100_/A _19290_/Y _19291_/Y vssd1 vssd1 vccd1 vccd1 _23524_/D sky130_fd_sc_hd__o21ba_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _12723_/X _12725_/X _21271_/B _12728_/Y _12941_/A vssd1 vssd1 vccd1 vccd1
+ _12738_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_187_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12460__A2 _12185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18243_ _18244_/A vssd1 vssd1 vccd1 vccd1 _18243_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15455_ _15455_/A _15485_/D vssd1 vssd1 vccd1 vccd1 _15457_/A sky130_fd_sc_hd__nand2_1
X_12667_ _12794_/B _12667_/B vssd1 vssd1 vccd1 vccd1 _13177_/B sky130_fd_sc_hd__nand2_2
XFILLER_187_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1099 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14406_ _14407_/A _15120_/B _14407_/C _14344_/B vssd1 vssd1 vccd1 vccd1 _14406_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__13122__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18174_ _18170_/Y _18171_/X _18173_/X vssd1 vssd1 vccd1 vccd1 _18176_/B sky130_fd_sc_hd__a21o_1
X_11618_ _11604_/X _18798_/B _11618_/C vssd1 vssd1 vccd1 vccd1 _12168_/A sky130_fd_sc_hd__and3b_2
XFILLER_168_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19676__A1 _19859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15386_ _15329_/A _15330_/A _15328_/Y vssd1 vssd1 vccd1 vccd1 _15386_/X sky130_fd_sc_hd__o21a_1
X_12598_ _13052_/A vssd1 vssd1 vccd1 vccd1 _12929_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17125_ _17125_/A _17125_/B vssd1 vssd1 vccd1 vccd1 _17298_/B sky130_fd_sc_hd__nand2_1
X_14337_ _13933_/A _14263_/Y _15075_/A _14183_/A _14260_/Y vssd1 vssd1 vccd1 vccd1
+ _14353_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_171_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17529__A _23526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17056_ _17964_/C _16142_/B _14730_/D vssd1 vssd1 vccd1 vccd1 _17444_/A sky130_fd_sc_hd__o21ai_2
XFILLER_143_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14268_ _14796_/A vssd1 vssd1 vccd1 vccd1 _15195_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16007_ _16004_/X _16005_/Y _16006_/Y vssd1 vssd1 vccd1 vccd1 _16008_/C sky130_fd_sc_hd__o21ai_1
X_13219_ _23319_/Q vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_994 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _14199_/A vssd1 vssd1 vccd1 vccd1 _14883_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13792__A _22064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_997 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _17958_/A vssd1 vssd1 vccd1 vccd1 _18211_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18939__B1 _19381_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16909_ _16911_/B _16908_/A _16913_/B vssd1 vssd1 vccd1 vccd1 _16909_/Y sky130_fd_sc_hd__a21oi_1
X_17889_ _16665_/X _17029_/X _17406_/B _17406_/A _17723_/B vssd1 vssd1 vccd1 vccd1
+ _17889_/Y sky130_fd_sc_hd__o2111ai_4
XANTENNA__17414__D _17414_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16414__A1 _16066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19628_ _19625_/A _19447_/B _19626_/X _19627_/X vssd1 vssd1 vccd1 vccd1 _19916_/C
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_26_628 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19559_ _19557_/X _19558_/X _19552_/B _19552_/C vssd1 vssd1 vccd1 vccd1 _19559_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__12436__C1 _19703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12987__B1 _20464_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17509__A4 _18376_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22570_ _22577_/A _22577_/B _22564_/X _22563_/Y vssd1 vssd1 vccd1 vccd1 _22573_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_90_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21171__B1 _20957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21521_ _21521_/A _21521_/B vssd1 vssd1 vccd1 vccd1 _21522_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17390__A2 _17323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21452_ _21510_/A _21510_/B _21510_/C vssd1 vssd1 vccd1 vccd1 _21463_/B sky130_fd_sc_hd__nand3_1
XFILLER_182_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20403_ _20403_/A _20403_/B vssd1 vssd1 vccd1 vccd1 _20405_/A sky130_fd_sc_hd__xnor2_1
XFILLER_119_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21383_ _21383_/A _21383_/B _21383_/C vssd1 vssd1 vccd1 vccd1 _21465_/A sky130_fd_sc_hd__nand3_2
XFILLER_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11962__A1 _11916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22064__B _22064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23122_ _23122_/A vssd1 vssd1 vccd1 vccd1 _23385_/D sky130_fd_sc_hd__clkbuf_1
X_20334_ _20335_/A _20363_/B vssd1 vssd1 vccd1 vccd1 _20336_/A sky130_fd_sc_hd__and2_1
XFILLER_135_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15153__B2 _15253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16062__B _16062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20265_ _20265_/A _20265_/B _20265_/C _20366_/C vssd1 vssd1 vccd1 vccd1 _20268_/A
+ sky130_fd_sc_hd__or4_1
X_23053_ _23110_/S vssd1 vssd1 vccd1 vccd1 _23062_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__13703__A2 _22388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22004_ _21999_/Y _22001_/Y _22003_/X _21920_/X vssd1 vssd1 vccd1 vccd1 _22076_/B
+ sky130_fd_sc_hd__o2bb2ai_2
X_20196_ _20207_/B _20196_/B _20196_/C _20196_/D vssd1 vssd1 vccd1 vccd1 _20196_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_163_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17605__C _20055_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22906_ _22906_/A vssd1 vssd1 vccd1 vccd1 _23289_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_1_1_0_bq_clk_i_A clkbuf_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22837_ _22792_/X _22797_/C _22836_/Y vssd1 vssd1 vccd1 vccd1 _22839_/A sky130_fd_sc_hd__o21a_1
XANTENNA__18158__A1 _17889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15422__A _15422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13570_ _13563_/A _22380_/C _13563_/C _22278_/B _13497_/A vssd1 vssd1 vccd1 vccd1
+ _13573_/A sky130_fd_sc_hd__a32o_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22768_ _22717_/A _22718_/X _22766_/Y vssd1 vssd1 vccd1 vccd1 _22789_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12442__A2 _12103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12521_ _18559_/A _18559_/B _12522_/C vssd1 vssd1 vccd1 vccd1 _12534_/A sky130_fd_sc_hd__a21oi_1
XFILLER_13_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21719_ _21723_/C _21719_/B vssd1 vssd1 vccd1 vccd1 _23556_/D sky130_fd_sc_hd__xor2_1
XFILLER_9_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22699_ _22700_/D _22566_/A _22566_/B _22700_/C _22790_/A vssd1 vssd1 vccd1 vccd1
+ _22701_/A sky130_fd_sc_hd__a32o_1
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15095_/X _15170_/Y _15179_/C _15239_/Y vssd1 vssd1 vccd1 vccd1 _15245_/B
+ sky130_fd_sc_hd__o211ai_2
X_12452_ _12447_/Y _12448_/X _12445_/C vssd1 vssd1 vccd1 vccd1 _18497_/B sky130_fd_sc_hd__o21ai_1
XFILLER_123_1050 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15171_ _15171_/A _15171_/B _15233_/C vssd1 vssd1 vccd1 vccd1 _15171_/Y sky130_fd_sc_hd__nand3_1
XFILLER_153_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12383_ _12368_/B _12366_/Y _12368_/A _12382_/X vssd1 vssd1 vccd1 vccd1 _12383_/Y
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__12781__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14122_ _14116_/X _14118_/X _14121_/Y vssd1 vssd1 vccd1 vccd1 _14133_/A sky130_fd_sc_hd__o21ai_1
XFILLER_180_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18930_ _18929_/X _18878_/Y _18886_/Y _18897_/D _18904_/Y vssd1 vssd1 vccd1 vccd1
+ _19075_/A sky130_fd_sc_hd__a32oi_4
X_14053_ _23496_/Q vssd1 vssd1 vccd1 vccd1 _14760_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_122_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ _12725_/A _12854_/Y _13002_/Y _13003_/Y vssd1 vssd1 vccd1 vccd1 _13004_/X
+ sky130_fd_sc_hd__a22o_1
X_18861_ _18862_/A _18862_/B _18862_/C vssd1 vssd1 vccd1 vccd1 _18863_/A sky130_fd_sc_hd__a21oi_1
XFILLER_133_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17812_ _17924_/A _17807_/Y _17662_/A _17669_/X vssd1 vssd1 vccd1 vccd1 _17814_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__17841__B1 _17414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18792_ _11736_/A _12409_/A _12413_/A _18971_/A vssd1 vssd1 vccd1 vccd1 _18792_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17743_ _17741_/X _17742_/X _18778_/A _17243_/D vssd1 vssd1 vccd1 vccd1 _17750_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14955_ _14957_/B _14957_/A vssd1 vssd1 vccd1 vccd1 _14956_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22193__A2 _22192_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13906_ _14023_/C vssd1 vssd1 vccd1 vccd1 _14191_/B sky130_fd_sc_hd__clkbuf_2
X_17674_ _17498_/B _17498_/C _17498_/A _17502_/C _17502_/A vssd1 vssd1 vccd1 vccd1
+ _17674_/X sky130_fd_sc_hd__a32o_1
X_14886_ _14886_/A _14886_/B _14886_/C vssd1 vssd1 vccd1 vccd1 _14887_/B sky130_fd_sc_hd__nand3_1
XFILLER_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19413_ _19413_/A _19413_/B _19413_/C vssd1 vssd1 vccd1 vccd1 _19437_/A sky130_fd_sc_hd__nand3_1
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16625_ _16812_/A vssd1 vssd1 vccd1 vccd1 _16625_/X sky130_fd_sc_hd__buf_2
X_13837_ _13646_/B _13646_/C _13646_/A _13671_/B _13671_/C vssd1 vssd1 vccd1 vccd1
+ _13839_/B sky130_fd_sc_hd__a32oi_4
XFILLER_51_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12956__A _21054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19344_ _19218_/X _17643_/A _19194_/X _19201_/A vssd1 vssd1 vccd1 vccd1 _19345_/C
+ sky130_fd_sc_hd__o31a_1
X_16556_ _16545_/Y _16555_/Y _16500_/Y _16503_/Y vssd1 vssd1 vccd1 vccd1 _16556_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13768_ _13257_/A _13765_/X _13769_/A _13767_/Y _13663_/C vssd1 vssd1 vccd1 vccd1
+ _13768_/Y sky130_fd_sc_hd__o2111ai_4
XANTENNA__11641__B1 _11915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15507_ _15419_/C _15419_/D _15446_/D _15536_/A vssd1 vssd1 vccd1 vccd1 _15513_/C
+ sky130_fd_sc_hd__a31o_1
X_12719_ _12923_/C _13138_/D vssd1 vssd1 vccd1 vccd1 _12776_/B sky130_fd_sc_hd__nand2_1
X_19275_ _19275_/A _19275_/B _19275_/C vssd1 vssd1 vccd1 vccd1 _19275_/Y sky130_fd_sc_hd__nand3_4
X_16487_ _16416_/X _16420_/Y _16426_/Y _16427_/X vssd1 vssd1 vccd1 vccd1 _16488_/A
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__21988__B _21988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13699_ _13698_/B _13587_/B _13578_/Y _13590_/Y vssd1 vssd1 vccd1 vccd1 _13730_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_176_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18226_ _18226_/A _18226_/B vssd1 vssd1 vccd1 vccd1 _18268_/A sky130_fd_sc_hd__xnor2_1
XFILLER_15_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15438_ _15438_/A _15438_/B vssd1 vssd1 vccd1 vccd1 _15439_/B sky130_fd_sc_hd__xor2_4
XFILLER_175_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_639 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18157_ _18163_/A _18157_/B _18157_/C _18157_/D vssd1 vssd1 vccd1 vccd1 _18157_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_157_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17259__A _17259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _15369_/A _15369_/B vssd1 vssd1 vccd1 vccd1 _15370_/A sky130_fd_sc_hd__and2_1
XFILLER_8_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17108_ _19662_/C _17108_/B _19485_/A _17259_/A vssd1 vssd1 vccd1 vccd1 _17112_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__16868__D1 _17226_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18088_ _18163_/A _18088_/B _18088_/C _18161_/C vssd1 vssd1 vccd1 vccd1 _18090_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_172_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16332__B1 _16330_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17039_ _17039_/A _17039_/B vssd1 vssd1 vccd1 vccd1 _17039_/Y sky130_fd_sc_hd__nand2_2
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19806__D1 _20055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22956__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20050_ _20209_/A _17600_/A _20049_/Y vssd1 vssd1 vccd1 vccd1 _20050_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__19193__B _19700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18624__A2 _18931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater110 _23298_/CLK vssd1 vssd1 vccd1 vccd1 _23295_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater121 _23397_/CLK vssd1 vssd1 vccd1 vccd1 _23391_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater132 _23339_/CLK vssd1 vssd1 vccd1 vccd1 _23345_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater143 _23437_/CLK vssd1 vssd1 vccd1 vccd1 _23435_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater154 _23430_/CLK vssd1 vssd1 vccd1 vccd1 _23431_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17045__D1 _16499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17722__A _17722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ _21295_/B vssd1 vssd1 vccd1 vccd1 _21497_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_723 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ _20883_/A vssd1 vssd1 vccd1 vccd1 _23542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22622_ _22623_/B _22623_/C _22623_/A vssd1 vssd1 vccd1 vccd1 _22818_/A sky130_fd_sc_hd__a21o_1
XFILLER_35_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19649__A _19649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22553_ _22553_/A _22554_/A _22553_/C _22553_/D vssd1 vssd1 vccd1 vccd1 _22649_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_167_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21504_ _21504_/A _21504_/B vssd1 vssd1 vccd1 vccd1 _21554_/B sky130_fd_sc_hd__nor2_1
XANTENNA__15374__A1 _15422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22484_ _22484_/A vssd1 vssd1 vccd1 vccd1 _22484_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21435_ _21502_/A _21440_/C _21435_/C _21497_/A vssd1 vssd1 vccd1 vccd1 _21435_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_182_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21366_ _21502_/D _21386_/A _21293_/Y _21300_/X vssd1 vssd1 vccd1 vccd1 _21377_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23105_ _23105_/A vssd1 vssd1 vccd1 vccd1 _23378_/D sky130_fd_sc_hd__clkbuf_1
X_20317_ _20317_/A _20317_/B _20317_/C vssd1 vssd1 vccd1 vccd1 _20317_/X sky130_fd_sc_hd__and3_1
XFILLER_163_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16801__A _16815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21297_ _21293_/Y _21295_/Y _21296_/X vssd1 vssd1 vccd1 vccd1 _21298_/C sky130_fd_sc_hd__a21bo_1
XFILLER_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22947__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18076__B1 _18001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23036_ _23348_/Q input30/X _23038_/S vssd1 vssd1 vccd1 vccd1 _23037_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20248_ _20189_/B _20189_/C _20189_/A vssd1 vssd1 vccd1 vccd1 _20248_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__19812__A1 _19190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1043 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20363__A_N _20335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19534__D _19534_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11945__A _23591_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20179_ _20172_/A _20172_/B _20170_/Y vssd1 vssd1 vccd1 vccd1 _20179_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_78 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21907__C1 _22043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17632__A _17712_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14740_ _14734_/X _11798_/A _14738_/X vssd1 vssd1 vccd1 vccd1 _23263_/D sky130_fd_sc_hd__a21o_1
XFILLER_85_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _11948_/X _11951_/X _12066_/A vssd1 vssd1 vccd1 vccd1 _11952_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16929__A2 _16662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _23400_/Q _14640_/X _14647_/X _23432_/Q _14670_/X vssd1 vssd1 vccd1 vccd1
+ _14671_/X sky130_fd_sc_hd__a221o_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11883_ _11883_/A vssd1 vssd1 vccd1 vccd1 _11883_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16410_ _18503_/B vssd1 vssd1 vccd1 vccd1 _17406_/B sky130_fd_sc_hd__buf_4
X_13622_ _21752_/A vssd1 vssd1 vccd1 vccd1 _22292_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17390_ _16529_/C _17323_/X _17324_/X _17549_/A _17392_/A vssd1 vssd1 vccd1 vccd1
+ _17810_/C sky130_fd_sc_hd__a32o_1
XANTENNA__13612__A1 _13552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16341_ _16340_/C _16340_/A _16340_/B vssd1 vssd1 vccd1 vccd1 _16341_/X sky130_fd_sc_hd__a21o_1
XFILLER_198_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13553_ _13553_/A vssd1 vssd1 vccd1 vccd1 _13553_/X sky130_fd_sc_hd__buf_2
XFILLER_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19060_ _19060_/A _19060_/B vssd1 vssd1 vccd1 vccd1 _19063_/B sky130_fd_sc_hd__nand2_1
X_12504_ _23593_/Q vssd1 vssd1 vccd1 vccd1 _23260_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_73_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15365__A1 _14097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16272_ _16275_/A _16281_/C _16281_/D vssd1 vssd1 vccd1 vccd1 _16272_/Y sky130_fd_sc_hd__nand3_1
X_13484_ _13483_/B _13483_/C _13264_/C vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__a21bo_1
XFILLER_173_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12179__A1 _12167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18011_ _18016_/C _17391_/B _17391_/C _20164_/C _17899_/B vssd1 vssd1 vccd1 vccd1
+ _18013_/C sky130_fd_sc_hd__a32o_1
X_15223_ _15298_/B vssd1 vssd1 vccd1 vccd1 _15455_/A sky130_fd_sc_hd__clkbuf_2
X_12435_ _12435_/A _12435_/B vssd1 vssd1 vccd1 vccd1 _19703_/A sky130_fd_sc_hd__nand2_4
XFILLER_172_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19500__B1 _20209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20217__B _20217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15154_ _15267_/B _15267_/C _15488_/A _14020_/Y vssd1 vssd1 vccd1 vccd1 _15154_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_12366_ _12366_/A vssd1 vssd1 vccd1 vccd1 _12366_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14105_ _14105_/A vssd1 vssd1 vccd1 vccd1 _15001_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19962_ _19860_/X _19943_/Y _19960_/Y _19944_/Y vssd1 vssd1 vccd1 vccd1 _19963_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15085_ _15488_/A _15085_/B _15085_/C vssd1 vssd1 vccd1 vccd1 _15085_/X sky130_fd_sc_hd__or3_1
XFILLER_141_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12297_ _12297_/A _12297_/B _12297_/C _12297_/D vssd1 vssd1 vccd1 vccd1 _12298_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22938__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18913_ _18902_/A _18903_/A _18914_/C vssd1 vssd1 vccd1 vccd1 _18913_/X sky130_fd_sc_hd__a21o_1
X_14036_ _14075_/A _14261_/A _14790_/C vssd1 vssd1 vccd1 vccd1 _14039_/A sky130_fd_sc_hd__nand3_2
XANTENNA__23060__A0 _14070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output75_A _14714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18606__A2 _18604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19893_ _19893_/A _19893_/B _19897_/A _19897_/B vssd1 vssd1 vccd1 vccd1 _19894_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_171_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11855__A _16365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18844_ _18844_/A _18844_/B _18844_/C _18844_/D vssd1 vssd1 vccd1 vccd1 _18845_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18775_ _18969_/A _18966_/A _18966_/B vssd1 vssd1 vccd1 vccd1 _18775_/Y sky130_fd_sc_hd__a21oi_1
X_15987_ _15858_/B _15969_/X _15995_/A _16181_/A _15993_/A vssd1 vssd1 vccd1 vccd1
+ _15999_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_83_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17726_ _19674_/B vssd1 vssd1 vccd1 vccd1 _19951_/D sky130_fd_sc_hd__buf_2
XANTENNA__19031__A2 _19218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14938_ _14938_/A _14938_/B vssd1 vssd1 vccd1 vccd1 _14939_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17657_ _17657_/A _17657_/B _17657_/C vssd1 vssd1 vccd1 vccd1 _17658_/C sky130_fd_sc_hd__nand3_1
XFILLER_24_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14869_ _14970_/B vssd1 vssd1 vccd1 vccd1 _14883_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23115__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11590__A _23598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16608_ _16608_/A vssd1 vssd1 vccd1 vccd1 _16647_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_51_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_992 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17588_ _20142_/A vssd1 vssd1 vccd1 vccd1 _18077_/A sky130_fd_sc_hd__buf_2
XFILLER_32_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19327_ _19805_/A _19327_/B _19804_/A vssd1 vssd1 vccd1 vccd1 _19478_/A sky130_fd_sc_hd__nand3_2
XFILLER_91_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16539_ _16539_/A _16539_/B _16539_/C vssd1 vssd1 vccd1 vccd1 _16539_/X sky130_fd_sc_hd__and3_1
XFILLER_32_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18373__A _18373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19258_ _19256_/X _19257_/Y _19245_/X _19254_/Y vssd1 vssd1 vccd1 vccd1 _19259_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_31_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18209_ _18209_/A vssd1 vssd1 vccd1 vccd1 _18298_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_164_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19189_ _19189_/A vssd1 vssd1 vccd1 vccd1 _19189_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21220_ _21218_/X _21219_/Y _21215_/A vssd1 vssd1 vccd1 vccd1 _21221_/C sky130_fd_sc_hd__o21bai_2
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21151_ _20884_/X _20885_/X _20996_/X _20998_/Y vssd1 vssd1 vccd1 vccd1 _21151_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_172_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22929__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20102_ _20102_/A _20102_/B vssd1 vssd1 vccd1 vccd1 _20106_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23051__A0 _13911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13964__B _14331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21082_ _21082_/A _21082_/B _21082_/C vssd1 vssd1 vccd1 vccd1 _21083_/B sky130_fd_sc_hd__nand3_4
XFILLER_99_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20033_ _20031_/X _20207_/A _20029_/Y vssd1 vssd1 vccd1 vccd1 _20033_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17266__D1 _20049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_712 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13980__A _23502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20797__B _23297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21984_ _21984_/A _21984_/B _21984_/C _21984_/D vssd1 vssd1 vccd1 vccd1 _21984_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_840 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ _21169_/A _21277_/A _21050_/C _21177_/B vssd1 vssd1 vccd1 vccd1 _20940_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_148_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16068__A _19659_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23106__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17584__A2 _17565_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _20862_/A _20862_/B _20863_/A vssd1 vssd1 vccd1 vccd1 _20872_/A sky130_fd_sc_hd__o21ai_1
XFILLER_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22605_ _22605_/A _22633_/A vssd1 vssd1 vccd1 vccd1 _22610_/A sky130_fd_sc_hd__nand2_1
X_23585_ _23588_/CLK _23585_/D vssd1 vssd1 vccd1 vccd1 _23585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18533__A1 _11851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20797_ _23296_/Q _23297_/Q _23298_/Q vssd1 vssd1 vccd1 vccd1 _20897_/D sky130_fd_sc_hd__nor3_1
XFILLER_195_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22536_ _22536_/A _22536_/B vssd1 vssd1 vccd1 vccd1 _23566_/D sky130_fd_sc_hd__xor2_4
XFILLER_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22467_ _13495_/X _22757_/B _22567_/A vssd1 vssd1 vccd1 vccd1 _22468_/A sky130_fd_sc_hd__o21ai_1
XFILLER_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12220_ _12531_/A _12531_/B _12531_/C vssd1 vssd1 vccd1 vccd1 _12220_/Y sky130_fd_sc_hd__nand3_2
XFILLER_185_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21418_ _21418_/A _21418_/B _21418_/C vssd1 vssd1 vccd1 vccd1 _21418_/Y sky130_fd_sc_hd__nand3_1
XFILLER_182_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22398_ _22400_/A _22400_/B _22412_/A _22400_/D vssd1 vssd1 vccd1 vccd1 _22398_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_120_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12581__A1 _20799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_992 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17627__A _17627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ _12146_/X _12147_/X _12149_/X _19010_/A _19700_/B vssd1 vssd1 vccd1 vccd1
+ _12151_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_155_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21349_ _23566_/Q _21349_/B vssd1 vssd1 vccd1 vccd1 _21352_/A sky130_fd_sc_hd__xor2_1
XFILLER_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16531__A _16531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12082_ _23256_/B _11947_/A _23258_/B _16807_/A vssd1 vssd1 vccd1 vccd1 _18600_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_123_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13874__B _21971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23019_ _23340_/Q input21/X _23023_/S vssd1 vssd1 vccd1 vccd1 _23020_/A sky130_fd_sc_hd__mux2_1
X_15910_ _16209_/A vssd1 vssd1 vccd1 vccd1 _15910_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_314 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16890_ _16893_/A _16890_/B _16893_/C vssd1 vssd1 vccd1 vccd1 _16890_/X sky130_fd_sc_hd__and3_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _16126_/A _15841_/B _16612_/A vssd1 vssd1 vccd1 vccd1 _15975_/A sky130_fd_sc_hd__nand3_4
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15822__A2 _11883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _18560_/A vssd1 vssd1 vccd1 vccd1 _18728_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15772_ _15612_/A _15612_/B _12241_/A vssd1 vssd1 vccd1 vccd1 _15772_/X sky130_fd_sc_hd__a21o_2
X_12984_ _12984_/A _12984_/B vssd1 vssd1 vccd1 vccd1 _13106_/A sky130_fd_sc_hd__nor2_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22699__A3 _22566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23514__D input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17511_ _17504_/Y _17677_/C _17510_/Y vssd1 vssd1 vccd1 vccd1 _17700_/A sky130_fd_sc_hd__o21ai_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14723_ _23594_/Q vssd1 vssd1 vccd1 vccd1 _16800_/D sky130_fd_sc_hd__clkbuf_2
X_11935_ _11935_/A vssd1 vssd1 vccd1 vccd1 _11935_/X sky130_fd_sc_hd__clkbuf_4
X_18491_ _19499_/A vssd1 vssd1 vccd1 vccd1 _19670_/B sky130_fd_sc_hd__clkbuf_4
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17442_ _17433_/X _17437_/X _17580_/A vssd1 vssd1 vccd1 vccd1 _17446_/A sky130_fd_sc_hd__o21ai_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _21853_/A vssd1 vssd1 vccd1 vccd1 _21852_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _11864_/X _11865_/X _19363_/A _19363_/B vssd1 vssd1 vccd1 vccd1 _11866_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13358_/X _13602_/A _13603_/X _13394_/B vssd1 vssd1 vccd1 vccd1 _21752_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_14_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17373_ _16988_/Y _16989_/Y _16777_/Y _16998_/C vssd1 vssd1 vccd1 vccd1 _17374_/B
+ sky130_fd_sc_hd__o211a_1
X_14585_ input50/X _14549_/X _14547_/X _12675_/X vssd1 vssd1 vccd1 vccd1 _14585_/X
+ sky130_fd_sc_hd__a22o_1
X_11797_ _16049_/D _18859_/C _11788_/Y _11803_/A vssd1 vssd1 vccd1 vccd1 _11805_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16706__A _16706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19721__B1 _12324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19112_ _18941_/B _17581_/A _18778_/B _19113_/C _19262_/A vssd1 vssd1 vccd1 vccd1
+ _19116_/A sky130_fd_sc_hd__a32o_2
X_16324_ _16322_/X _16323_/Y _16313_/B _16313_/C vssd1 vssd1 vccd1 vccd1 _16324_/Y
+ sky130_fd_sc_hd__a22oi_4
X_13536_ _13537_/A _13536_/B _13536_/C vssd1 vssd1 vccd1 vccd1 _13755_/C sky130_fd_sc_hd__nand3_1
XFILLER_174_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15889__A2 _12223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19043_ _19043_/A vssd1 vssd1 vccd1 vccd1 _19047_/A sky130_fd_sc_hd__clkbuf_2
X_16255_ _16240_/Y _16251_/X _16242_/A _16242_/B vssd1 vssd1 vccd1 vccd1 _16255_/X
+ sky130_fd_sc_hd__o211a_1
X_13467_ _13660_/A _21925_/B _13660_/C vssd1 vssd1 vccd1 vccd1 _13467_/X sky130_fd_sc_hd__and3_1
XANTENNA__21050__C _21050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15206_ _15221_/A _15277_/B _15222_/A vssd1 vssd1 vccd1 vccd1 _15282_/A sky130_fd_sc_hd__a21o_1
XFILLER_127_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12418_ _19180_/D _19123_/C _12455_/C _12455_/D vssd1 vssd1 vccd1 vccd1 _12423_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12021__B1 _18755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11569__B _23583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16186_ _23424_/Q _23425_/Q vssd1 vssd1 vccd1 vccd1 _16667_/C sky130_fd_sc_hd__nor2_2
X_13398_ _23472_/Q vssd1 vssd1 vccd1 vccd1 _13600_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_142_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15137_ _15136_/B _15136_/C _15074_/Y vssd1 vssd1 vccd1 vccd1 _15140_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__21292__C1 _21431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12349_ _12366_/A _12348_/B _12348_/C vssd1 vssd1 vccd1 vccd1 _12372_/B sky130_fd_sc_hd__a21o_1
XFILLER_141_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19945_ _20142_/C vssd1 vssd1 vccd1 vccd1 _20371_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15068_ _14957_/B _14957_/A _15063_/A _15067_/X _15065_/Y vssd1 vssd1 vccd1 vccd1
+ _15068_/X sky130_fd_sc_hd__o221a_1
XFILLER_101_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11585__A _16593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ _14120_/B vssd1 vssd1 vccd1 vccd1 _14901_/A sky130_fd_sc_hd__buf_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19876_ _19939_/A _19876_/B _19876_/C vssd1 vssd1 vccd1 vccd1 _19876_/X sky130_fd_sc_hd__and3_1
XFILLER_110_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17263__A1 _17586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17263__B2 _17454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18827_ _18844_/A _18844_/B vssd1 vssd1 vccd1 vccd1 _18872_/A sky130_fd_sc_hd__nand2_2
XFILLER_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18758_ _11766_/A _18604_/A _18765_/A vssd1 vssd1 vccd1 vccd1 _18758_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__19004__A2 _19190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17709_ _17667_/A _17666_/B _17666_/A vssd1 vssd1 vccd1 vccd1 _17709_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18689_ _18673_/X _17643_/X _18674_/X _18675_/X _18688_/Y vssd1 vssd1 vccd1 vccd1
+ _18689_/X sky130_fd_sc_hd__o311a_1
XFILLER_64_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20720_ _20718_/Y _20719_/X _20618_/Y _20700_/X vssd1 vssd1 vccd1 vccd1 _20854_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19199__A _19662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20651_ _12675_/X _12704_/X _12711_/Y _12705_/X _23452_/Q vssd1 vssd1 vccd1 vccd1
+ _20652_/B sky130_fd_sc_hd__o311a_1
XFILLER_149_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23370_ _23372_/CLK _23370_/D vssd1 vssd1 vccd1 vccd1 _23370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20582_ _21493_/C vssd1 vssd1 vccd1 vccd1 _21387_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22321_ _22314_/A _22314_/B _22291_/Y _22313_/X vssd1 vssd1 vccd1 vccd1 _22324_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_178_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22252_ _22252_/A _23274_/Q _22252_/C vssd1 vssd1 vccd1 vccd1 _22451_/C sky130_fd_sc_hd__nand3_1
XFILLER_145_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21203_ _12785_/X _21061_/X _12862_/X _21545_/A vssd1 vssd1 vccd1 vccd1 _21203_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16829__B2 _15856_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22183_ _22388_/C _22160_/B _22182_/X vssd1 vssd1 vccd1 vccd1 _22183_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_172_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21134_ _21134_/A _21134_/B _21134_/C vssd1 vssd1 vccd1 vccd1 _21153_/B sky130_fd_sc_hd__nand3_1
XFILLER_132_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12315__A1 _12353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21065_ _21065_/A vssd1 vssd1 vccd1 vccd1 _21196_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16057__A2 _16055_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20016_ _20108_/B _20111_/A _20108_/A vssd1 vssd1 vccd1 vccd1 _20016_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_171_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23184__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19381__B _19381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20320__B _20320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21967_ _13870_/A _13870_/B _21858_/D vssd1 vssd1 vccd1 vccd1 _21981_/C sky130_fd_sc_hd__o21ai_4
XFILLER_73_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16214__C1 _17753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11720_/A vssd1 vssd1 vccd1 vccd1 _11798_/A sky130_fd_sc_hd__clkbuf_2
X_20918_ _20495_/A _14615_/X _21047_/B _12571_/X vssd1 vssd1 vccd1 vccd1 _20918_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_70_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21898_ _22029_/A _21898_/B _21898_/C _22020_/B vssd1 vssd1 vccd1 vccd1 _21905_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21432__A _21432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11649_/X _11721_/A _23587_/Q vssd1 vssd1 vccd1 vccd1 _15704_/B sky130_fd_sc_hd__a21o_2
XFILLER_187_539 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20849_ _20849_/A _20849_/B vssd1 vssd1 vccd1 vccd1 _20849_/Y sky130_fd_sc_hd__nand2_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16526__A _16526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14370_ _14310_/Y _14311_/X _14369_/X vssd1 vssd1 vccd1 vccd1 _14847_/A sky130_fd_sc_hd__a21o_1
XFILLER_167_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23568_ _23575_/CLK _23568_/D vssd1 vssd1 vccd1 vccd1 _23568_/Q sky130_fd_sc_hd__dfxtp_1
X_11582_ _11582_/A _23590_/Q _11739_/A vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__nand3_1
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12773__B _12845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13321_ _13394_/B vssd1 vssd1 vccd1 vccd1 _13483_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_11_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22519_ _22609_/A _22607_/A _22607_/B vssd1 vssd1 vccd1 vccd1 _22524_/C sky130_fd_sc_hd__a21o_1
XFILLER_13_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23499_ _23499_/CLK _23499_/D vssd1 vssd1 vccd1 vccd1 _23499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ _15920_/A _15678_/Y _12018_/X _12020_/X _15682_/D vssd1 vssd1 vccd1 vccd1
+ _16310_/B sky130_fd_sc_hd__o221a_1
XFILLER_183_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22066__A1 _13642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13252_ _23320_/Q _23319_/Q _23318_/Q vssd1 vssd1 vccd1 vccd1 _13344_/A sky130_fd_sc_hd__nor3_2
XFILLER_143_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15740__A1 _15864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12203_ _12203_/A _12203_/B _12203_/C vssd1 vssd1 vccd1 vccd1 _12203_/Y sky130_fd_sc_hd__nand3_4
XFILLER_109_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13183_ _13181_/A _20563_/A _20563_/B _13181_/C vssd1 vssd1 vccd1 vccd1 _13186_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_135_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23509__D input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ _11849_/C _11849_/A _19308_/B _12133_/Y _19363_/B vssd1 vssd1 vccd1 vccd1
+ _12134_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_123_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17991_ _12088_/X _18002_/A _18157_/D _18157_/B vssd1 vssd1 vccd1 vccd1 _17991_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13503__B1 _22392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19730_ _19730_/A _19730_/B vssd1 vssd1 vccd1 vccd1 _19731_/B sky130_fd_sc_hd__nor2_1
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16942_ _16948_/A _16948_/B _16948_/C vssd1 vssd1 vccd1 vccd1 _16942_/X sky130_fd_sc_hd__and3_1
X_12065_ _11719_/X _12061_/Y _12391_/C vssd1 vssd1 vccd1 vccd1 _12542_/A sky130_fd_sc_hd__o21ai_2
XFILLER_111_539 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16048__A2 _11792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20919__A3 _21050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19661_ _18476_/X _18484_/X _19846_/A _19659_/C vssd1 vssd1 vccd1 vccd1 _19662_/A
+ sky130_fd_sc_hd__o211a_1
X_16873_ _16893_/A _16890_/B _16873_/C vssd1 vssd1 vccd1 vccd1 _16873_/X sky130_fd_sc_hd__and3_1
XFILLER_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12013__B _18859_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18993__A1 _16032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18612_ _12167_/X _12168_/X _18080_/A _18605_/Y vssd1 vssd1 vccd1 vccd1 _18615_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__18993__B2 _18440_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15605__A _15605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15824_ _16020_/A _16020_/B _16020_/C vssd1 vssd1 vccd1 vccd1 _16062_/B sky130_fd_sc_hd__nand3_4
X_19592_ _19592_/A _19592_/B _19592_/C vssd1 vssd1 vccd1 vccd1 _19609_/B sky130_fd_sc_hd__nand3_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12609__A2 _20495_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12948__B _21054_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _18721_/A _18541_/A _12478_/B _18524_/B vssd1 vssd1 vccd1 vccd1 _18553_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15755_ _15735_/C _15662_/B _23416_/Q _15624_/A _15665_/B vssd1 vssd1 vccd1 vccd1
+ _15757_/A sky130_fd_sc_hd__o311ai_4
X_12967_ _21079_/A vssd1 vssd1 vccd1 vccd1 _21295_/B sky130_fd_sc_hd__buf_2
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _11918_/A _11918_/B _16802_/B _16141_/A vssd1 vssd1 vccd1 vccd1 _11959_/A
+ sky130_fd_sc_hd__nand4_2
X_14706_ _23345_/Q _14689_/X _14694_/X _23313_/Q _14699_/X vssd1 vssd1 vccd1 vccd1
+ _14706_/X sky130_fd_sc_hd__a221o_1
XFILLER_166_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18474_ _18474_/A vssd1 vssd1 vccd1 vccd1 _18474_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ _12899_/B _12899_/C _12899_/A vssd1 vssd1 vccd1 vccd1 _13044_/A sky130_fd_sc_hd__a21o_1
X_15686_ _15686_/A _15686_/B _16187_/C vssd1 vssd1 vccd1 vccd1 _15686_/X sky130_fd_sc_hd__and3_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _17425_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17426_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11849_ _11849_/A _18657_/C _11849_/C vssd1 vssd1 vccd1 vccd1 _18474_/A sky130_fd_sc_hd__nand3_2
X_14637_ _23331_/Q _14636_/X _14547_/A _23299_/Q _14587_/X vssd1 vssd1 vccd1 vccd1
+ _14637_/X sky130_fd_sc_hd__a221o_1
XANTENNA__15978__C _16314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15340__A _15402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17356_ _17361_/B _17514_/A _17359_/B vssd1 vssd1 vccd1 vccd1 _17357_/B sky130_fd_sc_hd__nand3_1
X_14568_ input47/X _14518_/X _14547_/X _12601_/B vssd1 vssd1 vccd1 vccd1 _14568_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12793__A1 _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16307_ _16389_/A _16322_/B _16402_/B _16323_/A vssd1 vssd1 vccd1 vccd1 _16313_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_13519_ _13519_/A _13519_/B _13519_/C vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__nand3_1
XFILLER_173_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17287_ _17284_/X _17286_/X _17276_/A vssd1 vssd1 vccd1 vccd1 _17287_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_147_959 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14499_ _14846_/A _14846_/B _14847_/A _14847_/B vssd1 vssd1 vccd1 vccd1 _14853_/A
+ sky130_fd_sc_hd__nand4_1
X_19026_ _19026_/A _19026_/B _19026_/C vssd1 vssd1 vccd1 vccd1 _19138_/A sky130_fd_sc_hd__nand3_2
X_16238_ _16236_/X _15926_/X _15929_/Y _16251_/B vssd1 vssd1 vccd1 vccd1 _16253_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_133_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16171__A _17062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16169_ _16170_/A _16650_/A _16169_/C vssd1 vssd1 vccd1 vccd1 _16169_/Y sky130_fd_sc_hd__nand3_2
XFILLER_173_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21280__A2 _21453_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_815 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19928_ _19928_/A _19928_/B _19928_/C _19928_/D vssd1 vssd1 vccd1 vccd1 _19929_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19482__A _19482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19859_ _19859_/A vssd1 vssd1 vccd1 vccd1 _20210_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_56_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22870_ _22529_/A _22849_/X _22868_/Y _22848_/Y vssd1 vssd1 vccd1 vccd1 _22878_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_23_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21821_ _21810_/Y _21813_/X _21824_/C vssd1 vssd1 vccd1 vccd1 _21844_/A sky130_fd_sc_hd__o21bai_2
XFILLER_97_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15445__A1_N _15446_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16049__C _17414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21752_ _21752_/A _21752_/B _21909_/C vssd1 vssd1 vccd1 vccd1 _21753_/B sky130_fd_sc_hd__and3_1
XFILLER_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20703_ _20553_/A _20701_/X _20702_/Y vssd1 vssd1 vccd1 vccd1 _20703_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16211__A2 _15655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21683_ _21650_/A _21650_/B _21631_/Y vssd1 vssd1 vccd1 vccd1 _21704_/A sky130_fd_sc_hd__a21oi_1
XFILLER_24_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14792__C _23502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_bq_clk_i_A clkbuf_4_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23422_ _23427_/CLK _23422_/D vssd1 vssd1 vccd1 vccd1 _23422_/Q sky130_fd_sc_hd__dfxtp_1
X_20634_ _20634_/A _20634_/B vssd1 vssd1 vccd1 vccd1 _20635_/C sky130_fd_sc_hd__nand2_1
XFILLER_149_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23353_ _23365_/CLK _23353_/D vssd1 vssd1 vccd1 vccd1 _23353_/Q sky130_fd_sc_hd__dfxtp_1
X_20565_ _20565_/A _20704_/B _20773_/D _20565_/D vssd1 vssd1 vccd1 vccd1 _20566_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_166_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16514__A3 _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22304_ _22300_/Y _22301_/Y _22303_/Y vssd1 vssd1 vccd1 vccd1 _22403_/A sky130_fd_sc_hd__a21o_1
XFILLER_192_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23284_ _23492_/CLK _23284_/D vssd1 vssd1 vccd1 vccd1 _23284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20496_ _20782_/A vssd1 vssd1 vccd1 vccd1 _20496_/X sky130_fd_sc_hd__buf_2
XFILLER_4_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22235_ _22090_/C _22086_/A _22228_/Y _22234_/Y vssd1 vssd1 vccd1 vccd1 _22242_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_106_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22166_ _22166_/A _22166_/B _22166_/C vssd1 vssd1 vccd1 vccd1 _22166_/Y sky130_fd_sc_hd__nand3_4
XFILLER_133_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21117_ _21159_/A _21228_/A _21159_/B vssd1 vssd1 vccd1 vccd1 _21119_/B sky130_fd_sc_hd__nand3_1
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22097_ _21874_/A _21874_/B _22096_/X vssd1 vssd1 vccd1 vccd1 _22099_/C sky130_fd_sc_hd__o21ai_4
XANTENNA__17227__A1 _16604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21048_ _21048_/A _21048_/B vssd1 vssd1 vccd1 vccd1 _21181_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14779__C_N _14246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13870_ _13870_/A _13870_/B vssd1 vssd1 vccd1 vccd1 _13870_/Y sky130_fd_sc_hd__nor2_2
XFILLER_28_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ _12754_/A _13151_/C _12770_/C _12820_/X vssd1 vssd1 vccd1 vccd1 _12837_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22999_ _23331_/Q input11/X _23001_/S vssd1 vssd1 vccd1 vccd1 _23000_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15540_ _15540_/A _15540_/B vssd1 vssd1 vccd1 vccd1 _15540_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12752_ _20962_/A _20681_/C _20962_/C vssd1 vssd1 vccd1 vccd1 _12754_/A sky130_fd_sc_hd__nand3_2
XANTENNA__12472__B1 _12151_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_854 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11703_ _11686_/B _11676_/X _11672_/Y vssd1 vssd1 vccd1 vccd1 _11704_/B sky130_fd_sc_hd__o21ai_1
X_15471_ _15471_/A _15501_/A _15471_/C vssd1 vssd1 vccd1 vccd1 _15501_/B sky130_fd_sc_hd__nand3_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _23293_/Q _12683_/B vssd1 vssd1 vccd1 vccd1 _12683_/Y sky130_fd_sc_hd__nand2_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14213__A1 _14207_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17025_/A _16982_/X _16994_/D vssd1 vssd1 vccd1 vccd1 _17210_/X sky130_fd_sc_hd__o21a_1
X_14422_ _14422_/A _14422_/B _14422_/C vssd1 vssd1 vccd1 vccd1 _14495_/D sky130_fd_sc_hd__nand3_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12224__B1 _12090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ _11634_/A _11634_/B vssd1 vssd1 vccd1 vccd1 _11634_/Y sky130_fd_sc_hd__nand2_1
X_18190_ _18245_/A _18126_/A _18209_/A vssd1 vssd1 vccd1 vccd1 _18191_/B sky130_fd_sc_hd__a21o_1
XANTENNA__15961__A1 _11916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17141_ _16908_/X _17307_/A _17898_/D _17140_/Y _19653_/A vssd1 vssd1 vccd1 vccd1
+ _17145_/B sky130_fd_sc_hd__o2111ai_1
X_14353_ _14353_/A _14353_/B _14353_/C vssd1 vssd1 vccd1 vccd1 _14353_/X sky130_fd_sc_hd__and3_1
XFILLER_7_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13304_ _23323_/Q vssd1 vssd1 vccd1 vccd1 _13304_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17072_ _17089_/A _17089_/B _17067_/X _17071_/X vssd1 vssd1 vccd1 vccd1 _17221_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14284_ _14284_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14285_/A sky130_fd_sc_hd__nand2_1
XFILLER_143_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13235_ _13659_/B vssd1 vssd1 vccd1 vccd1 _13563_/A sky130_fd_sc_hd__clkbuf_2
X_16023_ _16021_/Y _16022_/Y _15895_/C vssd1 vssd1 vccd1 vccd1 _16347_/C sky130_fd_sc_hd__o21ai_2
XFILLER_108_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13166_ _13166_/A _13177_/A vssd1 vssd1 vccd1 vccd1 _13181_/C sky130_fd_sc_hd__nor2_1
XANTENNA__15477__B1 _15527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11750__A2 _11740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12117_ _17133_/C _19709_/A _19165_/C _18849_/C vssd1 vssd1 vccd1 vccd1 _12117_/Y
+ sky130_fd_sc_hd__nand4_1
X_17974_ _19967_/C _20133_/B _17974_/C _17974_/D vssd1 vssd1 vccd1 vccd1 _17986_/D
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19207__A2 _11841_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13097_ _13133_/C vssd1 vssd1 vccd1 vccd1 _20583_/A sky130_fd_sc_hd__buf_4
XFILLER_69_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19713_ _19713_/A _19713_/B _19713_/C vssd1 vssd1 vccd1 vccd1 _19716_/B sky130_fd_sc_hd__nand3_1
X_16925_ _17133_/A vssd1 vssd1 vccd1 vccd1 _17391_/B sky130_fd_sc_hd__clkbuf_2
X_12048_ _11975_/Y _11976_/Y _12035_/Y _12047_/Y vssd1 vssd1 vccd1 vccd1 _12205_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15229__B1 _14834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19644_ _19575_/A _19575_/B _19578_/A _19643_/Y vssd1 vssd1 vccd1 vccd1 _19686_/A
+ sky130_fd_sc_hd__a31o_1
X_16856_ _16856_/A _16856_/B _16856_/C _16856_/D vssd1 vssd1 vccd1 vccd1 _16856_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_133_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15807_ _15807_/A vssd1 vssd1 vccd1 vccd1 _17860_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11582__B _23590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19575_ _19575_/A _19575_/B _19578_/A _19578_/B vssd1 vssd1 vccd1 vccd1 _19734_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16787_ _16752_/Y _16787_/B _16787_/C vssd1 vssd1 vccd1 vccd1 _17026_/B sky130_fd_sc_hd__nand3b_2
X_13999_ _14331_/A _14790_/B _14331_/C _14149_/A _14796_/B vssd1 vssd1 vccd1 vccd1
+ _14002_/A sky130_fd_sc_hd__a32o_1
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20895__B _23299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18526_ _12483_/Y _12484_/Y _18524_/Y _18525_/X vssd1 vssd1 vccd1 vccd1 _18526_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ _15738_/A vssd1 vssd1 vccd1 vccd1 _15862_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20525__A1 _12674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21072__A _21072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18457_ _19803_/A _18453_/X _19969_/A _16526_/A _18634_/A vssd1 vssd1 vccd1 vccd1
+ _18458_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_34_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15669_ _17233_/A _16198_/C _17766_/B vssd1 vssd1 vccd1 vccd1 _15669_/X sky130_fd_sc_hd__and3_1
XANTENNA__16166__A _19381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17941__A2 _18208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17408_ _17642_/A vssd1 vssd1 vccd1 vccd1 _17408_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12215__B1 _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18388_ _18388_/A _18388_/B _18413_/A _18388_/D vssd1 vssd1 vccd1 vccd1 _18392_/A
+ sky130_fd_sc_hd__or4_1
XANTENNA__15952__A1 _15742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17339_ _17298_/B _17126_/X _17127_/Y _17128_/Y vssd1 vssd1 vccd1 vccd1 _17339_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_bq_clk_i clkbuf_2_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_20350_ _20359_/C _20359_/D vssd1 vssd1 vccd1 vccd1 _20352_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19196__B _19196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19009_ _18872_/A _18871_/Y _18844_/D vssd1 vssd1 vccd1 vccd1 _19148_/B sky130_fd_sc_hd__o21ai_2
XFILLER_175_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20281_ _20264_/X _20231_/C _20279_/X _20280_/Y vssd1 vssd1 vccd1 vccd1 _20285_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17457__A1 _17285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22020_ _22144_/A _22020_/B _22144_/C _22021_/A vssd1 vssd1 vccd1 vccd1 _22026_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_115_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17209__A1 _17943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22922_ _22922_/A vssd1 vssd1 vccd1 vccd1 _23296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22853_ _22847_/Y _22850_/Y _22852_/Y vssd1 vssd1 vccd1 vccd1 _22856_/B sky130_fd_sc_hd__a21boi_4
XFILLER_72_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21804_ _21804_/A _21804_/B vssd1 vssd1 vccd1 vccd1 _21805_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12454__B1 _18511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22784_ _22784_/A _22820_/B vssd1 vssd1 vccd1 vccd1 _22786_/A sky130_fd_sc_hd__nor2_2
XANTENNA__13651__C1 _22226_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19382__A1 _19380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21735_ _23328_/Q _21745_/A vssd1 vssd1 vccd1 vccd1 _21898_/C sky130_fd_sc_hd__nand2_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21666_ _21666_/A _21666_/B vssd1 vssd1 vccd1 vccd1 _21666_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23405_ _23409_/CLK _23405_/D vssd1 vssd1 vccd1 vccd1 _23405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20617_ _20597_/C _20614_/Y _20615_/Y _20616_/Y vssd1 vssd1 vccd1 vccd1 _20751_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_138_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21597_ _21597_/A _21597_/B vssd1 vssd1 vccd1 vccd1 _21641_/B sky130_fd_sc_hd__nor2_2
XFILLER_193_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23336_ _23336_/CLK _23336_/D vssd1 vssd1 vccd1 vccd1 _23336_/Q sky130_fd_sc_hd__dfxtp_1
X_20548_ _20548_/A vssd1 vssd1 vccd1 vccd1 _20553_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16523__B _16523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23267_ _23584_/CLK _23267_/D vssd1 vssd1 vccd1 vccd1 _23267_/Q sky130_fd_sc_hd__dfxtp_4
X_20479_ _20479_/A vssd1 vssd1 vccd1 vccd1 _20479_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13020_ _23296_/Q vssd1 vssd1 vccd1 vccd1 _20481_/B sky130_fd_sc_hd__buf_4
XANTENNA__12770__C _12770_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22218_ _22218_/A _22218_/B vssd1 vssd1 vccd1 vccd1 _22220_/A sky130_fd_sc_hd__nand2_1
XFILLER_152_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23198_ _15674_/C input34/X _23206_/S vssd1 vssd1 vccd1 vccd1 _23199_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17635__A _17635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16120__A1 _15971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22149_ _22474_/C _22160_/B _22162_/B vssd1 vssd1 vccd1 vccd1 _22149_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_95 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input37_A wb_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14971_ _23363_/Q _15115_/B _15115_/C vssd1 vssd1 vccd1 vccd1 _15171_/A sky130_fd_sc_hd__nand3b_1
XFILLER_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16710_ _16710_/A vssd1 vssd1 vccd1 vccd1 _16712_/A sky130_fd_sc_hd__inv_2
X_13922_ _14189_/A _14027_/A _14078_/A _13922_/D vssd1 vssd1 vccd1 vccd1 _13927_/A
+ sky130_fd_sc_hd__nand4_4
X_17690_ _18207_/A _18208_/A _17538_/X _17527_/C _17945_/B vssd1 vssd1 vccd1 vccd1
+ _17693_/B sky130_fd_sc_hd__o221ai_1
XANTENNA__12693__B1 _12692_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18412__A3 _20317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12498__B _23592_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15226__A3 _15075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16641_ _16641_/A _16641_/B vssd1 vssd1 vccd1 vccd1 _16641_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13853_ _13853_/A _13853_/B _13853_/C vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__nand3_1
XFILLER_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14434__A1 _14068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19360_ _12324_/X _17976_/A _19357_/Y _19614_/B vssd1 vssd1 vccd1 vccd1 _19361_/B
+ sky130_fd_sc_hd__o31ai_2
XFILLER_16_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ _13176_/A _20528_/C _13176_/C vssd1 vssd1 vccd1 vccd1 _12805_/B sky130_fd_sc_hd__nand3_1
X_16572_ _16757_/C _16572_/B vssd1 vssd1 vccd1 vccd1 _16573_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13784_ _13784_/A vssd1 vssd1 vccd1 vccd1 _21744_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18311_ _18302_/A _18254_/B _18254_/C _18154_/A vssd1 vssd1 vccd1 vccd1 _18314_/A
+ sky130_fd_sc_hd__a31o_1
X_15523_ _15503_/A _15503_/B _15502_/A vssd1 vssd1 vccd1 vccd1 _15525_/A sky130_fd_sc_hd__a21oi_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19291_ _19104_/A _19290_/B _19290_/A vssd1 vssd1 vccd1 vccd1 _19291_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12735_ _12634_/X _12722_/X _12733_/A vssd1 vssd1 vccd1 vccd1 _12738_/A sky130_fd_sc_hd__o21ai_1
XFILLER_71_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18242_ _18242_/A _18242_/B vssd1 vssd1 vccd1 vccd1 _18244_/A sky130_fd_sc_hd__nand2_1
XFILLER_176_818 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15934__A1 _16781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15454_ _15424_/A _15424_/C _15424_/B vssd1 vssd1 vccd1 vccd1 _15457_/B sky130_fd_sc_hd__a21boi_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12618_/A _20493_/D _14655_/A vssd1 vssd1 vccd1 vccd1 _12794_/B sky130_fd_sc_hd__o21ai_1
XFILLER_188_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_870 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14405_ _14405_/A _14405_/B _14405_/C vssd1 vssd1 vccd1 vccd1 _14405_/Y sky130_fd_sc_hd__nand3_1
X_11617_ _12100_/C vssd1 vssd1 vccd1 vccd1 _18798_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_187_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18173_ _18219_/D _18101_/B _18217_/A _18172_/X vssd1 vssd1 vccd1 vccd1 _18173_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13122__B _13122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15385_ _15330_/A _15329_/A _15328_/Y _15383_/X _15384_/Y vssd1 vssd1 vccd1 vccd1
+ _15385_/Y sky130_fd_sc_hd__o2111ai_4
X_12597_ _12601_/A _12601_/C _12601_/B vssd1 vssd1 vccd1 vccd1 _13052_/A sky130_fd_sc_hd__a21o_2
XFILLER_7_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17124_ _17124_/A _17124_/B vssd1 vssd1 vccd1 vccd1 _17125_/B sky130_fd_sc_hd__nand2_1
XFILLER_128_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23209__A0 _15605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14336_ _14793_/C vssd1 vssd1 vccd1 vccd1 _15075_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_144_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17055_ _17055_/A vssd1 vssd1 vccd1 vccd1 _17443_/A sky130_fd_sc_hd__buf_2
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14267_ _14086_/B _14094_/X _14863_/A _14108_/Y vssd1 vssd1 vccd1 vccd1 _14267_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_109_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17248__C _17248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13218_ _23333_/Q vssd1 vssd1 vccd1 vccd1 _22018_/A sky130_fd_sc_hd__buf_2
XFILLER_48_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16006_ _16248_/A _16249_/B vssd1 vssd1 vccd1 vccd1 _16006_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14198_ _13942_/X _14107_/A _14197_/Y vssd1 vssd1 vccd1 vccd1 _14934_/A sky130_fd_sc_hd__o21ai_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17545__A _19675_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13196_/B _13135_/B _13129_/X _13136_/Y vssd1 vssd1 vccd1 vccd1 _13149_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13792__B _22064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17957_ _17928_/A _17928_/B _17836_/Y vssd1 vssd1 vccd1 vccd1 _17957_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18939__A1 _18755_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16908_ _16908_/A vssd1 vssd1 vccd1 vccd1 _16908_/X sky130_fd_sc_hd__clkbuf_2
X_17888_ _17888_/A _18016_/B _19957_/A _18016_/D vssd1 vssd1 vccd1 vccd1 _18017_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_38_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19627_ _19638_/A _19627_/B _19638_/B _19638_/C vssd1 vssd1 vccd1 vccd1 _19627_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__16414__A2 _16408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16839_ _16822_/X _16838_/Y _17073_/A vssd1 vssd1 vccd1 vccd1 _16839_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18376__A _20366_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23589__CLK _23598_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19558_ _12243_/X _17763_/A _19119_/Y _19547_/X vssd1 vssd1 vccd1 vccd1 _19558_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18509_ _18500_/X _11926_/X _18508_/Y vssd1 vssd1 vccd1 vccd1 _18510_/D sky130_fd_sc_hd__o21ai_1
X_19489_ _11926_/X _19668_/A _19486_/A vssd1 vssd1 vccd1 vccd1 _19492_/A sky130_fd_sc_hd__o21ai_1
XFILLER_181_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21520_ _21521_/B _21521_/A vssd1 vssd1 vccd1 vccd1 _21570_/A sky130_fd_sc_hd__and2_1
XANTENNA__17390__A3 _17324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21451_ _21510_/B _21510_/C _21510_/A vssd1 vssd1 vccd1 vccd1 _21463_/A sky130_fd_sc_hd__a21o_1
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20402_ _20428_/B _20428_/C _20401_/X vssd1 vssd1 vccd1 vccd1 _20403_/B sky130_fd_sc_hd__o21bai_1
XFILLER_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19000__A _19163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21382_ _21383_/B _21383_/C _21383_/A vssd1 vssd1 vccd1 vccd1 _21391_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20146__A _20146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15689__B1 _15664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23121_ _11743_/A input32/X _23123_/S vssd1 vssd1 vccd1 vccd1 _23122_/A sky130_fd_sc_hd__mux2_1
X_20333_ _20287_/C _20332_/X _20284_/X vssd1 vssd1 vccd1 vccd1 _20363_/B sky130_fd_sc_hd__a21boi_2
XFILLER_190_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16062__C _16073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23052_ _23052_/A vssd1 vssd1 vccd1 vccd1 _23354_/D sky130_fd_sc_hd__clkbuf_1
X_20264_ _20221_/X _20223_/Y _18001_/X _20368_/D _20164_/B vssd1 vssd1 vccd1 vccd1
+ _20264_/X sky130_fd_sc_hd__a2111o_1
XFILLER_1_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22361__A _22564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__D _16141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22003_ _13642_/X _22420_/B _22420_/C _21922_/A _21922_/B vssd1 vssd1 vccd1 vccd1
+ _22003_/X sky130_fd_sc_hd__o32a_1
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17455__A _17845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13983__A _23502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16102__A1 _16089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20195_ _19775_/Y _19782_/X _19783_/X vssd1 vssd1 vccd1 vccd1 _20196_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12599__A _23449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17605__D _20055_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19670__A _19670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22905_ _12678_/C input32/X _22907_/S vssd1 vssd1 vccd1 vccd1 _22906_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22836_ _22836_/A _22836_/B vssd1 vssd1 vccd1 vccd1 _22836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22767_ _22710_/A _22709_/A _22800_/C _22766_/Y vssd1 vssd1 vccd1 vccd1 _22767_/X
+ sky130_fd_sc_hd__o31a_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_695 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ _18540_/C _12520_/B vssd1 vssd1 vccd1 vccd1 _12522_/C sky130_fd_sc_hd__or2_2
XFILLER_72_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21718_ _21716_/X _21711_/B _21717_/Y _21723_/B vssd1 vssd1 vccd1 vccd1 _21719_/B
+ sky130_fd_sc_hd__o31ai_1
XFILLER_9_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22698_ _22537_/X _22729_/C _22697_/X vssd1 vssd1 vccd1 vccd1 _22698_/Y sky130_fd_sc_hd__o21bai_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12443_/B _12443_/C _12443_/A vssd1 vssd1 vccd1 vccd1 _12451_/Y sky130_fd_sc_hd__a21oi_2
X_21649_ _21666_/A _21666_/B _21649_/C vssd1 vssd1 vccd1 vccd1 _21650_/B sky130_fd_sc_hd__nand3_1
XFILLER_185_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15170_ _15316_/A _15317_/A _15238_/C vssd1 vssd1 vccd1 vccd1 _15170_/Y sky130_fd_sc_hd__nand3_2
XFILLER_138_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12382_ _12363_/B _12376_/X _12381_/X vssd1 vssd1 vccd1 vccd1 _12382_/X sky130_fd_sc_hd__o21ba_1
XFILLER_138_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14121_ _14121_/A _14121_/B vssd1 vssd1 vccd1 vccd1 _14121_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23319_ input5/X _23319_/D vssd1 vssd1 vccd1 vccd1 _23319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ _14017_/X _14050_/X _15085_/C vssd1 vssd1 vccd1 vccd1 _14911_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__18618__B1 _18617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_21 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13003_ _20473_/A _13003_/B _20473_/C vssd1 vssd1 vccd1 vccd1 _13003_/Y sky130_fd_sc_hd__nand3_1
XFILLER_134_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18860_ _18952_/D _19664_/B _18677_/Y _18859_/X vssd1 vssd1 vccd1 vccd1 _18862_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_106_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17811_ _17806_/B _17810_/X _17805_/A _17805_/B vssd1 vssd1 vccd1 vccd1 _17924_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__23517__D input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17841__A1 _17742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18791_ _18475_/A _18484_/A _18973_/C _18478_/A vssd1 vssd1 vccd1 vccd1 _18971_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17742_ _17742_/A vssd1 vssd1 vccd1 vccd1 _17742_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_130_1011 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14954_ _14954_/A _14954_/B vssd1 vssd1 vccd1 vccd1 _14957_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12666__B1 _14655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1085 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13905_ _23352_/Q vssd1 vssd1 vccd1 vccd1 _14023_/C sky130_fd_sc_hd__inv_2
XFILLER_78_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17673_ _17673_/A _17673_/B vssd1 vssd1 vccd1 vccd1 _17705_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14885_ _14753_/Y _14760_/X _14756_/Y vssd1 vssd1 vccd1 vccd1 _14885_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19412_ _19254_/A _19245_/A _19257_/Y _19256_/X vssd1 vssd1 vccd1 vccd1 _19413_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_16624_ _17249_/A _17250_/A _16805_/A _16799_/A vssd1 vssd1 vccd1 vccd1 _16812_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13836_ _13836_/A _13842_/A vssd1 vssd1 vccd1 vccd1 _13839_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _19350_/A _19325_/Y _19339_/X _19342_/Y vssd1 vssd1 vccd1 vccd1 _19471_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_16555_ _16531_/A _16544_/Y _16543_/X _16553_/X _16554_/Y vssd1 vssd1 vccd1 vccd1
+ _16555_/Y sky130_fd_sc_hd__a32oi_2
XFILLER_62_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13767_ _13520_/A _13256_/A _13766_/Y vssd1 vssd1 vccd1 vccd1 _13767_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_189_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14229__A _14230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15506_ _15499_/A _15498_/A _15497_/Y vssd1 vssd1 vccd1 vccd1 _15521_/B sky130_fd_sc_hd__o21a_1
XFILLER_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19274_ _19442_/A _19106_/B _19268_/X _19273_/Y vssd1 vssd1 vccd1 vccd1 _19294_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_12718_ _12718_/A _12718_/B _12718_/C vssd1 vssd1 vccd1 vccd1 _13138_/D sky130_fd_sc_hd__nand3_2
XFILLER_149_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11641__B2 _19196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16486_ _16763_/B vssd1 vssd1 vccd1 vccd1 _16486_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20900__A1 _12674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21988__C _21992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13698_ _13698_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13698_/Y sky130_fd_sc_hd__nand2_1
X_18225_ _18223_/X _18225_/B vssd1 vssd1 vccd1 vccd1 _18226_/B sky130_fd_sc_hd__and2b_1
X_15437_ _15437_/A _15437_/B vssd1 vssd1 vccd1 vccd1 _15438_/B sky130_fd_sc_hd__nand2_2
XFILLER_50_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12649_ _20628_/C vssd1 vssd1 vccd1 vccd1 _20781_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_157_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18156_ _18156_/A _18156_/B vssd1 vssd1 vccd1 vccd1 _18242_/B sky130_fd_sc_hd__nand2_1
XANTENNA__22653__A1 _13547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17259__B _18607_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15368_ _15366_/Y _15365_/X _15360_/X _15308_/D vssd1 vssd1 vccd1 vccd1 _15379_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17107_ _17107_/A _17235_/A _17243_/B vssd1 vssd1 vccd1 vccd1 _17112_/B sky130_fd_sc_hd__and3_1
XANTENNA__20664__B1 _12692_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_748 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14319_ _14459_/D _15356_/A _14459_/A _15082_/D vssd1 vssd1 vccd1 vccd1 _14319_/Y
+ sky130_fd_sc_hd__a22oi_4
X_18087_ _20217_/A _17960_/B _18016_/D _18079_/A _20215_/A vssd1 vssd1 vccd1 vccd1
+ _18088_/C sky130_fd_sc_hd__a32o_1
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15299_ _15299_/A _15299_/B vssd1 vssd1 vccd1 vccd1 _15388_/B sky130_fd_sc_hd__nor2_1
XFILLER_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17038_ _17249_/A _17250_/A _15968_/A _17569_/A vssd1 vssd1 vccd1 vccd1 _17039_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_144_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19806__C1 _20055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12354__C1 _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19193__C _19193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22169__B1 _22280_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater100 _23503_/Q vssd1 vssd1 vccd1 vccd1 _14797_/B sky130_fd_sc_hd__clkbuf_2
X_18989_ _18989_/A _18989_/B vssd1 vssd1 vccd1 vccd1 _19509_/A sky130_fd_sc_hd__nand2_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater111 _23300_/CLK vssd1 vssd1 vccd1 vccd1 _23298_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater122 _23381_/CLK vssd1 vssd1 vccd1 vccd1 _23397_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater133 _23359_/CLK vssd1 vssd1 vccd1 vccd1 _23363_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater144 _23377_/CLK vssd1 vssd1 vccd1 vccd1 _23437_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater155 _23327_/CLK vssd1 vssd1 vccd1 vccd1 _23430_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20951_ _20984_/B _20984_/C vssd1 vssd1 vccd1 vccd1 _20977_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17596__B1 _17605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16619__A _16619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20882_ _20882_/A _20882_/B vssd1 vssd1 vccd1 vccd1 _20883_/A sky130_fd_sc_hd__and2_1
XANTENNA__11880__A1 _11799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22621_ _23278_/Q vssd1 vssd1 vccd1 vccd1 _22623_/A sky130_fd_sc_hd__inv_2
XFILLER_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22552_ _22550_/Y _22551_/Y _22501_/A vssd1 vssd1 vccd1 vccd1 _22589_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__19649__B _19649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21503_ _21502_/B _21502_/C _21635_/A _20786_/Y vssd1 vssd1 vccd1 vccd1 _21504_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_166_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22483_ _22493_/A vssd1 vssd1 vccd1 vccd1 _22545_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18272__C _19425_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21434_ _21359_/B _21635_/C _21431_/X _21433_/Y vssd1 vssd1 vccd1 vccd1 _21434_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_181_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16073__B _16073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19087__D _19263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21365_ _21365_/A vssd1 vssd1 vccd1 vccd1 _21386_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23104_ _23378_/Q input27/X _23106_/S vssd1 vssd1 vccd1 vccd1 _23105_/A sky130_fd_sc_hd__mux2_1
X_20316_ _18211_/A _20365_/A _20269_/B _18324_/A vssd1 vssd1 vccd1 vccd1 _20322_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19384__B _19568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21296_ _20906_/X _20907_/X _21302_/A _20908_/X vssd1 vssd1 vccd1 vccd1 _21296_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23035_ _23035_/A vssd1 vssd1 vccd1 vccd1 _23347_/D sky130_fd_sc_hd__clkbuf_1
X_20247_ _20252_/C _20247_/B _20252_/A vssd1 vssd1 vccd1 vccd1 _20307_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__20958__A1 _20957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19812__A2 _12518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16087__B1 _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20958__B2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17823__A1 _17535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17284__C1 _17974_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_86 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20178_ _20173_/Y _20176_/Y _20177_/Y vssd1 vssd1 vccd1 vccd1 _20181_/A sky130_fd_sc_hd__a21oi_2
XFILLER_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14637__A1 _23331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14637__B2 _23299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13218__A _23333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21907__B1 _21913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ _11951_/A vssd1 vssd1 vccd1 vccd1 _11951_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_123_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _23368_/Q _14667_/X _14669_/X vssd1 vssd1 vccd1 vccd1 _14670_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11882_ _11882_/A vssd1 vssd1 vccd1 vccd1 _11882_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19328__A1 _16604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13621_ _13610_/Y _13609_/X _13620_/X vssd1 vssd1 vccd1 vccd1 _13621_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13073__B1 _12902_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22819_ _22783_/B _23281_/Q _22821_/B _22743_/B _22626_/A vssd1 vssd1 vccd1 vccd1
+ _22819_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_77_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13612__A2 _13599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16340_ _16340_/A _16340_/B _16340_/C vssd1 vssd1 vccd1 vccd1 _16340_/Y sky130_fd_sc_hd__nand3_1
X_13552_ _13552_/A vssd1 vssd1 vccd1 vccd1 _22474_/A sky130_fd_sc_hd__buf_2
XFILLER_197_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16547__D1 _16458_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12503_ _12497_/A _17964_/A _11721_/A vssd1 vssd1 vccd1 vccd1 _12514_/B sky130_fd_sc_hd__o21ai_2
XFILLER_185_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13483_ _13264_/C _13483_/B _13483_/C vssd1 vssd1 vccd1 vccd1 _13485_/A sky130_fd_sc_hd__nand3b_2
X_16271_ _16585_/A vssd1 vssd1 vccd1 vccd1 _16281_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_185_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18010_ _12088_/X _18276_/C _17860_/Y _17859_/Y vssd1 vssd1 vccd1 vccd1 _18013_/B
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__12179__A2 _12168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15222_ _15222_/A vssd1 vssd1 vccd1 vccd1 _15222_/Y sky130_fd_sc_hd__inv_2
X_12434_ _12121_/B _11980_/Y _12095_/Y _14646_/A vssd1 vssd1 vccd1 vccd1 _12435_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_138_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23284__CLK _23492_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19500__A1 _16523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19500__B2 _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12365_ _12364_/A _12364_/B _12364_/C vssd1 vssd1 vccd1 vccd1 _12368_/B sky130_fd_sc_hd__a21o_1
XANTENNA__15117__A2 _15233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15153_ _15109_/X _15110_/X _15017_/D _15082_/B _15253_/B vssd1 vssd1 vccd1 vccd1
+ _15267_/C sky130_fd_sc_hd__a32o_1
XFILLER_126_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14104_ _14261_/A vssd1 vssd1 vccd1 vccd1 _14105_/A sky130_fd_sc_hd__inv_2
X_19961_ _19944_/Y _19864_/C _19960_/Y vssd1 vssd1 vccd1 vccd1 _19963_/A sky130_fd_sc_hd__a21oi_2
X_15084_ _15084_/A vssd1 vssd1 vccd1 vccd1 _15488_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12296_ _12266_/Y _12339_/C _12339_/B vssd1 vssd1 vccd1 vccd1 _12298_/B sky130_fd_sc_hd__o21ai_1
XFILLER_113_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18912_ _19090_/A _18912_/B _19090_/C vssd1 vssd1 vccd1 vccd1 _18912_/Y sky130_fd_sc_hd__nand3_1
X_14035_ _14035_/A vssd1 vssd1 vccd1 vccd1 _14790_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_113_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23060__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19892_ _19896_/A _19897_/C vssd1 vssd1 vccd1 vccd1 _19894_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_120 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14512__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18843_ _18647_/C _18647_/A _18647_/B _18669_/C _18665_/C vssd1 vssd1 vccd1 vccd1
+ _18845_/B sky130_fd_sc_hd__a32oi_1
XFILLER_110_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18774_ _18774_/A vssd1 vssd1 vccd1 vccd1 _19073_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15986_ _15986_/A vssd1 vssd1 vccd1 vccd1 _16181_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17725_ _17589_/Y _17719_/X _17720_/Y _17724_/Y vssd1 vssd1 vccd1 vccd1 _17725_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__23036__S _23038_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14937_ _14805_/B _14928_/B _14934_/X vssd1 vssd1 vccd1 vccd1 _14938_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__21374__A1 _13177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17656_ _17656_/A _17656_/B _17656_/C vssd1 vssd1 vccd1 vccd1 _17658_/B sky130_fd_sc_hd__nand3_1
X_14868_ _15111_/B _15112_/C _15112_/D _14868_/D vssd1 vssd1 vccd1 vccd1 _14868_/Y
+ sky130_fd_sc_hd__nand4b_2
XFILLER_90_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19319__A1 _19172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16607_ _16607_/A _16647_/B vssd1 vssd1 vccd1 vccd1 _16655_/B sky130_fd_sc_hd__nand2_1
X_13819_ _13819_/A _13819_/B vssd1 vssd1 vccd1 vccd1 _13819_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17587_ _17587_/A vssd1 vssd1 vccd1 vccd1 _20138_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14799_ _14795_/Y _14796_/Y _14797_/X _14798_/Y vssd1 vssd1 vccd1 vccd1 _14934_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19326_ _18440_/X _18439_/X _19017_/A _19805_/A vssd1 vssd1 vccd1 vccd1 _19482_/A
+ sky130_fd_sc_hd__o211ai_4
X_16538_ _16539_/A _16539_/B _16539_/C vssd1 vssd1 vccd1 vccd1 _16538_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18542__A2 _18524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19257_ _19257_/A _19257_/B vssd1 vssd1 vccd1 vccd1 _19257_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16469_ _16469_/A _16469_/B _16517_/B _16517_/C vssd1 vssd1 vccd1 vccd1 _16483_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19188__C _19188_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20408__B _20408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18208_ _18208_/A vssd1 vssd1 vccd1 vccd1 _18208_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19188_ _19188_/A _19188_/B _19188_/C vssd1 vssd1 vccd1 vccd1 _19189_/A sky130_fd_sc_hd__nand3_1
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18139_ _18139_/A _18139_/B _18139_/C _18139_/D vssd1 vssd1 vccd1 vccd1 _18140_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19485__A _19485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1022 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12207__A _12207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_662 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21150_ _21014_/X _21002_/Y _21148_/Y _21149_/Y vssd1 vssd1 vccd1 vccd1 _21150_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__16621__B _23595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20101_ _20011_/B _20011_/C _20011_/A vssd1 vssd1 vccd1 vccd1 _20102_/B sky130_fd_sc_hd__a21boi_1
XFILLER_132_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23051__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21081_ _21082_/A _21082_/B _21082_/C vssd1 vssd1 vccd1 vccd1 _21083_/A sky130_fd_sc_hd__a21o_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21062__B1 _12692_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20032_ _20032_/A _20032_/B vssd1 vssd1 vccd1 vccd1 _20207_/A sky130_fd_sc_hd__nor2_1
XANTENNA__17266__C1 _17243_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14619__A1 _18997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17733__A _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19558__A1 _12243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20797__C _23298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21983_ _21891_/Y _13553_/X _21892_/X _21798_/C vssd1 vssd1 vccd1 vccd1 _21983_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11781__A _15718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20934_ _20934_/A _20934_/B vssd1 vssd1 vccd1 vccd1 _20940_/C sky130_fd_sc_hd__nand2_1
XFILLER_82_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ _21157_/C vssd1 vssd1 vccd1 vccd1 _20865_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22604_ _22605_/A _22633_/A _22633_/B vssd1 vssd1 vccd1 vccd1 _22631_/A sky130_fd_sc_hd__and3_1
X_23584_ _23584_/CLK _23584_/D vssd1 vssd1 vccd1 vccd1 _23584_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20796_ _20799_/A _20641_/A _21047_/C _21046_/A vssd1 vssd1 vccd1 vccd1 _21036_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_169_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18533__A2 _11852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22535_ _22454_/A _22454_/B _22450_/A vssd1 vssd1 vccd1 vccd1 _22536_/B sky130_fd_sc_hd__o21ai_4
XFILLER_194_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_606 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22466_ _22566_/A _22566_/B vssd1 vssd1 vccd1 vccd1 _22757_/B sky130_fd_sc_hd__nand2_2
XFILLER_120_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21417_ _21411_/A _21411_/B _21410_/Y vssd1 vssd1 vccd1 vccd1 _21418_/C sky130_fd_sc_hd__o21ai_1
XFILLER_182_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22397_ _22288_/B _22288_/A _22289_/B _22395_/Y vssd1 vssd1 vccd1 vccd1 _22400_/D
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__12117__A _17133_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12150_ _19193_/C vssd1 vssd1 vccd1 vccd1 _19700_/B sky130_fd_sc_hd__buf_4
X_21348_ _21542_/A _21341_/Y _21347_/X vssd1 vssd1 vccd1 vccd1 _21349_/B sky130_fd_sc_hd__o21ai_2
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20334__A _20335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16531__B _16558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11956__A _17626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _11916_/X _11947_/C _12070_/Y _11961_/A vssd1 vssd1 vccd1 vccd1 _18600_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21279_ _21369_/A _21370_/A _21279_/C _21279_/D vssd1 vssd1 vccd1 vccd1 _21279_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_151_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23018_ _23018_/A vssd1 vssd1 vccd1 vccd1 _23339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17643__A _17643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15840_ _15852_/A _15843_/A _15759_/X _15754_/X vssd1 vssd1 vccd1 vccd1 _15941_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15771_ _16070_/B _15746_/Y _15760_/Y _15770_/X vssd1 vssd1 vccd1 vccd1 _15890_/A
+ sky130_fd_sc_hd__o2bb2ai_4
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12983_ _12977_/B _12977_/C _12977_/A vssd1 vssd1 vccd1 vccd1 _12984_/B sky130_fd_sc_hd__a21oi_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _17514_/A _17514_/D vssd1 vssd1 vccd1 vccd1 _17510_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11691__A _18849_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _23595_/Q _23596_/Q vssd1 vssd1 vccd1 vccd1 _16795_/B sky130_fd_sc_hd__nor2_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18490_ _18490_/A vssd1 vssd1 vccd1 vccd1 _19499_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _12089_/A _11926_/X _11966_/B vssd1 vssd1 vccd1 vccd1 _11934_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _16479_/X _17733_/A _17433_/X _17437_/X _17580_/A vssd1 vssd1 vccd1 vccd1
+ _17441_/Y sky130_fd_sc_hd__o221ai_4
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21108__A1 _21159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ _22028_/B vssd1 vssd1 vccd1 vccd1 _21853_/A sky130_fd_sc_hd__buf_2
XFILLER_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11865_ _11896_/B vssd1 vssd1 vccd1 vccd1 _11865_/X sky130_fd_sc_hd__buf_4
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _22022_/A _13602_/Y _13603_/X vssd1 vssd1 vccd1 vccd1 _21752_/A sky130_fd_sc_hd__o21bai_4
X_17372_ _17372_/A _17372_/B vssd1 vssd1 vccd1 vccd1 _17698_/A sky130_fd_sc_hd__nor2_1
X_14584_ _13379_/X _14532_/X _14580_/X _14583_/X vssd1 vssd1 vccd1 vccd1 _14584_/X
+ sky130_fd_sc_hd__a211o_1
X_11796_ _11847_/A _11764_/A _12016_/A vssd1 vssd1 vccd1 vccd1 _11803_/A sky130_fd_sc_hd__o21ai_1
X_19111_ _19138_/A _19138_/B _19139_/A vssd1 vssd1 vccd1 vccd1 _19409_/A sky130_fd_sc_hd__a21boi_2
XANTENNA__16706__B _16706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16323_ _16323_/A _16402_/B vssd1 vssd1 vccd1 vccd1 _16323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ _13535_/A _13535_/B vssd1 vssd1 vccd1 vccd1 _13536_/C sky130_fd_sc_hd__nor2_1
XFILLER_186_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14507__A _15964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19042_ _19138_/A _19139_/A _19138_/B vssd1 vssd1 vccd1 vccd1 _19042_/X sky130_fd_sc_hd__and3_1
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13411__A _13804_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16254_ _16254_/A _16254_/B _16254_/C _16254_/D vssd1 vssd1 vccd1 vccd1 _16258_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_173_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13466_ _13466_/A vssd1 vssd1 vccd1 vccd1 _21892_/A sky130_fd_sc_hd__buf_2
XFILLER_12_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21050__D _21050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15205_ _15204_/Y _15080_/X _15134_/B vssd1 vssd1 vccd1 vccd1 _15222_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__12021__A1 _12018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ _11705_/Y _19804_/A _18788_/A _15699_/A vssd1 vssd1 vccd1 vccd1 _12455_/D
+ sky130_fd_sc_hd__nand4b_2
XFILLER_154_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16185_ _16194_/B vssd1 vssd1 vccd1 vccd1 _16662_/A sky130_fd_sc_hd__clkbuf_2
X_13397_ _13620_/C vssd1 vssd1 vccd1 vccd1 _22420_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15136_ _15074_/Y _15136_/B _15136_/C vssd1 vssd1 vccd1 vccd1 _15140_/C sky130_fd_sc_hd__nand3b_1
XFILLER_182_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12348_ _12366_/A _12348_/B _12348_/C vssd1 vssd1 vccd1 vccd1 _12372_/A sky130_fd_sc_hd__nand3_1
XFILLER_99_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15338__A _15338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19944_ _19943_/Y _19860_/X _19656_/B vssd1 vssd1 vccd1 vccd1 _19944_/Y sky130_fd_sc_hd__a21oi_1
X_12279_ _12279_/A vssd1 vssd1 vccd1 vccd1 _12279_/X sky130_fd_sc_hd__buf_4
X_15067_ _15067_/A _15067_/B _15067_/C vssd1 vssd1 vccd1 vccd1 _15067_/X sky130_fd_sc_hd__and3_1
XFILLER_4_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21044__B1 _12634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ _14077_/C _14017_/X _13939_/A _14588_/A vssd1 vssd1 vccd1 vccd1 _14120_/B
+ sky130_fd_sc_hd__o211ai_4
X_19875_ _19939_/A _19876_/B _19833_/X vssd1 vssd1 vccd1 vccd1 _19875_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20898__B _23300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17263__A2 _17587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18826_ _11814_/A _18452_/A _12105_/Y _18835_/A _19029_/A vssd1 vssd1 vccd1 vccd1
+ _18844_/B sky130_fd_sc_hd__o221ai_4
XFILLER_68_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18757_ _18599_/B _18755_/Y _18932_/B _18601_/A vssd1 vssd1 vccd1 vccd1 _18765_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_95_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15969_ _16860_/A _16860_/C _17041_/B _16160_/A vssd1 vssd1 vccd1 vccd1 _15969_/X
+ sky130_fd_sc_hd__and4_2
XANTENNA__12697__A _23451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17708_ _17806_/A _17806_/B _17810_/B vssd1 vssd1 vccd1 vccd1 _17708_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_64_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18688_ _18880_/A _18784_/B vssd1 vssd1 vccd1 vccd1 _18688_/Y sky130_fd_sc_hd__nand2_1
X_17639_ _16408_/X _18002_/A _17634_/A vssd1 vssd1 vccd1 vccd1 _17641_/B sky130_fd_sc_hd__o21ai_1
XFILLER_1_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20650_ _20649_/Y _20646_/Y _20645_/Y _12754_/A vssd1 vssd1 vccd1 vccd1 _20652_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__19199__B _19543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13024__C _20669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19309_ _19309_/A _19309_/B vssd1 vssd1 vccd1 vccd1 _19309_/Y sky130_fd_sc_hd__nand2_1
X_20581_ _20886_/A vssd1 vssd1 vccd1 vccd1 _21493_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22320_ _22319_/Y _22200_/C _22214_/Y _22205_/Y vssd1 vssd1 vccd1 vccd1 _22324_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_143_1087 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22251_ _22455_/A _22445_/B _22247_/Y vssd1 vssd1 vccd1 vccd1 _22252_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__17728__A _19951_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21202_ _21202_/A _21202_/B _21307_/B vssd1 vssd1 vccd1 vccd1 _21206_/A sky130_fd_sc_hd__nand3_1
XFILLER_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22182_ _22560_/A _22560_/B _13430_/A vssd1 vssd1 vccd1 vccd1 _22182_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21133_ _21125_/A _21125_/B _21126_/Y vssd1 vssd1 vccd1 vccd1 _21153_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__19228__B1 _19188_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21064_ _21545_/A _21061_/X _20962_/Y _21062_/X _21063_/Y vssd1 vssd1 vccd1 vccd1
+ _21064_/X sky130_fd_sc_hd__o311a_1
XANTENNA__19662__B _20142_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20015_ _20111_/A _20108_/A _20108_/B vssd1 vssd1 vccd1 vccd1 _20015_/X sky130_fd_sc_hd__a21bo_1
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18203__A1 _18154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20320__C _20320_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21966_ _22117_/D _21981_/B _21842_/A vssd1 vssd1 vccd1 vccd1 _21968_/A sky130_fd_sc_hd__a21boi_1
XFILLER_27_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16214__B1 _17753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _20917_/A vssd1 vssd1 vccd1 vccd1 _21358_/B sky130_fd_sc_hd__buf_2
X_21897_ _23330_/Q vssd1 vssd1 vccd1 vccd1 _22029_/A sky130_fd_sc_hd__inv_2
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16807__A _16807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11650_ _11739_/A vssd1 vssd1 vccd1 vccd1 _11721_/A sky130_fd_sc_hd__buf_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ _20770_/X _20772_/X _20776_/A vssd1 vssd1 vccd1 vccd1 _20849_/B sky130_fd_sc_hd__o21a_1
XANTENNA__21432__B _21432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11581_ _11648_/A _11918_/B _11624_/A _11593_/C vssd1 vssd1 vccd1 vccd1 _11582_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_23_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20779_ _20625_/B _20778_/A _20627_/Y vssd1 vssd1 vccd1 vccd1 _20779_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23567_ _23571_/CLK _23567_/D vssd1 vssd1 vccd1 vccd1 _23567_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_11_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13231__A _23333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13320_ _13320_/A vssd1 vssd1 vccd1 vccd1 _13320_/X sky130_fd_sc_hd__clkbuf_2
X_22518_ _22521_/C _22521_/A _22419_/Y _22756_/C _22517_/Y vssd1 vssd1 vccd1 vccd1
+ _22607_/B sky130_fd_sc_hd__a41o_1
XFILLER_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23498_ _23499_/CLK _23498_/D vssd1 vssd1 vccd1 vccd1 _23498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13251_ _23320_/Q _13259_/A _13224_/B _13394_/B _13253_/A vssd1 vssd1 vccd1 vccd1
+ _13660_/C sky130_fd_sc_hd__o311ai_4
X_22449_ _22447_/A _22447_/B _23276_/Q vssd1 vssd1 vccd1 vccd1 _22450_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__15740__A2 _17626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22263__B _22263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ _12387_/A _12387_/B _12059_/D vssd1 vssd1 vccd1 vccd1 _12203_/C sky130_fd_sc_hd__o21ai_2
XFILLER_89_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13182_ _13168_/B _13186_/C _20775_/A _13180_/X _13181_/X vssd1 vssd1 vccd1 vccd1
+ _13191_/D sky130_fd_sc_hd__a41o_1
XFILLER_182_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12133_ _11882_/A _11883_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _12133_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__23015__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17990_ _18157_/D _18157_/B _17960_/X vssd1 vssd1 vccd1 vccd1 _17990_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16941_ _16948_/B _16948_/C _16948_/A vssd1 vssd1 vccd1 vccd1 _16941_/Y sky130_fd_sc_hd__a21oi_1
X_12064_ _12388_/B _12064_/B _12064_/C vssd1 vssd1 vccd1 vccd1 _12391_/C sky130_fd_sc_hd__nand3b_2
XFILLER_81_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19660_ _11936_/X _19499_/A _19659_/Y vssd1 vssd1 vccd1 vccd1 _19674_/C sky130_fd_sc_hd__o21ai_2
X_16872_ _15882_/X _16382_/A _16871_/X _16601_/B vssd1 vssd1 vccd1 vccd1 _16873_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_38_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18611_ _18534_/Y _18607_/X _18532_/Y vssd1 vssd1 vccd1 vccd1 _18615_/A sky130_fd_sc_hd__a21boi_2
XANTENNA__16453__B1 _16356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12013__C _12306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18993__A2 _16033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_bq_clk_i clkbuf_3_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_15823_ _15699_/Y _15785_/A _16451_/B _15822_/X vssd1 vssd1 vccd1 vccd1 _16020_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_19591_ _19587_/X _19589_/X _19590_/Y vssd1 vssd1 vccd1 vccd1 _19592_/C sky130_fd_sc_hd__o21ai_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _12478_/B _18524_/B _18721_/A _18721_/B vssd1 vssd1 vccd1 vccd1 _18902_/B
+ sky130_fd_sc_hd__a211oi_2
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15754_/A vssd1 vssd1 vccd1 vccd1 _15754_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12310__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ _20669_/C vssd1 vssd1 vccd1 vccd1 _21079_/A sky130_fd_sc_hd__buf_2
XANTENNA__20001__A1 _19941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _23408_/Q _14693_/X _14698_/X _23440_/Q _14704_/X vssd1 vssd1 vccd1 vccd1
+ _14705_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ _18473_/A vssd1 vssd1 vccd1 vccd1 _18473_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11917_ _23589_/Q _23590_/Q vssd1 vssd1 vccd1 vccd1 _16141_/A sky130_fd_sc_hd__nor2_4
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16756__A1 _16757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15685_ _15685_/A vssd1 vssd1 vccd1 vccd1 _15686_/B sky130_fd_sc_hd__clkbuf_4
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12900_/A _13034_/A _12893_/Y _12894_/X vssd1 vssd1 vccd1 vccd1 _12901_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_178_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17424_ _17959_/B _19949_/D _17959_/A vssd1 vssd1 vccd1 vccd1 _17425_/B sky130_fd_sc_hd__and3_1
XANTENNA__18508__A1_N _18675_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _22968_/D vssd1 vssd1 vccd1 vccd1 _14636_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11848_ _11848_/A vssd1 vssd1 vccd1 vccd1 _11848_/X sky130_fd_sc_hd__buf_4
XFILLER_159_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17200_/B _17354_/Y _17200_/C vssd1 vssd1 vccd1 vccd1 _17357_/A sky130_fd_sc_hd__o21ai_1
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14567_ _15762_/A _14516_/X _14564_/X _14566_/X vssd1 vssd1 vccd1 vccd1 _14567_/X
+ sky130_fd_sc_hd__o22a_1
X_11779_ _11882_/A _11883_/A vssd1 vssd1 vccd1 vccd1 _18972_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_787 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16306_ _16306_/A vssd1 vssd1 vccd1 vccd1 _16323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13518_ _13517_/A _13517_/C _13517_/B vssd1 vssd1 vccd1 vccd1 _13519_/C sky130_fd_sc_hd__a21o_1
XFILLER_186_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17286_ _12088_/A _17285_/X _17260_/A _17260_/B _17265_/Y vssd1 vssd1 vccd1 vccd1
+ _17286_/X sky130_fd_sc_hd__o221a_1
XFILLER_118_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21996__C _22510_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14498_ _14498_/A _14498_/B vssd1 vssd1 vccd1 vccd1 _14847_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19025_ _17627_/A _11670_/X _19020_/Y _19018_/X vssd1 vssd1 vccd1 vccd1 _19026_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_162_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ _16237_/A vssd1 vssd1 vccd1 vccd1 _16251_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23254__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13449_ _23475_/Q vssd1 vssd1 vccd1 vccd1 _21921_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_127_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12980__A _12980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16168_ _16174_/C _16174_/B _16168_/C vssd1 vssd1 vccd1 vccd1 _16169_/C sky130_fd_sc_hd__nand3_1
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11596__A _19327_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23006__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15119_ _15319_/C _15109_/X _15110_/X _15120_/A _15120_/D vssd1 vssd1 vccd1 vccd1
+ _15164_/A sky130_fd_sc_hd__a32o_1
XFILLER_170_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16099_ _16424_/A _16424_/B vssd1 vssd1 vccd1 vccd1 _16099_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19927_ _19613_/Y _19638_/Y _19768_/A vssd1 vssd1 vccd1 vccd1 _19929_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__20702__A _20775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17283__A _20049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19858_ _19858_/A vssd1 vssd1 vccd1 vccd1 _19953_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16444__B1 _16225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18809_ _18844_/D vssd1 vssd1 vccd1 vccd1 _18872_/B sky130_fd_sc_hd__buf_2
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19789_ _19636_/Y _19459_/B _19788_/Y vssd1 vssd1 vccd1 vccd1 _19789_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__20791__A2 _20786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21820_ _21820_/A _21820_/B vssd1 vssd1 vccd1 vccd1 _21824_/C sky130_fd_sc_hd__xor2_1
XFILLER_37_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21751_ _13793_/B _21906_/A _21750_/Y vssd1 vssd1 vccd1 vccd1 _21753_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__16049__D _16049_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20543__A2 _13184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20702_ _20775_/A _23456_/Q vssd1 vssd1 vccd1 vccd1 _20702_/Y sky130_fd_sc_hd__nand2_1
XFILLER_196_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21682_ _21666_/Y _21647_/Y _21646_/A _21673_/Y vssd1 vssd1 vccd1 vccd1 _21704_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_52_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20633_ _20475_/B _20783_/A _20793_/A _20627_/Y vssd1 vssd1 vccd1 vccd1 _20635_/B
+ sky130_fd_sc_hd__o211ai_1
X_23421_ _23424_/CLK _23421_/D vssd1 vssd1 vccd1 vccd1 _23421_/Q sky130_fd_sc_hd__dfxtp_1
X_23352_ _23352_/CLK _23352_/D vssd1 vssd1 vccd1 vccd1 _23352_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13981__A1 _13972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20564_ _13055_/X _13060_/X _13061_/Y _13070_/B vssd1 vssd1 vccd1 vccd1 _20565_/A
+ sky130_fd_sc_hd__o31ai_1
XFILLER_20_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22364__A _22487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22303_ _22012_/Y _22171_/Y _22302_/X _22173_/Y vssd1 vssd1 vccd1 vccd1 _22303_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_109_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23283_ _23510_/CLK _23283_/D vssd1 vssd1 vccd1 vccd1 _23283_/Q sky130_fd_sc_hd__dfxtp_1
X_20495_ _20495_/A _23297_/Q _20495_/C vssd1 vssd1 vccd1 vccd1 _20782_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12890__A _13052_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22234_ _22234_/A _22234_/B _22234_/C vssd1 vssd1 vccd1 vccd1 _22234_/Y sky130_fd_sc_hd__nand3_1
XFILLER_118_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22165_ _22474_/A _22754_/B _22040_/B _22271_/A _22160_/Y vssd1 vssd1 vccd1 vccd1
+ _22166_/C sky130_fd_sc_hd__o221ai_4
XFILLER_182_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21116_ _21159_/A _21228_/A _21159_/B vssd1 vssd1 vccd1 vccd1 _21119_/A sky130_fd_sc_hd__a21o_1
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22096_ _22830_/B _22096_/B _22096_/C vssd1 vssd1 vccd1 vccd1 _22096_/X sky130_fd_sc_hd__or3_1
XFILLER_160_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17227__A2 _17409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21047_ _21047_/A _21047_/B _21047_/C vssd1 vssd1 vccd1 vccd1 _21048_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19621__B1 _18373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12820_ _12622_/X _12624_/X _12765_/A vssd1 vssd1 vccd1 vccd1 _12820_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22998_ _22998_/A vssd1 vssd1 vccd1 vccd1 _23330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18727__A2 _18723_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12751_ _20473_/C vssd1 vssd1 vccd1 vccd1 _20962_/C sky130_fd_sc_hd__buf_2
XANTENNA__12472__B2 _12093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21949_ _21936_/Y _21941_/Y _21890_/X _21894_/X vssd1 vssd1 vccd1 vccd1 _21949_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_27_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16738__B2 _16724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11702_ _11610_/C _11606_/X _11773_/C _11677_/X vssd1 vssd1 vccd1 vccd1 _11704_/A
+ sky130_fd_sc_hd__o211ai_1
X_15470_ _15471_/A _15501_/A _15471_/C vssd1 vssd1 vccd1 vccd1 _15472_/A sky130_fd_sc_hd__a21o_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _23291_/Q _12873_/C _23292_/Q vssd1 vssd1 vccd1 vccd1 _12682_/Y sky130_fd_sc_hd__nor3_2
XANTENNA__15410__A1 _15225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14213__A2 _14212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14421_ _14422_/B _14422_/C _14422_/A vssd1 vssd1 vccd1 vccd1 _14495_/C sky130_fd_sc_hd__a21o_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12224__A1 _12222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11633_ _23590_/Q vssd1 vssd1 vccd1 vccd1 _11633_/Y sky130_fd_sc_hd__inv_2
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17140_ _17140_/A _17140_/B vssd1 vssd1 vccd1 vccd1 _17140_/Y sky130_fd_sc_hd__nand2_2
XFILLER_11_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14352_ _14420_/A _14352_/B vssd1 vssd1 vccd1 vccd1 _14416_/B sky130_fd_sc_hd__nor2_1
XFILLER_168_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ _13303_/A _13303_/B _13303_/C vssd1 vssd1 vccd1 vccd1 _13538_/B sky130_fd_sc_hd__nor3_2
XFILLER_156_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17071_ _12086_/A _16355_/A _17068_/X _17069_/X _17070_/X vssd1 vssd1 vccd1 vccd1
+ _17071_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14283_ _14358_/C _14349_/C _14349_/D vssd1 vssd1 vccd1 vccd1 _14283_/X sky130_fd_sc_hd__and3_1
XFILLER_183_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16272__A _16275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16022_ _16022_/A vssd1 vssd1 vccd1 vccd1 _16022_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13234_ _22022_/A _13221_/A _13233_/Y vssd1 vssd1 vccd1 vccd1 _13659_/B sky130_fd_sc_hd__o21ai_2
XFILLER_6_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22995__A0 _14614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17466__A2 _17465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ _20773_/C _12979_/A _20773_/A _21440_/B _13158_/A vssd1 vssd1 vccd1 vccd1
+ _13169_/C sky130_fd_sc_hd__a32o_1
XFILLER_156_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18663__B2 _18656_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ _19364_/A vssd1 vssd1 vccd1 vccd1 _19709_/A sky130_fd_sc_hd__clkbuf_4
X_17973_ _19113_/C vssd1 vssd1 vccd1 vccd1 _20133_/B sky130_fd_sc_hd__buf_2
X_13096_ _21455_/B vssd1 vssd1 vccd1 vccd1 _21554_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19712_ _19547_/X _19537_/X _19538_/X _19542_/X vssd1 vssd1 vccd1 vccd1 _19713_/C
+ sky130_fd_sc_hd__a2bb2oi_1
X_16924_ _16935_/A _16930_/B _16922_/Y _16923_/X vssd1 vssd1 vccd1 vccd1 _16924_/Y
+ sky130_fd_sc_hd__o2bb2ai_4
X_12047_ _12015_/Y _12027_/Y _12033_/Y _12049_/A vssd1 vssd1 vccd1 vccd1 _12047_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19612__B1 _19381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1042 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19643_ _19524_/A _19524_/C _19524_/B vssd1 vssd1 vccd1 vccd1 _19643_/Y sky130_fd_sc_hd__a21oi_2
X_16855_ _11853_/A _11921_/Y _17092_/A _16856_/C _16856_/D vssd1 vssd1 vccd1 vccd1
+ _17095_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16977__A1 _16663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12678__C _12678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15806_ _15804_/Y _15621_/X _16213_/A vssd1 vssd1 vccd1 vccd1 _15807_/A sky130_fd_sc_hd__a21boi_2
X_19574_ _19572_/X _19573_/X _19588_/B _19587_/A vssd1 vssd1 vccd1 vccd1 _19574_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16786_ _16198_/X _16194_/Y _16744_/A _16744_/B _16749_/A vssd1 vssd1 vccd1 vccd1
+ _16787_/C sky130_fd_sc_hd__o2111ai_2
XANTENNA__12040__A _18481_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13998_ _14246_/A _14149_/A _14796_/B _14795_/C vssd1 vssd1 vccd1 vccd1 _14003_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_65_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18525_ _12399_/X _12400_/X _12445_/Y _12449_/Y vssd1 vssd1 vccd1 vccd1 _18525_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15737_ _15864_/A _15729_/X _14553_/X vssd1 vssd1 vccd1 vccd1 _15738_/A sky130_fd_sc_hd__o21a_2
X_12949_ _20905_/C _12981_/B _20966_/A _20966_/B vssd1 vssd1 vccd1 vccd1 _12949_/Y
+ sky130_fd_sc_hd__nand4_2
XANTENNA__16447__A _16447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18456_ _18456_/A vssd1 vssd1 vccd1 vccd1 _18634_/A sky130_fd_sc_hd__buf_2
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15668_ _15668_/A vssd1 vssd1 vccd1 vccd1 _17766_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17407_ _16684_/X _16683_/X _11951_/X _11948_/X _17233_/A vssd1 vssd1 vccd1 vccd1
+ _17407_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_18_1130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14619_ _18997_/B _14544_/X _14612_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _14619_/X
+ sky130_fd_sc_hd__a211o_1
X_18387_ _18384_/A _18385_/X _18411_/B vssd1 vssd1 vccd1 vccd1 _18388_/D sky130_fd_sc_hd__a21o_1
XANTENNA__12215__B2 _12214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15952__A2 _16447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15599_ _15715_/A vssd1 vssd1 vccd1 vccd1 _15599_/X sky130_fd_sc_hd__buf_2
XFILLER_53_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17338_ _17337_/A _17337_/B _17331_/A _17331_/B vssd1 vssd1 vccd1 vccd1 _17341_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17154__A1 _12323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11974__B1 _12289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17269_ _16638_/X _16639_/X _16311_/X vssd1 vssd1 vccd1 vccd1 _17269_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19008_ _19043_/A _19044_/A _19007_/Y vssd1 vssd1 vccd1 vccd1 _19148_/A sky130_fd_sc_hd__a21o_1
X_20280_ _20328_/A _20328_/B _20328_/C vssd1 vssd1 vccd1 vccd1 _20280_/Y sky130_fd_sc_hd__nor3_1
XFILLER_162_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22986__A0 _13349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19493__A _19543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17457__A2 _17600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17311__D1 _16529_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20213__A1 _19700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12151__B1 _12149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22921_ _20481_/B input8/X _22929_/S vssd1 vssd1 vccd1 vccd1 _22922_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18837__A _19703_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14979__B1 _14089_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22852_ _22845_/Y _22848_/Y _22851_/Y vssd1 vssd1 vccd1 vccd1 _22852_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15640__A1 _11864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21803_ _21805_/C _21805_/B _21804_/A _21804_/B vssd1 vssd1 vccd1 vccd1 _21803_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12454__A1 _19512_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13651__B1 _22553_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22783_ _23281_/Q _22783_/B vssd1 vssd1 vccd1 vccd1 _22820_/B sky130_fd_sc_hd__nor2_1
XANTENNA__22910__A0 _12608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19382__A2 _19381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21734_ _13358_/A _13784_/A _21745_/A vssd1 vssd1 vccd1 vccd1 _21898_/B sky130_fd_sc_hd__o21ai_2
XFILLER_24_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19119__C1 _17595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21665_ _21665_/A _21665_/B vssd1 vssd1 vccd1 vccd1 _21665_/Y sky130_fd_sc_hd__nand2_1
XFILLER_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23404_ _23435_/CLK _23404_/D vssd1 vssd1 vccd1 vccd1 _23404_/Q sky130_fd_sc_hd__dfxtp_1
X_20616_ _12987_/Y _20459_/Y _13202_/A vssd1 vssd1 vccd1 vccd1 _20616_/Y sky130_fd_sc_hd__a21oi_2
X_21596_ _21595_/C _21633_/A _21594_/B _21594_/A vssd1 vssd1 vccd1 vccd1 _21597_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20547_ _20548_/A _20553_/B _20547_/C vssd1 vssd1 vccd1 vccd1 _20547_/X sky130_fd_sc_hd__and3_1
X_23335_ _23429_/CLK _23335_/D vssd1 vssd1 vccd1 vccd1 _23335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16523__C _16523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20478_ _20621_/A vssd1 vssd1 vccd1 vccd1 _20625_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_23266_ _23584_/CLK _23266_/D vssd1 vssd1 vccd1 vccd1 _23266_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22977__A0 _13253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12770__D _21054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22217_ _22208_/X _22209_/X _22210_/Y _22216_/X vssd1 vssd1 vccd1 vccd1 _22231_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_180_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19842__B1 _19494_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23197_ _23254_/S vssd1 vssd1 vccd1 vccd1 _23206_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_193_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22148_ _22569_/A _22270_/C _22569_/C vssd1 vssd1 vccd1 vccd1 _22162_/B sky130_fd_sc_hd__and3_1
XFILLER_117_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22079_ _21936_/B _21994_/Y _21995_/Y _22075_/Y _22078_/Y vssd1 vssd1 vccd1 vccd1
+ _22093_/C sky130_fd_sc_hd__o2111ai_4
X_14970_ _23362_/Q _14970_/B vssd1 vssd1 vccd1 vccd1 _15115_/C sky130_fd_sc_hd__nand2_1
XFILLER_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18948__A2 _19261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ _23357_/Q _14077_/C vssd1 vssd1 vccd1 vccd1 _13922_/D sky130_fd_sc_hd__nor2_1
XANTENNA__18169__D _18172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16640_ _16638_/X _16639_/X _16064_/A vssd1 vssd1 vccd1 vccd1 _16640_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13852_ _13857_/A _13857_/B vssd1 vssd1 vccd1 vccd1 _13853_/C sky130_fd_sc_hd__nor2_1
XFILLER_90_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22269__A _22566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19358__C1 _17443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14434__A2 _14069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ _13051_/C vssd1 vssd1 vccd1 vccd1 _13176_/C sky130_fd_sc_hd__clkbuf_2
X_16571_ _16759_/B _16759_/C _16763_/B _16570_/Y vssd1 vssd1 vccd1 vccd1 _16768_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13783_ _13783_/A _13783_/B _13783_/C vssd1 vssd1 vccd1 vccd1 _13784_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12795__A _13051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14985__A3 _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22901__A0 _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18310_ _18304_/Y _18306_/Y _18302_/Y _18417_/D vssd1 vssd1 vccd1 vccd1 _18315_/A
+ sky130_fd_sc_hd__o211ai_1
X_15522_ _15522_/A _15522_/B vssd1 vssd1 vccd1 vccd1 _15525_/B sky130_fd_sc_hd__or2_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19290_ _19290_/A _19290_/B vssd1 vssd1 vccd1 vccd1 _19290_/Y sky130_fd_sc_hd__nand2_1
X_12734_ _12734_/A _12734_/B _12734_/C vssd1 vssd1 vccd1 vccd1 _12845_/A sky130_fd_sc_hd__nand3_2
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18241_ _18245_/A _18298_/C _18245_/C vssd1 vssd1 vccd1 vccd1 _18241_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15453_ _15453_/A vssd1 vssd1 vccd1 vccd1 _15462_/B sky130_fd_sc_hd__inv_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _20805_/C vssd1 vssd1 vccd1 vccd1 _13041_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__15934__A2 _15933_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_882 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14404_ _14403_/A _14403_/B _14354_/Y _14355_/X vssd1 vssd1 vccd1 vccd1 _14405_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_18172_ _18172_/A _20151_/C _18172_/C _18172_/D vssd1 vssd1 vccd1 vccd1 _18172_/X
+ sky130_fd_sc_hd__and4_1
X_11616_ _11758_/A vssd1 vssd1 vccd1 vccd1 _12100_/C sky130_fd_sc_hd__buf_2
X_15384_ _15383_/B _15383_/C _15383_/A vssd1 vssd1 vccd1 vccd1 _15384_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__22665__C1 _22664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ _12873_/C vssd1 vssd1 vccd1 vccd1 _12601_/B sky130_fd_sc_hd__clkbuf_4
X_17123_ _17302_/A _17301_/A _17123_/C vssd1 vssd1 vccd1 vccd1 _17124_/B sky130_fd_sc_hd__nand3_1
XANTENNA__17098__A _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14335_ _14381_/A _14381_/B _14333_/X _14334_/Y vssd1 vssd1 vccd1 vccd1 _14353_/B
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__23209__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14515__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17054_ _16625_/X _17252_/A _17039_/Y vssd1 vssd1 vccd1 vccd1 _17058_/A sky130_fd_sc_hd__o21ai_1
XFILLER_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11858__B _11912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14266_ _14429_/A vssd1 vssd1 vccd1 vccd1 _14876_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_171_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17248__D _20317_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16005_ _15946_/Y _15947_/X _16268_/A _15944_/Y vssd1 vssd1 vccd1 vccd1 _16005_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_143_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13217_ _22564_/C vssd1 vssd1 vccd1 vccd1 _22476_/C sky130_fd_sc_hd__buf_2
XANTENNA__18636__A1 _16044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14197_ _14886_/A _14774_/C _14886_/C vssd1 vssd1 vccd1 vccd1 _14197_/Y sky130_fd_sc_hd__nand3_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13148_ _13129_/X _13136_/Y _13135_/Y vssd1 vssd1 vccd1 vccd1 _13148_/X sky130_fd_sc_hd__a21bo_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17956_ _17956_/A vssd1 vssd1 vccd1 vccd1 _23589_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_13079_ _13079_/A _13079_/B vssd1 vssd1 vccd1 vccd1 _13079_/Y sky130_fd_sc_hd__nand2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11593__B _16807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16907_ _16898_/Y _16899_/X _16901_/Y _16906_/Y vssd1 vssd1 vccd1 vccd1 _16935_/A
+ sky130_fd_sc_hd__o211ai_4
X_17887_ _11948_/X _11951_/X _17960_/B vssd1 vssd1 vccd1 vccd1 _18016_/B sky130_fd_sc_hd__o21a_1
XFILLER_38_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19626_ _19613_/Y _19615_/X _19617_/Y vssd1 vssd1 vccd1 vccd1 _19626_/X sky130_fd_sc_hd__o21a_2
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16838_ _16627_/X _17039_/A _16814_/X vssd1 vssd1 vccd1 vccd1 _16838_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__23145__A0 _23396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18376__B _18376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19557_ _12053_/X _12509_/X _19203_/X _17600_/A vssd1 vssd1 vccd1 vccd1 _19557_/X
+ sky130_fd_sc_hd__o22a_1
X_16769_ _17011_/A _17011_/B vssd1 vssd1 vccd1 vccd1 _16776_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18508_ _18675_/C _18504_/Y _18503_/Y _12460_/Y vssd1 vssd1 vccd1 vccd1 _18508_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_181_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19488_ _19577_/A vssd1 vssd1 vccd1 vccd1 _19522_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17375__A1 _17535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18439_ _18439_/A vssd1 vssd1 vccd1 vccd1 _18439_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21450_ _21378_/A _21378_/B _21378_/C _21376_/B vssd1 vssd1 vccd1 vccd1 _21510_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_194_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401_ _20323_/C _20401_/B _20401_/C vssd1 vssd1 vccd1 vccd1 _20401_/X sky130_fd_sc_hd__and3b_1
XFILLER_30_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21381_ _21317_/A _21317_/C _21317_/D _21380_/Y vssd1 vssd1 vccd1 vccd1 _21383_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_147_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20146__B _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20332_ _20210_/C _20366_/A _20314_/X _20265_/B _20287_/B vssd1 vssd1 vccd1 vccd1
+ _20332_/X sky130_fd_sc_hd__o41a_1
X_23120_ _23120_/A vssd1 vssd1 vccd1 vccd1 _23384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_855 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15153__A3 _15017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23051_ _13911_/C input33/X _23051_/S vssd1 vssd1 vccd1 vccd1 _23052_/A sky130_fd_sc_hd__mux2_1
X_20263_ _20263_/A vssd1 vssd1 vccd1 vccd1 _20368_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_116_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22423__A2 _13431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22002_ _21925_/X _21922_/Y _21999_/Y _22001_/Y _21928_/X vssd1 vssd1 vccd1 vccd1
+ _22218_/A sky130_fd_sc_hd__o2111ai_4
XANTENNA__22361__B _22564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13983__B _23501_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20194_ _20207_/A _20117_/X _20196_/C _20193_/Y vssd1 vssd1 vccd1 vccd1 _20199_/B
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__17455__B _17586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_711 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12124__B1 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19670__B _19670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17063__B1 _16840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22904_ _22904_/A vssd1 vssd1 vccd1 vccd1 _23288_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__23533__CLK _23558_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22089__A _22089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22835_ _22834_/B _22834_/C _22834_/A vssd1 vssd1 vccd1 vccd1 _22836_/B sky130_fd_sc_hd__a21oi_1
XFILLER_72_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22766_ _22829_/A _22766_/B vssd1 vssd1 vccd1 vccd1 _22766_/Y sky130_fd_sc_hd__nand2_1
XFILLER_198_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21717_ _21717_/A _21717_/B vssd1 vssd1 vccd1 vccd1 _21717_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16815__A _16815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22697_ _22631_/Y _22683_/B _22683_/A vssd1 vssd1 vccd1 vccd1 _22697_/X sky130_fd_sc_hd__a21bo_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14038__C _14777_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21440__B _21440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ _12399_/X _12400_/X _12445_/Y _12449_/Y vssd1 vssd1 vccd1 vccd1 _12490_/A
+ sky130_fd_sc_hd__o211ai_2
X_21648_ _21632_/Y _21621_/Y _21647_/Y vssd1 vssd1 vccd1 vccd1 _21650_/A sky130_fd_sc_hd__o21ai_1
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12381_ _12381_/A _12381_/B _12381_/C vssd1 vssd1 vccd1 vccd1 _12381_/X sky130_fd_sc_hd__and3_1
X_21579_ _21579_/A _23570_/Q _21579_/C vssd1 vssd1 vccd1 vccd1 _21627_/C sky130_fd_sc_hd__nand3_1
XFILLER_165_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ _14120_/A _14120_/B _14384_/A vssd1 vssd1 vccd1 vccd1 _14121_/B sky130_fd_sc_hd__nand3_4
XFILLER_193_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23318_ _23321_/CLK _23318_/D vssd1 vssd1 vccd1 vccd1 _23318_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21870__B1 _22236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ _14017_/X _14094_/A _14031_/X vssd1 vssd1 vccd1 vccd1 _15085_/C sky130_fd_sc_hd__a21oi_2
XFILLER_4_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23249_ _23249_/A vssd1 vssd1 vccd1 vccd1 _23442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _12712_/X _12704_/A _12694_/A _12726_/Y _20781_/C vssd1 vssd1 vccd1 vccd1
+ _13002_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17810_ _17810_/A _17810_/B _17810_/C _17810_/D vssd1 vssd1 vccd1 vccd1 _17810_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__17841__A2 _17741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19028__D1 _19548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18790_ _18984_/A vssd1 vssd1 vccd1 vccd1 _18790_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17741_ _17741_/A vssd1 vssd1 vccd1 vccd1 _17741_/X sky130_fd_sc_hd__clkbuf_4
X_14953_ _14951_/X _14953_/B _14953_/C vssd1 vssd1 vccd1 vccd1 _14954_/B sky130_fd_sc_hd__nand3b_1
XFILLER_130_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13904_ _14013_/B vssd1 vssd1 vccd1 vccd1 _14191_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_1097 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17672_ _17662_/Y _17669_/X _17671_/X vssd1 vssd1 vccd1 vccd1 _17673_/B sky130_fd_sc_hd__o21ai_1
X_14884_ _15459_/B _14108_/Y _15459_/A _15001_/A _14178_/Y vssd1 vssd1 vccd1 vccd1
+ _14884_/X sky130_fd_sc_hd__o32a_1
X_19411_ _19409_/X _19410_/X _19422_/B _19406_/A vssd1 vssd1 vccd1 vccd1 _19413_/B
+ sky130_fd_sc_hd__o211ai_1
X_16623_ _16817_/A _16819_/A vssd1 vssd1 vccd1 vccd1 _16799_/A sky130_fd_sc_hd__nand2_1
X_13835_ _13820_/Y _13830_/Y _13834_/Y vssd1 vssd1 vccd1 vccd1 _13842_/A sky130_fd_sc_hd__o21ai_1
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12418__A1 _19180_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19342_ _19345_/A _19345_/B _19339_/C vssd1 vssd1 vccd1 vccd1 _19342_/Y sky130_fd_sc_hd__a21oi_1
X_16554_ _16554_/A _16554_/B vssd1 vssd1 vccd1 vccd1 _16554_/Y sky130_fd_sc_hd__nand2_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12969__A2 _12785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ _13766_/A _13766_/B _21883_/B vssd1 vssd1 vccd1 vccd1 _13766_/Y sky130_fd_sc_hd__nand3_1
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15505_ _15527_/B _15505_/B vssd1 vssd1 vccd1 vccd1 _23281_/D sky130_fd_sc_hd__xnor2_1
XFILLER_189_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19273_ _19442_/B vssd1 vssd1 vccd1 vccd1 _19273_/Y sky130_fd_sc_hd__inv_2
X_12717_ _12652_/X _12651_/X _12980_/A _12941_/A _12654_/Y vssd1 vssd1 vccd1 vccd1
+ _12718_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__13133__B _21548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11641__A2 _18675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16485_ _16495_/C _16482_/X _16495_/B vssd1 vssd1 vccd1 vccd1 _16763_/B sky130_fd_sc_hd__a21bo_2
X_13697_ _13697_/A _13697_/B _13697_/C vssd1 vssd1 vccd1 vccd1 _13759_/A sky130_fd_sc_hd__nand3_1
XFILLER_31_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20900__A2 _20471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18224_ _18170_/D _18170_/Y _18220_/X _18222_/X vssd1 vssd1 vccd1 vccd1 _18225_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_15_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21988__D _22663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15436_ _15391_/A _15391_/B _15435_/Y vssd1 vssd1 vccd1 vccd1 _15437_/A sky130_fd_sc_hd__o21ai_1
XFILLER_176_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12648_ _12648_/A vssd1 vssd1 vccd1 vccd1 _12648_/X sky130_fd_sc_hd__buf_2
XANTENNA__17109__B2 _17112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18155_ _18155_/A _18155_/B vssd1 vssd1 vccd1 vccd1 _18192_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14591__A1 _12113_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18857__A1 _11926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15367_ _15308_/D _15360_/X _15365_/X _15366_/Y vssd1 vssd1 vccd1 vccd1 _15379_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_172_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14245__A _14245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12579_ _13011_/C vssd1 vssd1 vccd1 vccd1 _12580_/A sky130_fd_sc_hd__buf_2
XFILLER_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17259__C _18607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17106_ _17106_/A _17106_/B _17106_/C vssd1 vssd1 vccd1 vccd1 _17118_/B sky130_fd_sc_hd__nand3_1
XANTENNA__20664__A1 _20639_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16868__B1 _15991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14318_ _14407_/C _15120_/B _14459_/A vssd1 vssd1 vccd1 vccd1 _14318_/Y sky130_fd_sc_hd__nand3_1
X_18086_ _12506_/A _12506_/B _18002_/A _17959_/Y vssd1 vssd1 vccd1 vccd1 _18088_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16332__A2 _16089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15298_ _15298_/A _15298_/B _15350_/C vssd1 vssd1 vccd1 vccd1 _15299_/B sky130_fd_sc_hd__and3_1
XFILLER_85_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17037_ _16953_/A _16953_/B _16953_/C _16954_/Y vssd1 vssd1 vccd1 vccd1 _17172_/A
+ sky130_fd_sc_hd__a31oi_1
X_14249_ _14433_/D _14797_/B _14003_/A _14002_/A vssd1 vssd1 vccd1 vccd1 _14253_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17394__A2_N _17305_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23556__CLK _23558_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _11840_/X _18813_/A _19156_/B vssd1 vssd1 vccd1 vccd1 _18989_/B sky130_fd_sc_hd__o21ai_1
XFILLER_86_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater101 _23500_/Q vssd1 vssd1 vccd1 vccd1 _14246_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_79_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater112 _23300_/CLK vssd1 vssd1 vccd1 vccd1 _23389_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__19034__A1 _12243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater123 _23349_/CLK vssd1 vssd1 vccd1 vccd1 _23381_/CLK sky130_fd_sc_hd__clkbuf_1
X_17939_ _17936_/X _17938_/Y _23529_/Q vssd1 vssd1 vccd1 vccd1 _18149_/D sky130_fd_sc_hd__o21bai_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13308__B _13377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater134 _23358_/CLK vssd1 vssd1 vccd1 vccd1 _23359_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater145 _23372_/CLK vssd1 vssd1 vccd1 vccd1 _23377_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17045__B1 _19381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater156 _23321_/CLK vssd1 vssd1 vccd1 vccd1 _23327_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_27_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20950_ _20950_/A _20950_/B _20950_/C vssd1 vssd1 vccd1 vccd1 _20984_/C sky130_fd_sc_hd__nand3_2
XFILLER_27_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19609_ _19609_/A _19609_/B vssd1 vssd1 vccd1 vccd1 _19609_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20881_ _21031_/A _21030_/B _20880_/A vssd1 vssd1 vccd1 vccd1 _20882_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11880__A2 _11801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22620_ _22629_/A _22629_/B _22629_/C _22529_/A vssd1 vssd1 vccd1 vccd1 _22623_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_59_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12290__C1 _12289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22551_ _22473_/B _22473_/A _22500_/C vssd1 vssd1 vccd1 vccd1 _22551_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_195_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19011__A _19011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21502_ _21502_/A _21502_/B _21502_/C _21502_/D vssd1 vssd1 vccd1 vccd1 _21504_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_22_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22482_ _22478_/X _22480_/Y _22489_/A vssd1 vssd1 vccd1 vccd1 _22493_/A sky130_fd_sc_hd__o21bai_1
XFILLER_10_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18848__A1 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21433_ _21433_/A _21433_/B vssd1 vssd1 vccd1 vccd1 _21433_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14582__A1 _11665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18848__B2 _11936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21301__C1 _21061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14582__B2 _15664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18850__A _19123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16859__B1 _16592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21364_ _21285_/C _21453_/B _21453_/C vssd1 vssd1 vccd1 vccd1 _21377_/B sky130_fd_sc_hd__nand3b_2
XFILLER_135_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20315_ _20366_/A _20314_/X _20265_/B _20366_/C _20274_/B vssd1 vssd1 vccd1 vccd1
+ _20331_/A sky130_fd_sc_hd__o41a_2
X_23103_ _23103_/A vssd1 vssd1 vccd1 vccd1 _23377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21295_ _21438_/A _21295_/B _21358_/C _21299_/A vssd1 vssd1 vccd1 vccd1 _21295_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_190_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19384__C _19569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16370__A _16370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20246_ _20246_/A vssd1 vssd1 vccd1 vccd1 _20252_/A sky130_fd_sc_hd__inv_2
XFILLER_116_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23034_ _23347_/Q input28/X _23034_/S vssd1 vssd1 vccd1 vccd1 _23035_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18076__A2 _17406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16087__A1 _16167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20958__A2 _12862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16087__B2 _15890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20177_ _20177_/A _20177_/B vssd1 vssd1 vccd1 vccd1 _20177_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_98 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14098__B1 _14097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15295__C1 _15353_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19025__A1 _17627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21907__A1 _22045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15714__A _16856_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _11947_/A _18434_/B _11947_/C vssd1 vssd1 vccd1 vccd1 _11951_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__11856__C1 _18481_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11961__B _23256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ _11788_/A _16462_/B _18952_/D _11803_/X _11880_/X vssd1 vssd1 vccd1 vccd1
+ _11881_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19328__A2 _12103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13620_ _13620_/A _13620_/B _13620_/C vssd1 vssd1 vccd1 vccd1 _13620_/X sky130_fd_sc_hd__or3_2
XFILLER_72_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22818_ _22818_/A _22818_/B _22818_/C _22821_/A vssd1 vssd1 vccd1 vccd1 _22818_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_60_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18536__B1 _12222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13551_ _13537_/A _13536_/B _13536_/C vssd1 vssd1 vccd1 vccd1 _13755_/B sky130_fd_sc_hd__a21o_1
XFILLER_186_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16547__C1 _16066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22749_ _22749_/A _22749_/B _22749_/C vssd1 vssd1 vccd1 vccd1 _22813_/B sky130_fd_sc_hd__nand3_1
XFILLER_186_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12502_ _17964_/C _17964_/A _15957_/C _16795_/C vssd1 vssd1 vccd1 vccd1 _12506_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_186_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16270_ _16586_/A _16586_/B _16270_/C vssd1 vssd1 vccd1 vccd1 _16585_/A sky130_fd_sc_hd__nand3_1
XFILLER_125_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13482_ _13482_/A _13482_/B vssd1 vssd1 vccd1 vccd1 _13482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15221_ _15221_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15221_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12433_ _18435_/A _12099_/D _12100_/B _12121_/A vssd1 vssd1 vccd1 vccd1 _12435_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19500__A2 _16523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15152_ _14184_/A _14184_/B _13960_/Y _14115_/Y vssd1 vssd1 vccd1 vccd1 _15267_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__20217__D _20217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ _12364_/A _12364_/B _12364_/C vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__nand3_1
XFILLER_193_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15117__A3 _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ _14090_/X _14098_/X _14164_/B vssd1 vssd1 vccd1 vccd1 _14139_/B sky130_fd_sc_hd__o21ai_1
XFILLER_154_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22713__C _22713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19960_ _19960_/A _20072_/C vssd1 vssd1 vccd1 vccd1 _19960_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15083_ _15356_/A _14243_/A _14901_/X _15082_/B _15017_/D vssd1 vssd1 vccd1 vccd1
+ _15083_/X sky130_fd_sc_hd__a32o_1
X_12295_ _12295_/A vssd1 vssd1 vccd1 vccd1 _12339_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23579__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23528__D _23528_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18911_ _12563_/A _12563_/B _12563_/C _19089_/B vssd1 vssd1 vccd1 vccd1 _18911_/X
+ sky130_fd_sc_hd__o31a_1
X_14034_ _23498_/Q vssd1 vssd1 vccd1 vccd1 _14261_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17095__B _17095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19891_ _19725_/C _19725_/A _19725_/B _19730_/B vssd1 vssd1 vccd1 vccd1 _19897_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18842_ _18803_/A _18844_/D _18841_/Y vssd1 vssd1 vccd1 vccd1 _18845_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12313__A _19653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14628__A2 _18799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18773_ _18773_/A _18773_/B _18773_/C _18773_/D vssd1 vssd1 vccd1 vccd1 _18774_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_121_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15985_ _15985_/A _15985_/B _15985_/C vssd1 vssd1 vccd1 vccd1 _15986_/A sky130_fd_sc_hd__nand3_1
X_17724_ _17724_/A _17724_/B vssd1 vssd1 vccd1 vccd1 _17724_/Y sky130_fd_sc_hd__nand2_1
X_14936_ _15044_/C _14936_/B vssd1 vssd1 vccd1 vccd1 _14938_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18000__A _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17655_ _17654_/Y _17481_/D _17481_/C vssd1 vssd1 vccd1 vccd1 _17658_/A sky130_fd_sc_hd__a21boi_1
X_14867_ _15094_/A _15094_/B _14867_/C vssd1 vssd1 vccd1 vccd1 _14904_/A sky130_fd_sc_hd__nand3_1
XFILLER_91_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19319__A2 _19172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16606_ _16604_/X _16311_/X _16128_/X _16124_/X _16605_/X vssd1 vssd1 vccd1 vccd1
+ _16647_/B sky130_fd_sc_hd__o32a_1
X_13818_ _13818_/A _13818_/B _21925_/B _21877_/A vssd1 vssd1 vccd1 vccd1 _13819_/B
+ sky130_fd_sc_hd__and4_1
X_17586_ _17586_/A vssd1 vssd1 vccd1 vccd1 _20138_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14798_ _14798_/A _14798_/B vssd1 vssd1 vccd1 vccd1 _14798_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18527__B1 _18526_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19325_ _19325_/A _19325_/B _19477_/A _19477_/B vssd1 vssd1 vccd1 vccd1 _19325_/Y
+ sky130_fd_sc_hd__nand4_2
X_16537_ _16749_/C _17445_/A _16445_/A _16536_/X vssd1 vssd1 vccd1 vccd1 _16564_/B
+ sky130_fd_sc_hd__a31oi_2
X_13749_ _13745_/Y _13747_/X _13748_/Y _13738_/X vssd1 vssd1 vccd1 vccd1 _13749_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19256_ _19256_/A _19256_/B _19256_/C vssd1 vssd1 vccd1 vccd1 _19256_/X sky130_fd_sc_hd__and3_1
X_16468_ _16539_/A _16539_/C _16539_/B vssd1 vssd1 vccd1 vccd1 _16518_/C sky130_fd_sc_hd__a21boi_2
XFILLER_177_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18207_ _18207_/A vssd1 vssd1 vccd1 vccd1 _18207_/X sky130_fd_sc_hd__clkbuf_2
X_15419_ _15419_/A _15419_/B _15419_/C _15419_/D vssd1 vssd1 vccd1 vccd1 _15420_/D
+ sky130_fd_sc_hd__nand4_2
XANTENNA__14564__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19187_ _19047_/B _19047_/A _19185_/X _19186_/Y vssd1 vssd1 vccd1 vccd1 _19188_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__19155__A_N _18799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16399_ _16399_/A vssd1 vssd1 vccd1 vccd1 _16399_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_980 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18138_ _18138_/A _18138_/B vssd1 vssd1 vccd1 vccd1 _18139_/D sky130_fd_sc_hd__nand2_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19485__B _19700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18069_ _17928_/A _17928_/B _17836_/Y _18129_/B vssd1 vssd1 vccd1 vccd1 _18069_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_144_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20100_ _20103_/C _20177_/B vssd1 vssd1 vccd1 vccd1 _20102_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21080_ _21430_/C _21196_/A _20953_/X _20963_/Y _20967_/B vssd1 vssd1 vccd1 vccd1
+ _21082_/C sky130_fd_sc_hd__a32o_1
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22920__A _22966_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16069__A1 _17248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20031_ _20031_/A vssd1 vssd1 vccd1 vccd1 _20031_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__21062__A1 _20639_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20404__A4 _20368_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15260__A1_N _14212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21982_ _21982_/A _21982_/B vssd1 vssd1 vccd1 vccd1 _22089_/B sky130_fd_sc_hd__nand2_2
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18766__B1 _12353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15253__B _15253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20933_ _20919_/Y _20929_/Y _20940_/B vssd1 vssd1 vccd1 vccd1 _20937_/B sky130_fd_sc_hd__o21ai_1
XFILLER_81_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20864_ _20851_/Y _20857_/Y _20859_/Y _20863_/Y vssd1 vssd1 vccd1 vccd1 _21157_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__21271__A _21387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22603_ _22601_/Y _22756_/C _13816_/A _22602_/Y vssd1 vssd1 vccd1 vccd1 _22633_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23583_ _23588_/CLK _23583_/D vssd1 vssd1 vccd1 vccd1 _23583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16365__A _16365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20795_ _23299_/Q vssd1 vssd1 vccd1 vccd1 _21047_/C sky130_fd_sc_hd__clkinv_2
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22534_ _22530_/Y _22532_/Y _22533_/X vssd1 vssd1 vccd1 vccd1 _22536_/A sky130_fd_sc_hd__o21a_1
XFILLER_195_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_bq_clk_i clkbuf_4_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _23559_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14555__A1 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19479__D1 _18479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14555__B2 _13226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22465_ _22700_/A _22554_/A _22553_/D _22465_/D vssd1 vssd1 vccd1 vccd1 _22465_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_183_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_618 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21416_ _21616_/A _21617_/A _21346_/X _21340_/Y _21411_/Y vssd1 vssd1 vccd1 vccd1
+ _21418_/B sky130_fd_sc_hd__o221ai_2
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1044 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22396_ _22289_/B _22289_/Y _22395_/Y vssd1 vssd1 vccd1 vccd1 _22412_/A sky130_fd_sc_hd__a21o_1
XFILLER_191_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12117__B _19709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21347_ _21342_/Y _21343_/Y _21346_/X _21247_/X vssd1 vssd1 vccd1 vccd1 _21347_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20334__B _20363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12080_ _18778_/C _12080_/B _18163_/A vssd1 vssd1 vccd1 vccd1 _12231_/A sky130_fd_sc_hd__and3_1
XFILLER_150_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21278_ _21278_/A _21448_/B _21502_/A vssd1 vssd1 vccd1 vccd1 _21278_/X sky130_fd_sc_hd__and3_1
X_23017_ _23339_/Q input20/X _23023_/S vssd1 vssd1 vccd1 vccd1 _23018_/A sky130_fd_sc_hd__mux2_1
X_20229_ _20229_/A _20229_/B _20229_/C vssd1 vssd1 vccd1 vccd1 _20231_/B sky130_fd_sc_hd__and3_1
XFILLER_89_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15770_ _12207_/A _15883_/A _15843_/A _15852_/A _15754_/A vssd1 vssd1 vccd1 vccd1
+ _15770_/X sky130_fd_sc_hd__o221a_1
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12982_ _12981_/X _12955_/Y _12972_/A vssd1 vssd1 vccd1 vccd1 _12984_/A sky130_fd_sc_hd__o21ai_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _14729_/A vssd1 vssd1 vccd1 vccd1 _18435_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_input12_A wb_dat_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _18859_/A _18859_/D _12260_/C _18531_/A vssd1 vssd1 vccd1 vccd1 _11966_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18755__A _18755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _17440_/A vssd1 vssd1 vccd1 vccd1 _17580_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_62 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _15114_/B vssd1 vssd1 vccd1 vccd1 _15338_/A sky130_fd_sc_hd__buf_4
XFILLER_73_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11864_ _11896_/A vssd1 vssd1 vccd1 vccd1 _11864_/X sky130_fd_sc_hd__buf_4
XANTENNA__21108__A2 _21109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22277__A _22364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _23327_/Q vssd1 vssd1 vccd1 vccd1 _13603_/X sky130_fd_sc_hd__clkbuf_4
X_17371_ _17522_/B _17522_/C _17522_/D _17832_/A vssd1 vssd1 vccd1 vccd1 _17372_/B
+ sky130_fd_sc_hd__a31oi_2
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ input49/X _14549_/A _14545_/A _14031_/X _14582_/X vssd1 vssd1 vccd1 vccd1
+ _14583_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16275__A _16275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11795_ _12145_/B _19157_/C _12145_/A vssd1 vssd1 vccd1 vccd1 _12016_/A sky130_fd_sc_hd__nand3_4
XFILLER_159_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19110_ _19075_/C _19075_/B _19075_/A _19087_/A _19082_/X vssd1 vssd1 vccd1 vccd1
+ _19275_/A sky130_fd_sc_hd__a32o_1
X_16322_ _16389_/A _16322_/B vssd1 vssd1 vccd1 vccd1 _16322_/X sky130_fd_sc_hd__or2_1
XANTENNA__20509__B _20509_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13534_ _13544_/A _13544_/B _13545_/A vssd1 vssd1 vccd1 vccd1 _13535_/B sky130_fd_sc_hd__a21oi_1
XFILLER_186_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19041_ _19040_/X _20081_/B _19031_/X _18958_/C _19033_/A vssd1 vssd1 vccd1 vccd1
+ _19041_/X sky130_fd_sc_hd__o311a_1
XFILLER_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16253_ _16253_/A _16253_/B vssd1 vssd1 vccd1 vccd1 _16254_/D sky130_fd_sc_hd__nand2_1
X_13465_ _13465_/A vssd1 vssd1 vccd1 vccd1 _13465_/X sky130_fd_sc_hd__buf_2
XANTENNA__15743__B1 _15662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18490__A _18490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12308__A _12308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15204_ _15132_/A _15132_/B _15132_/C vssd1 vssd1 vccd1 vccd1 _15204_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21816__B1 _22420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12416_ _12410_/Y _18653_/C _18997_/A vssd1 vssd1 vccd1 vccd1 _18788_/A sky130_fd_sc_hd__a21o_2
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16184_ _15932_/A _15933_/Y _15937_/A vssd1 vssd1 vccd1 vccd1 _16194_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__12021__A2 _12020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13396_ _13620_/B vssd1 vssd1 vccd1 vccd1 _22420_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15135_ _15134_/C _15134_/B _15080_/X vssd1 vssd1 vccd1 vccd1 _15136_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__21292__A1 _20502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ _17546_/C _19903_/C _19261_/C _16528_/B vssd1 vssd1 vccd1 vccd1 _12348_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__15619__A _23429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14523__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output80_A _14572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19943_ _19943_/A _19943_/B vssd1 vssd1 vccd1 vccd1 _19943_/Y sky130_fd_sc_hd__nand2_1
X_15066_ _15067_/A _15064_/X _15065_/Y _14959_/C vssd1 vssd1 vccd1 vccd1 _15066_/Y
+ sky130_fd_sc_hd__a22oi_4
X_12278_ _16437_/A vssd1 vssd1 vccd1 vccd1 _12279_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_142_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14242__B _15082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14017_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14017_/X sky130_fd_sc_hd__buf_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21044__B2 _21635_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19874_ _19874_/A _19874_/B _20003_/A _19888_/D vssd1 vssd1 vccd1 vccd1 _19879_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12043__A _19323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18825_ _18825_/A _18825_/B vssd1 vssd1 vccd1 vccd1 _18844_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17263__A3 _16056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18756_ _18756_/A _18756_/B _19364_/B vssd1 vssd1 vccd1 vccd1 _18932_/B sky130_fd_sc_hd__nand3_4
XFILLER_49_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13285__A1 _13465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15968_ _15968_/A vssd1 vssd1 vccd1 vccd1 _17041_/B sky130_fd_sc_hd__buf_2
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17707_ _17426_/A _17557_/Y _17487_/B _17553_/Y vssd1 vssd1 vccd1 vccd1 _17810_/B
+ sky130_fd_sc_hd__o211ai_2
X_14919_ _14923_/C vssd1 vssd1 vccd1 vccd1 _14926_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18687_ _18687_/A _18687_/B _18687_/C vssd1 vssd1 vccd1 vccd1 _18784_/B sky130_fd_sc_hd__nand3_2
X_15899_ _15899_/A vssd1 vssd1 vccd1 vccd1 _15899_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17638_ _17454_/Y _17467_/X _17460_/B _17457_/Y vssd1 vssd1 vccd1 vccd1 _17641_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17569_ _17569_/A vssd1 vssd1 vccd1 vccd1 _20317_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_143_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19173__B1 _19670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19308_ _19652_/A _19308_/B _19308_/C vssd1 vssd1 vccd1 vccd1 _19309_/B sky130_fd_sc_hd__nand3_1
XFILLER_177_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20580_ _20578_/X _20736_/B _20576_/Y _20568_/Y vssd1 vssd1 vccd1 vccd1 _20580_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20138__C _20320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19239_ _19217_/X _19222_/X _19189_/X _19228_/X vssd1 vssd1 vccd1 vccd1 _19239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22250_ _21850_/A _21850_/B _22247_/Y _22445_/B vssd1 vssd1 vccd1 vccd1 _22252_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17728__B _17885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21201_ _21191_/Y _21192_/Y _21431_/C _21196_/A _21194_/Y vssd1 vssd1 vccd1 vccd1
+ _21307_/B sky130_fd_sc_hd__o2111ai_4
XANTENNA__21283__A1 _21440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22181_ _22028_/A _21853_/A _22141_/C vssd1 vssd1 vccd1 vccd1 _22560_/B sky130_fd_sc_hd__a21o_2
XANTENNA__21283__B2 _21276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_994 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21132_ _21132_/A _21132_/B vssd1 vssd1 vccd1 vccd1 _21132_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16070__D _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21063_ _12815_/B _21061_/X _20960_/Y vssd1 vssd1 vccd1 vccd1 _21063_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_48_16 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19662__C _19662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20014_ _19040_/X _18373_/A _20013_/Y _20013_/A vssd1 vssd1 vccd1 vccd1 _20108_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_154_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input4_A wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23184__C input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19381__D _19381_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11792__A _11792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23274__CLK _23492_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21965_ _21965_/A _21965_/B _21965_/C vssd1 vssd1 vccd1 vccd1 _21981_/B sky130_fd_sc_hd__nand3_4
XFILLER_55_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16214__A1 _12018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17411__B1 _17410_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _20916_/A vssd1 vssd1 vccd1 vccd1 _21358_/A sky130_fd_sc_hd__buf_2
XANTENNA__17962__A1 _18211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21896_ _21896_/A vssd1 vssd1 vccd1 vccd1 _22045_/A sky130_fd_sc_hd__buf_2
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14776__A1 _14245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ _20847_/A _20847_/B vssd1 vssd1 vccd1 vccd1 _20849_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_744 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23566_ _23566_/CLK _23566_/D vssd1 vssd1 vccd1 vccd1 _23566_/Q sky130_fd_sc_hd__dfxtp_1
X_11580_ _23589_/Q vssd1 vssd1 vccd1 vccd1 _11593_/C sky130_fd_sc_hd__clkinv_2
XFILLER_11_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20778_ _20778_/A vssd1 vssd1 vccd1 vccd1 _20778_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14528__A1 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22517_ _22405_/A _22418_/X _22420_/X vssd1 vssd1 vccd1 vccd1 _22517_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23497_ _23499_/CLK _23497_/D vssd1 vssd1 vccd1 vccd1 _23497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12539__B1 _12227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_747 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13250_ _23321_/Q vssd1 vssd1 vccd1 vccd1 _13253_/A sky130_fd_sc_hd__clkbuf_4
X_22448_ _23276_/Q _22448_/B vssd1 vssd1 vccd1 vccd1 _22450_/A sky130_fd_sc_hd__nand2_1
XFILLER_129_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12201_ _12057_/A _12057_/C _12057_/B vssd1 vssd1 vccd1 vccd1 _12387_/B sky130_fd_sc_hd__a21oi_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13181_ _13181_/A _13181_/B _13181_/C vssd1 vssd1 vccd1 vccd1 _13181_/X sky130_fd_sc_hd__and3_1
X_22379_ _22381_/B vssd1 vssd1 vccd1 vccd1 _22637_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_191_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19219__A1 _19218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ _18445_/B vssd1 vssd1 vccd1 vccd1 _19308_/B sky130_fd_sc_hd__buf_4
XFILLER_135_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22560__A _22560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16940_ _16939_/Y _16708_/A _16706_/A vssd1 vssd1 vccd1 vccd1 _16948_/A sky130_fd_sc_hd__o21ai_2
X_12063_ _12254_/A _12392_/C _12253_/A vssd1 vssd1 vccd1 vccd1 _12388_/B sky130_fd_sc_hd__a21boi_1
XFILLER_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20080__A _20080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16871_ _16604_/A _16315_/A _16058_/A _11926_/A vssd1 vssd1 vccd1 vccd1 _16871_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12798__A _23455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16453__A1 _16370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15256__A2 _15353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18610_ _18620_/A vssd1 vssd1 vccd1 vccd1 _18931_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12013__D _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16453__B2 _16225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15822_ _11882_/X _11883_/X _15716_/B _15712_/D vssd1 vssd1 vccd1 vccd1 _15822_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19590_ _19475_/X _19527_/Y _19583_/Y vssd1 vssd1 vccd1 vccd1 _19590_/Y sky130_fd_sc_hd__o21ai_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18541_ _18541_/A vssd1 vssd1 vccd1 vccd1 _18721_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15753_ _15753_/A _15753_/B vssd1 vssd1 vccd1 vccd1 _15754_/A sky130_fd_sc_hd__nand2_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _21193_/C vssd1 vssd1 vccd1 vccd1 _21358_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_94 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ _11916_/A vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__buf_2
XFILLER_18_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14704_ _23376_/Q _14688_/X _14703_/X vssd1 vssd1 vccd1 vccd1 _14704_/X sky130_fd_sc_hd__o21a_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ _11848_/X _12053_/A _12241_/A _18490_/A vssd1 vssd1 vccd1 vccd1 _18473_/A
+ sky130_fd_sc_hd__o22ai_2
X_15684_ _15712_/A vssd1 vssd1 vccd1 vccd1 _15686_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _12896_/A _12896_/B _12896_/C vssd1 vssd1 vccd1 vccd1 _12902_/C sky130_fd_sc_hd__nand3_2
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_536 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _17625_/B vssd1 vssd1 vccd1 vccd1 _17959_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14635_/A vssd1 vssd1 vccd1 vccd1 _14635_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11847_ _11847_/A vssd1 vssd1 vccd1 vccd1 _18500_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13422__A _13453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17354_ _16952_/Y _17191_/Y _17198_/Y _17189_/Y vssd1 vssd1 vccd1 vccd1 _17354_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_14566_ _13253_/A _14532_/X _14534_/X _14565_/X vssd1 vssd1 vccd1 vccd1 _14566_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11860_/A _11860_/B _11860_/C vssd1 vssd1 vccd1 vccd1 _11883_/A sky130_fd_sc_hd__nand3_1
XANTENNA__21501__A2 _21548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16305_ _16302_/Y _16303_/Y _16304_/Y vssd1 vssd1 vccd1 vccd1 _16306_/A sky130_fd_sc_hd__o21ai_1
X_13517_ _13517_/A _13517_/B _13517_/C vssd1 vssd1 vccd1 vccd1 _13519_/B sky130_fd_sc_hd__nand3_1
X_17285_ _17285_/A vssd1 vssd1 vccd1 vccd1 _17285_/X sky130_fd_sc_hd__buf_2
XFILLER_159_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14497_ _14497_/A _14497_/B _14497_/C vssd1 vssd1 vccd1 vccd1 _14498_/B sky130_fd_sc_hd__nand3_1
X_19024_ _19029_/A _19029_/D vssd1 vssd1 vccd1 vccd1 _19026_/B sky130_fd_sc_hd__nand2_1
X_16236_ _16236_/A _16236_/B _16236_/C vssd1 vssd1 vccd1 vccd1 _16236_/X sky130_fd_sc_hd__and3_1
XFILLER_173_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13448_ _13448_/A vssd1 vssd1 vccd1 vccd1 _13517_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16167_ _16641_/A _16641_/B _16167_/C _20062_/C vssd1 vssd1 vccd1 vccd1 _16650_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_142_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13379_ _23324_/Q vssd1 vssd1 vccd1 vccd1 _13379_/X sky130_fd_sc_hd__buf_2
XFILLER_170_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15118_ _15118_/A _15257_/B _15233_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15120_/D
+ sky130_fd_sc_hd__nand4_4
XANTENNA__12950__B1 _12674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16098_ _16093_/Y _16096_/Y _16072_/Y _16097_/Y vssd1 vssd1 vccd1 vccd1 _16424_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16692__A1 _16054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19926_ _19427_/X _19433_/Y _19439_/Y vssd1 vssd1 vccd1 vccd1 _19926_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15049_ _15049_/A _15049_/B _15049_/C vssd1 vssd1 vccd1 vccd1 _15053_/A sky130_fd_sc_hd__nand3_1
XANTENNA__16692__B2 _16684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20702__B _23456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19857_ _12279_/X _20263_/A _19853_/Y _19856_/Y vssd1 vssd1 vccd1 vccd1 _19873_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13019__D _20798_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16444__B2 _16479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18808_ _18808_/A _18808_/B _18808_/C vssd1 vssd1 vccd1 vccd1 _18844_/D sky130_fd_sc_hd__nand3_2
X_19788_ _19788_/A _19923_/A _19788_/C vssd1 vssd1 vccd1 vccd1 _19788_/Y sky130_fd_sc_hd__nand3_1
XFILLER_23_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21814__A _21987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18739_ _23540_/Q vssd1 vssd1 vccd1 vccd1 _18739_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16908__A _16908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21750_ _21747_/Y _21749_/Y _13791_/A vssd1 vssd1 vccd1 vccd1 _21750_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20701_ _20542_/A _20542_/B _20542_/C _20553_/C vssd1 vssd1 vccd1 vccd1 _20701_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21681_ _21691_/A _21691_/B _21691_/C vssd1 vssd1 vccd1 vccd1 _21688_/C sky130_fd_sc_hd__nand3_1
XFILLER_145_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23420_ _23424_/CLK _23420_/D vssd1 vssd1 vccd1 vccd1 _23420_/Q sky130_fd_sc_hd__dfxtp_1
X_20632_ _20632_/A _20632_/B vssd1 vssd1 vccd1 vccd1 _20635_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19697__A1 _19903_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23351_ _23352_/CLK _23351_/D vssd1 vssd1 vccd1 vccd1 _23351_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13051__B _23455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20563_ _20563_/A _20563_/B _23457_/Q vssd1 vssd1 vccd1 vccd1 _20566_/B sky130_fd_sc_hd__and3_1
XFILLER_149_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22364__B _22364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22302_ _22476_/A _22476_/B _22392_/C vssd1 vssd1 vccd1 vccd1 _22302_/X sky130_fd_sc_hd__and3_1
XFILLER_165_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15183__A1 _14212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23282_ _23510_/CLK _23282_/D vssd1 vssd1 vccd1 vccd1 _23282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20494_ _20798_/A _20897_/C _20798_/C _20494_/D vssd1 vssd1 vccd1 vccd1 _20495_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12890__B _13052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20059__A2 _18211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22233_ _22225_/A _22231_/B _22232_/X vssd1 vssd1 vccd1 vccd1 _22234_/C sky130_fd_sc_hd__a21o_1
XFILLER_173_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22164_ _22164_/A vssd1 vssd1 vccd1 vccd1 _22754_/B sky130_fd_sc_hd__buf_2
XFILLER_59_26 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21115_ _21115_/A _21115_/B vssd1 vssd1 vccd1 vccd1 _21159_/B sky130_fd_sc_hd__xor2_1
XFILLER_120_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22095_ _22754_/A vssd1 vssd1 vccd1 vccd1 _22830_/B sky130_fd_sc_hd__buf_2
XFILLER_8_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19621__A1 _18673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21046_ _21046_/A _21046_/B _23299_/Q vssd1 vssd1 vccd1 vccd1 _21048_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19621__B2 _12353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11901__D1 _16497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17093__D1 _16866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1078 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22997_ _21902_/B input10/X _23001_/S vssd1 vssd1 vccd1 vccd1 _22998_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _12997_/C vssd1 vssd1 vccd1 vccd1 _20473_/C sky130_fd_sc_hd__clkbuf_2
X_21948_ _21943_/X _21944_/X _21936_/Y _21941_/Y vssd1 vssd1 vccd1 vccd1 _21948_/Y
+ sky130_fd_sc_hd__o211ai_2
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11682_/Y _18859_/B _16674_/A vssd1 vssd1 vccd1 vccd1 _11717_/B sky130_fd_sc_hd__nand3b_4
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _23447_/Q vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__clkbuf_4
X_21879_ _21762_/Y _22126_/A _21783_/A vssd1 vssd1 vccd1 vccd1 _21984_/B sky130_fd_sc_hd__o21ai_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14420_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14422_/A sky130_fd_sc_hd__inv_2
XANTENNA__13242__A _23477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11632_ _23598_/Q vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__clkinv_4
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12224__A2 _12223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14351_ _14324_/A _14319_/Y _14318_/Y _14344_/B vssd1 vssd1 vccd1 vccd1 _14352_/B
+ sky130_fd_sc_hd__o211a_1
X_23549_ _23578_/CLK _23549_/D vssd1 vssd1 vccd1 vccd1 _23549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _13303_/A _13303_/C _13303_/B vssd1 vssd1 vccd1 vccd1 _13538_/A sky130_fd_sc_hd__o21a_1
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17070_ _17070_/A vssd1 vssd1 vccd1 vccd1 _17070_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15174__A1 _14181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14282_ _14361_/C _14361_/A _14282_/C vssd1 vssd1 vccd1 vccd1 _14349_/D sky130_fd_sc_hd__nand3_1
XFILLER_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16910__A2 _16908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16021_ _16073_/A _16073_/B _16020_/X vssd1 vssd1 vccd1 vccd1 _16021_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_183_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13233_ _23320_/Q vssd1 vssd1 vccd1 vccd1 _13233_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22995__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164_ _21172_/A vssd1 vssd1 vccd1 vccd1 _21440_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__19860__A1 _20081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12115_ _12114_/Y _11665_/Y _12118_/C vssd1 vssd1 vccd1 vccd1 _19364_/A sky130_fd_sc_hd__a21boi_4
XANTENNA__21379__A2_N _21376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17972_ _17972_/A vssd1 vssd1 vccd1 vccd1 _19113_/C sky130_fd_sc_hd__clkbuf_2
X_13095_ _21490_/B vssd1 vssd1 vccd1 vccd1 _21455_/B sky130_fd_sc_hd__buf_2
XANTENNA__23536__D _23536_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19711_ _12053_/X _17763_/A _19819_/A _19820_/A vssd1 vssd1 vccd1 vccd1 _19713_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12024__C _15718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16923_ _16923_/A _16923_/B _16923_/C vssd1 vssd1 vccd1 vccd1 _16923_/X sky130_fd_sc_hd__and3_1
X_12046_ _12046_/A _12046_/B vssd1 vssd1 vccd1 vccd1 _12049_/A sky130_fd_sc_hd__nand2_1
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19642_ _19475_/X _19527_/Y _19641_/Y vssd1 vssd1 vccd1 vccd1 _19733_/A sky130_fd_sc_hd__o21ai_1
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16854_ _16153_/B _16617_/X _16635_/B _16614_/Y vssd1 vssd1 vccd1 vccd1 _16879_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_37_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15805_ _16677_/C vssd1 vssd1 vccd1 vccd1 _16213_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19573_ _19573_/A _19573_/B _19573_/C vssd1 vssd1 vccd1 vccd1 _19573_/X sky130_fd_sc_hd__and3_1
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13997_ _13933_/A _13933_/B _13953_/Y _13996_/Y vssd1 vssd1 vccd1 vccd1 _13997_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16785_ _16744_/A _16744_/B _16784_/Y vssd1 vssd1 vccd1 vccd1 _16787_/B sky130_fd_sc_hd__a21o_1
XANTENNA__23172__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18524_ _18524_/A _18524_/B vssd1 vssd1 vccd1 vccd1 _18524_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15632__A _23429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15736_ _15736_/A vssd1 vssd1 vccd1 vccd1 _15862_/A sky130_fd_sc_hd__clkbuf_4
X_12948_ _13176_/A _21054_/C _13176_/C vssd1 vssd1 vccd1 vccd1 _12981_/B sky130_fd_sc_hd__and3_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23271__D _23271_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16729__A2 _16723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16447__B _16447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18455_ _18455_/A _18460_/A vssd1 vssd1 vccd1 vccd1 _19969_/A sky130_fd_sc_hd__nor2_4
XFILLER_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _12894_/B vssd1 vssd1 vccd1 vccd1 _12899_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15667_ _15920_/A _15920_/B _16667_/B _15918_/C vssd1 vssd1 vccd1 vccd1 _15668_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17406_ _17406_/A _17406_/B _17753_/A _17753_/B vssd1 vssd1 vccd1 vccd1 _17406_/Y
+ sky130_fd_sc_hd__nand4_4
X_14618_ _14614_/X _14550_/A _14526_/X _14615_/X _14617_/X vssd1 vssd1 vccd1 vccd1
+ _14618_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18386_ _18288_/A _18288_/B _18288_/C _18384_/A _18388_/B vssd1 vssd1 vccd1 vccd1
+ _18411_/B sky130_fd_sc_hd__a2111oi_1
XFILLER_18_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15598_ _15628_/A _15685_/A _15614_/A vssd1 vssd1 vccd1 vccd1 _15715_/A sky130_fd_sc_hd__nand3_2
XANTENNA__17139__C1 _15937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_90 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17337_ _17337_/A _17337_/B _17337_/C vssd1 vssd1 vccd1 vccd1 _17341_/A sky130_fd_sc_hd__nand3_1
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14549_ _14549_/A vssd1 vssd1 vccd1 vccd1 _14549_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17154__A2 _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11974__B2 _11942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17268_ _17275_/A _17275_/B _17268_/C vssd1 vssd1 vccd1 vccd1 _17268_/Y sky130_fd_sc_hd__nand3_1
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19007_ _19007_/A _19007_/B vssd1 vssd1 vccd1 vccd1 _19007_/Y sky130_fd_sc_hd__nand2_1
X_16219_ _16183_/X _16193_/Y _16199_/Y _16233_/B _16710_/A vssd1 vssd1 vccd1 vccd1
+ _16219_/Y sky130_fd_sc_hd__o2111ai_4
X_17199_ _16955_/X _17185_/Y _17198_/Y _17189_/Y vssd1 vssd1 vccd1 vccd1 _17200_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__22986__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17311__C1 _17307_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15807__A _15807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19909_ _19909_/A _19909_/B _19909_/C vssd1 vssd1 vccd1 vccd1 _19928_/D sky130_fd_sc_hd__nand3_1
XFILLER_69_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14430__B _15094_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20151__C _20151_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20213__A2 _19700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17614__B1 _17606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22920_ _22966_/S vssd1 vssd1 vccd1 vccd1 _22929_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_84_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14428__B1 _14181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16968__A2 _18277_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22851_ _22845_/Y _22848_/Y _23283_/Q vssd1 vssd1 vccd1 vccd1 _22851_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__23163__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21802_ _21801_/B _21801_/C _21801_/A vssd1 vssd1 vccd1 vccd1 _21804_/B sky130_fd_sc_hd__a21oi_1
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15640__A2 _11865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22782_ _22783_/B _23281_/Q vssd1 vssd1 vccd1 vccd1 _22784_/A sky130_fd_sc_hd__and2_1
XANTENNA__12454__A2 _19530_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22910__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21733_ _13615_/A _21916_/A _13797_/B _13793_/Y vssd1 vssd1 vccd1 vccd1 _21754_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__11662__B1 _11665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19949__A _19949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19119__B1 _12283_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18853__A _18959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21664_ _21630_/A _21666_/B _21614_/Y vssd1 vssd1 vccd1 vccd1 _21665_/B sky130_fd_sc_hd__a21oi_1
XFILLER_12_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23403_ _23434_/CLK _23403_/D vssd1 vssd1 vccd1 vccd1 _23403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20615_ _12987_/Y _20459_/Y _20605_/A vssd1 vssd1 vccd1 vccd1 _20615_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_165_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12757__A3 _20639_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__C1 _12608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21595_ _21633_/A _21595_/B _21595_/C vssd1 vssd1 vccd1 vccd1 _21597_/A sky130_fd_sc_hd__and3_1
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23334_ _23429_/CLK _23334_/D vssd1 vssd1 vccd1 vccd1 _23334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_330 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20546_ _20728_/A _20714_/A _20713_/B vssd1 vssd1 vccd1 vccd1 _20551_/B sky130_fd_sc_hd__nand3_1
XFILLER_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17550__C1 _19862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__23462__CLK _23462_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23265_ _23584_/CLK _23265_/D vssd1 vssd1 vccd1 vccd1 _23265_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20477_ _12632_/A _20471_/Y _20490_/A vssd1 vssd1 vccd1 vccd1 _20484_/B sky130_fd_sc_hd__o21ai_1
XFILLER_193_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22977__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22216_ _22214_/Y _22200_/Y _22215_/X vssd1 vssd1 vccd1 vccd1 _22216_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13182__A3 _20775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19842__A1 _19505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23196_ _23196_/A vssd1 vssd1 vccd1 vccd1 _23418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22147_ _22562_/C vssd1 vssd1 vccd1 vccd1 _22569_/C sky130_fd_sc_hd__buf_2
XANTENNA__15717__A _16856_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22078_ _22069_/Y _22074_/X _22076_/X _22077_/Y vssd1 vssd1 vccd1 vccd1 _22078_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__13237__A _23478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21029_ _21029_/A _21029_/B vssd1 vssd1 vccd1 vccd1 _21029_/X sky130_fd_sc_hd__and2_1
X_13920_ _23356_/Q vssd1 vssd1 vccd1 vccd1 _14077_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_19_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12693__A2 _12850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13851_ _13848_/Y _13849_/Y _13686_/A _21987_/B vssd1 vssd1 vccd1 vccd1 _13857_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19358__B1 _12185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23154__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22269__B _22566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ _13051_/A vssd1 vssd1 vccd1 vccd1 _13176_/A sky130_fd_sc_hd__clkbuf_2
X_16570_ _16570_/A _16570_/B vssd1 vssd1 vccd1 vccd1 _16570_/Y sky130_fd_sc_hd__nand2_1
X_13782_ _23327_/Q vssd1 vssd1 vccd1 vccd1 _13783_/A sky130_fd_sc_hd__inv_2
XANTENNA__22901__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15521_ _15520_/B _15521_/B vssd1 vssd1 vccd1 vccd1 _15522_/B sky130_fd_sc_hd__and2b_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _12733_/A _12733_/B vssd1 vssd1 vccd1 vccd1 _12734_/C sky130_fd_sc_hd__nand2_1
XANTENNA__19859__A _19859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18240_ _18240_/A _18349_/A vssd1 vssd1 vccd1 vccd1 _18245_/C sky130_fd_sc_hd__or2_1
X_15452_ _15371_/B _15451_/B _15446_/A _15451_/D _15451_/C vssd1 vssd1 vccd1 vccd1
+ _15453_/A sky130_fd_sc_hd__a32o_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12664_ _23452_/Q vssd1 vssd1 vccd1 vccd1 _20805_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_31_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14403_/A _14403_/B _14403_/C _14403_/D vssd1 vssd1 vccd1 vccd1 _14405_/B
+ sky130_fd_sc_hd__nand4_1
X_11615_ _23397_/Q vssd1 vssd1 vccd1 vccd1 _11758_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18171_ _17959_/A _18217_/A _17959_/B _18170_/A _18170_/D vssd1 vssd1 vccd1 vccd1
+ _18171_/X sky130_fd_sc_hd__a32o_1
XFILLER_168_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15383_ _15383_/A _15383_/B _15383_/C vssd1 vssd1 vccd1 vccd1 _15383_/X sky130_fd_sc_hd__or3_1
XFILLER_169_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12595_ _23290_/Q vssd1 vssd1 vccd1 vccd1 _12873_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__19297__C _19431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17122_ _17302_/A _17301_/A _17112_/B _17112_/A vssd1 vssd1 vccd1 vccd1 _17124_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_128_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14334_ _14797_/A _14886_/B _14797_/C _14386_/A _14751_/B vssd1 vssd1 vccd1 vccd1
+ _14334_/Y sky130_fd_sc_hd__a32oi_4
XANTENNA__20140__A1 _17600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17098__B _17098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17053_ _16627_/X _17039_/A _16811_/X _16814_/X vssd1 vssd1 vccd1 vccd1 _17053_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_14265_ _14039_/A _14260_/A _14009_/X _15231_/A _14049_/Y vssd1 vssd1 vccd1 vccd1
+ _14290_/B sky130_fd_sc_hd__o221ai_2
XANTENNA__19818__D1 _20146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12316__A _17134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16004_ _15725_/Y _15898_/X _16268_/A _15944_/Y vssd1 vssd1 vccd1 vccd1 _16004_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13216_ _23479_/Q vssd1 vssd1 vccd1 vccd1 _22564_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14196_ _15111_/A _15111_/B _14878_/A _14091_/A vssd1 vssd1 vccd1 vccd1 _14886_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_100_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13147_ _13147_/A _13147_/B _13147_/C vssd1 vssd1 vccd1 vccd1 _13199_/A sky130_fd_sc_hd__nand3_1
XFILLER_97_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18003__A _18003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _17955_/A _17955_/B vssd1 vssd1 vccd1 vccd1 _17956_/A sky130_fd_sc_hd__or2_1
X_13078_ _13078_/A _13078_/B vssd1 vssd1 vccd1 vccd1 _13079_/A sky130_fd_sc_hd__nand2_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18938__A _18938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16906_ _16360_/A _16194_/B _16913_/A vssd1 vssd1 vccd1 vccd1 _16906_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12029_ _12029_/A _12029_/B vssd1 vssd1 vccd1 vccd1 _12159_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12051__A _12051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17886_ _18016_/C _20164_/C _18079_/A _18161_/B _17724_/B vssd1 vssd1 vccd1 vccd1
+ _17886_/X sky130_fd_sc_hd__a41o_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_959 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19625_ _19625_/A _19625_/B _19768_/A _19625_/D vssd1 vssd1 vccd1 vccd1 _19916_/B
+ sky130_fd_sc_hd__nand4_4
X_16837_ _16837_/A _16837_/B _16837_/C vssd1 vssd1 vccd1 vccd1 _16845_/B sky130_fd_sc_hd__and3_1
XFILLER_20_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13618__D1 _13816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19349__B1 _19179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16458__A _16458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23145__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11890__A _19363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19556_ _19040_/X _17976_/A _19358_/Y _19554_/X _19532_/X vssd1 vssd1 vccd1 vccd1
+ _19556_/X sky130_fd_sc_hd__o311a_1
X_16768_ _16768_/A _16768_/B _17010_/A _17009_/A vssd1 vssd1 vccd1 vccd1 _17011_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18507_ _12460_/Y _18503_/Y _18505_/Y _19381_/D _19847_/C vssd1 vssd1 vccd1 vccd1
+ _18510_/C sky130_fd_sc_hd__o2111ai_1
X_15719_ _15719_/A _15719_/B vssd1 vssd1 vccd1 vccd1 _15723_/B sky130_fd_sc_hd__nand2_1
XFILLER_178_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19487_ _18656_/Y _19173_/X _19483_/Y _19486_/Y vssd1 vssd1 vccd1 vccd1 _19577_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__18673__A _18673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16699_ _16699_/A _16699_/B _16699_/C vssd1 vssd1 vccd1 vccd1 _16700_/A sky130_fd_sc_hd__nand3_1
XFILLER_94_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18438_ _18649_/A _19155_/C _18811_/B vssd1 vssd1 vccd1 vccd1 _18439_/A sky130_fd_sc_hd__and3_1
XFILLER_167_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18369_ _18264_/B _18319_/Y _18367_/Y vssd1 vssd1 vccd1 vccd1 _18370_/C sky130_fd_sc_hd__o21a_1
XFILLER_175_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20400_ _20400_/A _20400_/B vssd1 vssd1 vccd1 vccd1 _20401_/C sky130_fd_sc_hd__nand2_1
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15138__A1 _13985_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20131__A1 _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21380_ _21380_/A _21380_/B vssd1 vssd1 vccd1 vccd1 _21380_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19000__C _19308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20331_ _20331_/A _20331_/B vssd1 vssd1 vccd1 vccd1 _20335_/A sky130_fd_sc_hd__xnor2_2
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23050_ _23050_/A vssd1 vssd1 vccd1 vccd1 _23353_/D sky130_fd_sc_hd__clkbuf_1
X_20262_ _19785_/X _20205_/A _20208_/A _20250_/Y vssd1 vssd1 vccd1 vccd1 _20341_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_127_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22001_ _22121_/A _21892_/A _22000_/Y vssd1 vssd1 vccd1 vccd1 _22001_/Y sky130_fd_sc_hd__o21ai_2
X_20193_ _19785_/X _20205_/A _20206_/A _20252_/B vssd1 vssd1 vccd1 vccd1 _20193_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_142_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17455__C _17587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22903_ _12667_/B input29/X _22907_/S vssd1 vssd1 vccd1 vccd1 _22904_/A sky130_fd_sc_hd__mux2_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22089__B _22089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22834_ _22834_/A _22834_/B _22834_/C vssd1 vssd1 vccd1 vccd1 _22836_/A sky130_fd_sc_hd__and3_1
XFILLER_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_759 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18012__B1 _20081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11635__B1 _11633_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22765_ _22764_/A _22764_/B _22764_/C vssd1 vssd1 vccd1 vccd1 _22766_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18563__A1 _12522_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21716_ _23574_/Q _21716_/B _21716_/C vssd1 vssd1 vccd1 vccd1 _21716_/X sky130_fd_sc_hd__and3b_1
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20370__A1 _18335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22696_ _22611_/A _22611_/B _22685_/X vssd1 vssd1 vccd1 vccd1 _22729_/C sky130_fd_sc_hd__o21ai_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21647_ _21649_/C vssd1 vssd1 vccd1 vccd1 _21647_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12380_ _12377_/X _12378_/X _12379_/X _19082_/B _12327_/Y vssd1 vssd1 vccd1 vccd1
+ _12381_/A sky130_fd_sc_hd__a2111oi_2
XFILLER_197_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21578_ _21529_/X _21575_/Y _21694_/C _21614_/C _21614_/B vssd1 vssd1 vccd1 vccd1
+ _21579_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23317_ _23397_/CLK _23317_/D vssd1 vssd1 vccd1 vccd1 _23317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20529_ _20529_/A _20529_/B vssd1 vssd1 vccd1 vccd1 _20670_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14050_ _14050_/A vssd1 vssd1 vccd1 vccd1 _14050_/X sky130_fd_sc_hd__buf_2
XFILLER_158_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23248_ _23442_/Q input27/X _23250_/S vssd1 vssd1 vccd1 vccd1 _23249_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18618__A2 _18615_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16629__A1 _16064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ _13001_/A vssd1 vssd1 vccd1 vccd1 _13001_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17826__B1 _17943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23179_ _23179_/A vssd1 vssd1 vccd1 vccd1 _23411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input42_A x[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17740_ _17583_/B _17571_/Y _17575_/X _17566_/X vssd1 vssd1 vccd1 vccd1 _17759_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_48_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14952_ _14953_/B _14953_/C _14951_/X vssd1 vssd1 vccd1 vccd1 _14954_/A sky130_fd_sc_hd__a21bo_1
XFILLER_48_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13903_ _23350_/Q _23351_/Q vssd1 vssd1 vccd1 vccd1 _14013_/B sky130_fd_sc_hd__nor2_1
X_17671_ _17662_/A _17670_/Y _17668_/Y vssd1 vssd1 vccd1 vccd1 _17671_/X sky130_fd_sc_hd__a21bo_1
XFILLER_48_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14883_ _14883_/A _14883_/B _14883_/C vssd1 vssd1 vccd1 vccd1 _15459_/A sky130_fd_sc_hd__and3_1
XFILLER_48_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19410_ _19410_/A _19410_/B _19410_/C vssd1 vssd1 vccd1 vccd1 _19410_/X sky130_fd_sc_hd__and3_1
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16622_ _11960_/B _23595_/Q _16815_/D vssd1 vssd1 vccd1 vccd1 _16819_/A sky130_fd_sc_hd__a21oi_1
XFILLER_62_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13834_ _13834_/A _13834_/B _13834_/C vssd1 vssd1 vccd1 vccd1 _13834_/Y sky130_fd_sc_hd__nand3_2
XFILLER_47_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12418__A2 _19123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19341_ _19341_/A vssd1 vssd1 vccd1 vccd1 _19345_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16553_ _16554_/A _16554_/B _16551_/X _16552_/Y vssd1 vssd1 vccd1 vccd1 _16553_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ _13765_/A vssd1 vssd1 vccd1 vccd1 _13765_/X sky130_fd_sc_hd__buf_2
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ _15439_/B _15527_/A _15439_/A _15289_/C vssd1 vssd1 vccd1 vccd1 _15505_/B
+ sky130_fd_sc_hd__o31ai_1
X_19272_ _19298_/A _19298_/B _19272_/C vssd1 vssd1 vccd1 vccd1 _19442_/B sky130_fd_sc_hd__nand3_2
X_12716_ _21039_/B vssd1 vssd1 vccd1 vccd1 _12941_/A sky130_fd_sc_hd__buf_2
X_16484_ _16477_/B _16477_/C _16483_/Y _16518_/C vssd1 vssd1 vccd1 vccd1 _16495_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_13696_ _13698_/A _13698_/B _13593_/X vssd1 vssd1 vccd1 vccd1 _13697_/A sky130_fd_sc_hd__a21o_1
X_18223_ _18220_/X _18222_/X _18170_/D _18170_/Y vssd1 vssd1 vccd1 vccd1 _18223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15435_ _15435_/A _15435_/B vssd1 vssd1 vccd1 vccd1 _15435_/Y sky130_fd_sc_hd__nor2_1
X_12647_ _12637_/X _12640_/X _12724_/A vssd1 vssd1 vccd1 vccd1 _12648_/A sky130_fd_sc_hd__o21ai_1
XFILLER_15_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13430__A _13430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18154_ _18154_/A vssd1 vssd1 vccd1 vccd1 _18154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15366_ _15366_/A _15366_/B _15366_/C _15366_/D vssd1 vssd1 vccd1 vccd1 _15366_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12578_ _23289_/Q vssd1 vssd1 vccd1 vccd1 _13011_/C sky130_fd_sc_hd__clkinv_2
XFILLER_8_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16868__A1 _16592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17105_ _12208_/A _15655_/X _16856_/Y _17093_/Y _17096_/X vssd1 vssd1 vccd1 vccd1
+ _17106_/C sky130_fd_sc_hd__o221ai_1
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14317_ _14407_/D vssd1 vssd1 vccd1 vccd1 _15120_/B sky130_fd_sc_hd__clkbuf_2
X_18085_ _18085_/A _18085_/B vssd1 vssd1 vccd1 vccd1 _18106_/A sky130_fd_sc_hd__nand2_1
XFILLER_172_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15297_ _15455_/A _15350_/C _15298_/A vssd1 vssd1 vccd1 vccd1 _15299_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__16741__A _16741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17036_ _16749_/C _16917_/X _18335_/C _17035_/X vssd1 vssd1 vccd1 vccd1 _17036_/X
+ sky130_fd_sc_hd__a31o_1
X_14248_ _14245_/A _14245_/B _14347_/C vssd1 vssd1 vccd1 vccd1 _14248_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_125_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12354__A1 _12353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14179_ _14121_/B _14756_/A _14114_/X _14178_/Y _14174_/Y vssd1 vssd1 vccd1 vccd1
+ _14180_/C sky130_fd_sc_hd__o221ai_4
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20821__C1 _12692_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _11980_/Y _18812_/C _14646_/A _18998_/D vssd1 vssd1 vccd1 vccd1 _18989_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12106__A1 _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater102 _23497_/Q vssd1 vssd1 vccd1 vccd1 _14262_/A sky130_fd_sc_hd__clkbuf_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _18198_/C _18140_/B _17933_/X vssd1 vssd1 vccd1 vccd1 _17938_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__19034__A2 _17408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater113 _23391_/CLK vssd1 vssd1 vccd1 vccd1 _23300_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater124 _23444_/CLK vssd1 vssd1 vccd1 vccd1 _23347_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater135 _23352_/CLK vssd1 vssd1 vccd1 vccd1 _23358_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater146 _23307_/CLK vssd1 vssd1 vccd1 vccd1 _23372_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater157 _23321_/CLK vssd1 vssd1 vccd1 vccd1 _23325_/CLK sky130_fd_sc_hd__clkbuf_1
X_17869_ _17848_/X _17850_/Y _17852_/Y vssd1 vssd1 vccd1 vccd1 _17869_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_22_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16188__A _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19608_ _19598_/A _19598_/B _19598_/C _19607_/X vssd1 vssd1 vccd1 vccd1 _19609_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20880_ _20880_/A _21030_/B _21031_/A vssd1 vssd1 vccd1 vccd1 _20882_/A sky130_fd_sc_hd__nand3_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19539_ _19539_/A _19539_/B _19700_/C _19700_/D vssd1 vssd1 vccd1 vccd1 _19540_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22550_ _22493_/A _22544_/A _22493_/C vssd1 vssd1 vccd1 vccd1 _22550_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_107_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21501_ _21371_/C _21548_/B _21371_/B _21440_/C _21497_/A vssd1 vssd1 vccd1 vccd1
+ _21502_/C sky130_fd_sc_hd__a32o_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19011__B _19700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22481_ _22393_/B _22386_/Y _22567_/A _22283_/X vssd1 vssd1 vccd1 vccd1 _22489_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_22_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21432_ _21432_/A _21432_/B _21435_/C vssd1 vssd1 vccd1 vccd1 _21433_/B sky130_fd_sc_hd__nand3_1
XANTENNA__20104__A1 _19966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18848__A2 _11846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16859__A1 _15882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21363_ _21453_/B _21453_/C _21285_/C vssd1 vssd1 vccd1 vccd1 _21377_/A sky130_fd_sc_hd__a21bo_1
XFILLER_175_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23102_ _23377_/Q input26/X _23106_/S vssd1 vssd1 vccd1 vccd1 _23103_/A sky130_fd_sc_hd__mux2_1
X_20314_ _20366_/B vssd1 vssd1 vccd1 vccd1 _20314_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23054__A0 _14863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21294_ _21356_/A _21061_/X _21194_/B _21359_/A _21293_/Y vssd1 vssd1 vccd1 vccd1
+ _21298_/B sky130_fd_sc_hd__o221ai_1
XFILLER_122_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23033_ _23033_/A vssd1 vssd1 vccd1 vccd1 _23346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20245_ _20106_/C _20111_/C _20183_/B vssd1 vssd1 vccd1 vccd1 _20246_/A sky130_fd_sc_hd__a21oi_2
XFILLER_107_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18076__A3 _17406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16087__A2 _17414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20176_ _20176_/A _20176_/B _20176_/C vssd1 vssd1 vccd1 vccd1 _20176_/Y sky130_fd_sc_hd__nand3_1
XFILLER_118_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14098__A1 _14184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19025__A2 _11670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17036__A1 _16749_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11856__B1 _11807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16529__C _16529_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11880_ _11799_/X _11801_/X _18503_/C _18503_/D vssd1 vssd1 vccd1 vccd1 _11880_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22817_ _23282_/Q _22817_/B vssd1 vssd1 vccd1 vccd1 _22856_/D sky130_fd_sc_hd__or2_1
XANTENNA__21732__A _21732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__A2 _12906_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18536__A1 _11611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18536__B2 _12223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ _13697_/B _13697_/C vssd1 vssd1 vccd1 vccd1 _13550_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22748_ _22698_/Y _22731_/Y _22810_/B vssd1 vssd1 vccd1 vccd1 _22749_/C sky130_fd_sc_hd__o21bai_1
XFILLER_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12501_ _16620_/C vssd1 vssd1 vccd1 vccd1 _16795_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_41_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ _13634_/A _13634_/B _22159_/C vssd1 vssd1 vccd1 vccd1 _13482_/B sky130_fd_sc_hd__nand3_1
XFILLER_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22679_ _22675_/Y _22676_/Y _22678_/X vssd1 vssd1 vccd1 vccd1 _22679_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15220_ _15220_/A _15220_/B _15220_/C _15219_/B vssd1 vssd1 vccd1 vccd1 _15402_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_32_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12432_ _12432_/A vssd1 vssd1 vccd1 vccd1 _18435_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15770__A1 _12207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15151_ _15129_/A _15129_/B _15130_/C vssd1 vssd1 vccd1 vccd1 _15193_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__19500__A3 _19858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12363_ _12363_/A _12363_/B _12363_/C _12363_/D vssd1 vssd1 vccd1 vccd1 _12372_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_5_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _14099_/X _14976_/A _14101_/Y vssd1 vssd1 vccd1 vccd1 _14164_/B sky130_fd_sc_hd__a21oi_2
XFILLER_165_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23045__A0 _13945_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15082_ _15155_/A _15082_/B _15356_/A _15082_/D vssd1 vssd1 vccd1 vccd1 _15082_/Y
+ sky130_fd_sc_hd__nand4_2
X_12294_ _12297_/B _12297_/C _12292_/X _12293_/Y vssd1 vssd1 vccd1 vccd1 _12298_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_10_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18910_ _18910_/A _18910_/B _18910_/C vssd1 vssd1 vccd1 vccd1 _18921_/A sky130_fd_sc_hd__nand3_1
X_14033_ _14015_/B _14029_/X _14429_/A _14312_/B vssd1 vssd1 vccd1 vccd1 _14121_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19890_ _19897_/A _19897_/B vssd1 vssd1 vccd1 vccd1 _19896_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_72 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18841_ _18841_/A _18841_/B vssd1 vssd1 vccd1 vccd1 _18841_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18472__B1 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18772_ _18969_/A _18966_/A _18966_/B vssd1 vssd1 vccd1 vccd1 _18773_/D sky130_fd_sc_hd__nand3_2
X_15984_ _15843_/B _16123_/A _19017_/D _16840_/A _16172_/A vssd1 vssd1 vccd1 vccd1
+ _15985_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_94_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17723_ _17723_/A _17723_/B _17723_/C vssd1 vssd1 vccd1 vccd1 _17724_/B sky130_fd_sc_hd__and3_1
XFILLER_94_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14935_ _14936_/B _15044_/C _14805_/B _14928_/B _14934_/X vssd1 vssd1 vccd1 vccd1
+ _14939_/A sky130_fd_sc_hd__a221oi_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21374__A3 _21635_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13425__A _22521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17654_ _17654_/A _17654_/B vssd1 vssd1 vccd1 vccd1 _17654_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14866_ _14879_/C _14864_/Y _14970_/B _23362_/Q vssd1 vssd1 vccd1 vccd1 _15094_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19319__A3 _19172_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16605_ _15698_/A _15698_/B _17626_/A _16058_/A _11936_/X vssd1 vssd1 vccd1 vccd1
+ _16605_/X sky130_fd_sc_hd__o32a_1
X_13817_ _21764_/C _21877_/A _13818_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13819_/A
+ sky130_fd_sc_hd__a22oi_2
X_17585_ _17585_/A _17585_/B _17585_/C vssd1 vssd1 vccd1 vccd1 _17609_/B sky130_fd_sc_hd__nand3_4
XFILLER_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14797_ _14797_/A _14797_/B _14797_/C vssd1 vssd1 vccd1 vccd1 _14797_/X sky130_fd_sc_hd__and3_1
XFILLER_90_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19324_ _19491_/A _19491_/B _19314_/Y _19525_/A _19524_/A vssd1 vssd1 vccd1 vccd1
+ _19477_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16536_ _17035_/C _16536_/B _17450_/C _17326_/D vssd1 vssd1 vccd1 vccd1 _16536_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_189_764 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16538__B1 _16539_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13748_ _13715_/X _13748_/B _13748_/C vssd1 vssd1 vccd1 vccd1 _13748_/Y sky130_fd_sc_hd__nand3b_1
XANTENNA__17735__C1 _17259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19255_ _19236_/Y _19245_/X _19254_/Y vssd1 vssd1 vccd1 vccd1 _19259_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16467_ _16467_/A _16467_/B _16467_/C vssd1 vssd1 vccd1 vccd1 _16539_/B sky130_fd_sc_hd__nand3_2
XFILLER_176_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13679_ _13680_/A _13680_/B _13680_/C _13680_/D vssd1 vssd1 vccd1 vccd1 _13679_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18206_ _18206_/A _18262_/B vssd1 vssd1 vccd1 vccd1 _23592_/D sky130_fd_sc_hd__xor2_2
XFILLER_176_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15418_ _15446_/C _15419_/C _15419_/D _15419_/B _15446_/D vssd1 vssd1 vccd1 vccd1
+ _15420_/A sky130_fd_sc_hd__a32o_1
XFILLER_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19186_ _19186_/A _19186_/B vssd1 vssd1 vccd1 vccd1 _19186_/Y sky130_fd_sc_hd__nand2_1
X_16398_ _16398_/A vssd1 vssd1 vccd1 vccd1 _16398_/X sky130_fd_sc_hd__buf_2
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_992 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18137_ _18137_/A _18252_/A vssd1 vssd1 vccd1 vccd1 _18141_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15349_ _15298_/B _15109_/X _15110_/X _15348_/Y _15324_/A vssd1 vssd1 vccd1 vccd1
+ _15350_/A sky130_fd_sc_hd__a311o_1
XFILLER_89_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19485__C _19700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22192__B _22554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18068_ _18068_/A vssd1 vssd1 vccd1 vccd1 _23590_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17019_ _17019_/A _17019_/B _17019_/C vssd1 vssd1 vccd1 vccd1 _17381_/B sky130_fd_sc_hd__nand3_1
XFILLER_144_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12504__A _23593_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17266__A1 _17260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16069__A2 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20030_ _20028_/Y _20029_/Y _23549_/Q vssd1 vssd1 vccd1 vccd1 _20042_/A sky130_fd_sc_hd__a21boi_1
XFILLER_113_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20270__B1 _18211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_328 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13827__A1 _13495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21981_ _21981_/A _21981_/B _21981_/C vssd1 vssd1 vccd1 vccd1 _22106_/B sky130_fd_sc_hd__nand3_1
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18766__B2 _18604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13335__A _23323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20932_ _20778_/X _20934_/A _20783_/Y _20790_/B vssd1 vssd1 vccd1 vccd1 _20937_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16241__A2 _16281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20863_ _20863_/A _20885_/B vssd1 vssd1 vccd1 vccd1 _20863_/Y sky130_fd_sc_hd__nand2_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22602_ _22509_/A _22509_/B _22505_/B vssd1 vssd1 vccd1 vccd1 _22602_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__21271__B _21271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23582_ _23582_/CLK _23582_/D vssd1 vssd1 vccd1 vccd1 _23582_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12263__B1 _12214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20794_ _20794_/A _20794_/B _20794_/C vssd1 vssd1 vccd1 vccd1 _20819_/B sky130_fd_sc_hd__nand3_2
XFILLER_179_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16365__B _16821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22533_ _22532_/A _22530_/A _23277_/Q vssd1 vssd1 vccd1 vccd1 _22533_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_762 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19957__A _19957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__B1 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19479__C1 _18503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22464_ _22271_/A _22271_/B _22475_/B vssd1 vssd1 vccd1 vccd1 _22473_/A sky130_fd_sc_hd__o21ai_1
XFILLER_33_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21415_ _21415_/A vssd1 vssd1 vccd1 vccd1 _21617_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22395_ _22383_/X _22389_/Y _22394_/Y vssd1 vssd1 vccd1 vccd1 _22395_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_135_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15402__D_N _15442_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1056 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12117__C _19165_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21346_ _21346_/A vssd1 vssd1 vccd1 vccd1 _21346_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_878 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15504__A1 _15439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21277_ _21277_/A vssd1 vssd1 vccd1 vccd1 _21502_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22830__B _22830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23016_ _23016_/A vssd1 vssd1 vccd1 vccd1 _23338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20228_ _20283_/C _20283_/A _20283_/B vssd1 vssd1 vccd1 vccd1 _20228_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20159_ _20159_/A _20159_/B _20159_/C vssd1 vssd1 vccd1 vccd1 _20232_/A sky130_fd_sc_hd__nand3_2
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12143__B1_N _12104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _13186_/C _12981_/B _12981_/C vssd1 vssd1 vccd1 vccd1 _12981_/X sky130_fd_sc_hd__and3_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14491__A1 _14298_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19954__B1 _20081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _23413_/Q _14640_/A _14534_/X _23445_/Q _14719_/X vssd1 vssd1 vccd1 vccd1
+ _14720_/X sky130_fd_sc_hd__a221o_4
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ _12256_/A vssd1 vssd1 vccd1 vccd1 _18531_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22558__A _22558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18755__B _18755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14651_ _16657_/B vssd1 vssd1 vccd1 vccd1 _16780_/B sky130_fd_sc_hd__buf_6
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11863_ _12017_/A _12019_/A _11887_/C _11887_/A vssd1 vssd1 vccd1 vccd1 _12016_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15440__B1 _15439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19706__B1 _19218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _13602_/A _23324_/Q _13602_/C vssd1 vssd1 vccd1 vccd1 _13602_/Y sky130_fd_sc_hd__nor3_2
XANTENNA__20316__A1 _18211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17370_ _17832_/A _17522_/B _17522_/C _17522_/D vssd1 vssd1 vccd1 vccd1 _17372_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _11665_/A _23112_/D _23184_/D _15664_/A vssd1 vssd1 vccd1 vccd1 _14582_/X
+ sky130_fd_sc_hd__a22o_1
X_11794_ _18973_/C vssd1 vssd1 vccd1 vccd1 _19157_/C sky130_fd_sc_hd__buf_2
XFILLER_198_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16321_ _16321_/A _16321_/B vssd1 vssd1 vccd1 vccd1 _16397_/B sky130_fd_sc_hd__nand2_2
XFILLER_14_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13533_ _13544_/A _13544_/B _13545_/A vssd1 vssd1 vccd1 vccd1 _13535_/A sky130_fd_sc_hd__and3_1
XANTENNA__18771__A _18771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19040_ _19040_/A vssd1 vssd1 vccd1 vccd1 _19040_/X sky130_fd_sc_hd__buf_2
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13464_ _13513_/A _13517_/A _13517_/C vssd1 vssd1 vccd1 vccd1 _13476_/A sky130_fd_sc_hd__a21boi_1
X_16252_ _16240_/Y _16251_/X _16242_/A _16242_/B vssd1 vssd1 vccd1 vccd1 _16254_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16940__B1 _16706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15203_ _15203_/A _15203_/B _15277_/A vssd1 vssd1 vccd1 vccd1 _15277_/B sky130_fd_sc_hd__nand3_2
X_12415_ _19155_/B _19155_/C _12410_/C _18440_/A vssd1 vssd1 vccd1 vccd1 _19804_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_12_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13395_ _13323_/X _13338_/X _13354_/C _13354_/B _13394_/Y vssd1 vssd1 vccd1 vccd1
+ _13620_/B sky130_fd_sc_hd__a41oi_4
X_16183_ _16183_/A vssd1 vssd1 vccd1 vccd1 _16183_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_127_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15320__A1_N _15366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12346_ _12346_/A vssd1 vssd1 vccd1 vccd1 _16528_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__21292__A2 _20504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15134_ _15080_/X _15134_/B _15134_/C vssd1 vssd1 vccd1 vccd1 _15136_/B sky130_fd_sc_hd__nand3b_1
XFILLER_142_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12309__B2 _12508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19942_ _19888_/A _19888_/B _19888_/D vssd1 vssd1 vccd1 vccd1 _19942_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_175_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15065_ _15065_/A _15065_/B _15065_/C vssd1 vssd1 vccd1 vccd1 _15065_/Y sky130_fd_sc_hd__nand3_2
X_12277_ _12275_/Y _12276_/X _11805_/A vssd1 vssd1 vccd1 vccd1 _12297_/C sky130_fd_sc_hd__o21bai_2
XANTENNA__12324__A _12324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14016_ _14120_/A vssd1 vssd1 vccd1 vccd1 _14243_/A sky130_fd_sc_hd__buf_2
XANTENNA__14242__C _15415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output73_A _14708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19873_ _19873_/A _19873_/B _19873_/C vssd1 vssd1 vccd1 vccd1 _19888_/D sky130_fd_sc_hd__nand3_2
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18824_ _19011_/A _19019_/B _19539_/B vssd1 vssd1 vccd1 vccd1 _18825_/B sky130_fd_sc_hd__and3_1
XFILLER_110_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18755_ _18755_/A _18755_/B _18755_/C _18755_/D vssd1 vssd1 vccd1 vccd1 _18755_/Y
+ sky130_fd_sc_hd__nand4_4
X_15967_ _15998_/A _15998_/B vssd1 vssd1 vccd1 vccd1 _16000_/A sky130_fd_sc_hd__xnor2_4
XFILLER_67_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16208__C1 _16866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17706_ _17514_/C _17705_/Y _17686_/X _17541_/Y vssd1 vssd1 vccd1 vccd1 _17821_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_76_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14918_ _14918_/A _14918_/B _14918_/C vssd1 vssd1 vccd1 vccd1 _14923_/C sky130_fd_sc_hd__nand3_1
XFILLER_48_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18686_ _12214_/X _17627_/A _18677_/Y _18678_/Y vssd1 vssd1 vccd1 vccd1 _18687_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15898_ _15773_/Y _15775_/X _15946_/A vssd1 vssd1 vccd1 vccd1 _15898_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_707 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17637_ _17637_/A _17637_/B _17637_/C vssd1 vssd1 vccd1 vccd1 _17792_/A sky130_fd_sc_hd__nand3_2
X_14849_ _14846_/Y _14847_/Y _14845_/Y _14848_/X vssd1 vssd1 vccd1 vccd1 _14849_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17568_ _17435_/X _17434_/X _16056_/X _17567_/X vssd1 vssd1 vccd1 vccd1 _17575_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_189_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19173__A1 _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19199__D _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19307_ _12018_/X _12020_/X _19308_/C _19163_/A vssd1 vssd1 vccd1 vccd1 _19307_/Y
+ sky130_fd_sc_hd__o211ai_4
X_16519_ _16471_/Y _16518_/Y _16512_/Y vssd1 vssd1 vccd1 vccd1 _16519_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_17_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17499_ _17154_/X _17155_/X _17152_/B _17161_/B vssd1 vssd1 vccd1 vccd1 _17499_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19238_ _19060_/B _19057_/D _19066_/Y _19065_/X vssd1 vssd1 vccd1 vccd1 _19244_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_31_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20138__D _20320_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19169_ _11898_/X _19838_/A _19162_/A vssd1 vssd1 vccd1 vccd1 _19172_/A sky130_fd_sc_hd__o21ai_4
XFILLER_157_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21200_ _21194_/Y _21307_/A _21356_/A _12862_/X vssd1 vssd1 vccd1 vccd1 _21202_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_144_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18684__B1 _12464_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22180_ _14614_/X _22047_/B _22141_/C _21853_/A vssd1 vssd1 vccd1 vccd1 _22560_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__21283__A2 _21432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14433__B _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21131_ _21131_/A _21131_/B vssd1 vssd1 vccd1 vccd1 _21132_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22232__A1 _21988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21062_ _20639_/C _12689_/X _12640_/X _12692_/Y _13056_/X vssd1 vssd1 vccd1 vccd1
+ _21062_/X sky130_fd_sc_hd__a311o_1
XFILLER_28_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20013_ _20013_/A _20013_/B vssd1 vssd1 vccd1 vccd1 _20013_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19017__A _19017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11792__B _11792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14473__A1 _14108_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21964_ _21964_/A _21964_/B _21964_/C vssd1 vssd1 vccd1 vccd1 _21965_/C sky130_fd_sc_hd__nand3_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17411__A1 _17408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16214__A2 _12020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20915_ _20911_/X _20914_/Y _20909_/X _20900_/Y vssd1 vssd1 vccd1 vccd1 _20943_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21895_ _21753_/B _21750_/Y _21906_/A _13793_/B vssd1 vssd1 vccd1 vccd1 _21911_/A
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16376__A _19503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23569__CLK _23582_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20846_ _20846_/A _20847_/A _20847_/B vssd1 vssd1 vccd1 vccd1 _20846_/Y sky130_fd_sc_hd__nand3_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15973__A1 _15855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_55 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16095__B _16326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23565_ _23566_/CLK _23565_/D vssd1 vssd1 vccd1 vccd1 _23565_/Q sky130_fd_sc_hd__dfxtp_1
X_20777_ _20770_/X _20772_/X _21000_/B vssd1 vssd1 vccd1 vccd1 _20846_/A sky130_fd_sc_hd__o21ai_1
XFILLER_196_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22516_ _22516_/A _22516_/B _22516_/C _22516_/D vssd1 vssd1 vccd1 vccd1 _22607_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_156_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23496_ _23499_/CLK _23496_/D vssd1 vssd1 vccd1 vccd1 _23496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22447_ _22447_/A _22447_/B vssd1 vssd1 vccd1 vccd1 _22448_/B sky130_fd_sc_hd__nor2_1
XFILLER_183_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14624__A _23298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ _12227_/B _12200_/B vssd1 vssd1 vccd1 vccd1 _12387_/A sky130_fd_sc_hd__nand2_1
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22471__A1 _13470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ _13181_/A _13176_/C _13176_/A _13168_/A _13159_/X vssd1 vssd1 vccd1 vccd1
+ _13180_/X sky130_fd_sc_hd__a32o_1
X_22378_ _22381_/A vssd1 vssd1 vccd1 vccd1 _22637_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15439__B _15439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12131_ _12131_/A _12425_/A vssd1 vssd1 vccd1 vccd1 _12131_/Y sky130_fd_sc_hd__nor2_1
X_21329_ _21320_/Y _21328_/Y _21311_/A vssd1 vssd1 vccd1 vccd1 _21330_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__19219__A2 _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12144__A _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22560__B _22560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12062_ _12391_/B _12251_/B vssd1 vssd1 vccd1 vccd1 _12392_/C sky130_fd_sc_hd__nor2_1
XFILLER_150_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16870_ _16870_/A _16870_/B _16870_/C vssd1 vssd1 vccd1 vccd1 _16890_/B sky130_fd_sc_hd__nand3_2
XFILLER_1_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15256__A3 _15353_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15821_ _15821_/A vssd1 vssd1 vccd1 vccd1 _16451_/B sky130_fd_sc_hd__buf_2
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18540_ _18540_/A _18540_/B _18540_/C vssd1 vssd1 vccd1 vccd1 _18541_/A sky130_fd_sc_hd__and3_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_73 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _16856_/A _16856_/B _15968_/A vssd1 vssd1 vccd1 vccd1 _15753_/B sky130_fd_sc_hd__nand3_4
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _13119_/B vssd1 vssd1 vccd1 vccd1 _20563_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17402__A1 _17134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21192__A _21493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14703_ _23344_/Q _14689_/X _14694_/X _23312_/Q _14699_/X vssd1 vssd1 vccd1 vccd1
+ _14703_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11915_ _11915_/A vssd1 vssd1 vccd1 vccd1 _12089_/A sky130_fd_sc_hd__buf_2
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _18475_/A _18483_/A _18478_/A vssd1 vssd1 vccd1 vccd1 _18490_/A sky130_fd_sc_hd__o21ai_4
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15683_ _16030_/A _11654_/A _15682_/Y vssd1 vssd1 vccd1 vccd1 _15783_/A sky130_fd_sc_hd__o21ai_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16286__A _16860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12895_ _12893_/Y _12894_/X _12900_/A _13034_/A vssd1 vssd1 vccd1 vccd1 _12896_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_166_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _17625_/C vssd1 vssd1 vccd1 vccd1 _17959_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _14688_/A vssd1 vssd1 vccd1 vccd1 _14635_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11846_ _11846_/A vssd1 vssd1 vccd1 vccd1 _19218_/A sky130_fd_sc_hd__buf_2
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _17361_/B _17514_/A _17359_/B vssd1 vssd1 vccd1 vccd1 _17353_/Y sky130_fd_sc_hd__a21oi_4
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14565_ _14188_/C _14545_/A _14539_/X _11743_/A vssd1 vssd1 vccd1 vccd1 _14565_/X
+ sky130_fd_sc_hd__a22o_1
X_11777_ _11720_/A _11644_/C _11694_/X _11733_/Y _11634_/B vssd1 vssd1 vccd1 vccd1
+ _11882_/A sky130_fd_sc_hd__o311ai_4
XANTENNA__12319__A _18941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _12146_/X _12147_/X _15742_/X _16447_/B _12149_/A vssd1 vssd1 vccd1 vccd1
+ _16304_/Y sky130_fd_sc_hd__o221ai_1
X_13516_ _13516_/A _13516_/B vssd1 vssd1 vccd1 vccd1 _13517_/B sky130_fd_sc_hd__xor2_1
X_17284_ _17260_/Y _17263_/Y _17960_/A _17974_/D vssd1 vssd1 vccd1 vccd1 _17284_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_929 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14496_ _14496_/A _14496_/B vssd1 vssd1 vccd1 vccd1 _14497_/C sky130_fd_sc_hd__nand2_1
XFILLER_173_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19023_ _11814_/A _18452_/A _12105_/Y _18835_/A vssd1 vssd1 vccd1 vccd1 _19029_/D
+ sky130_fd_sc_hd__o22ai_4
XFILLER_173_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16235_ _16242_/B vssd1 vssd1 vccd1 vccd1 _16725_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13447_ _13458_/C _13447_/B _13447_/C vssd1 vssd1 vccd1 vccd1 _13448_/A sky130_fd_sc_hd__nand3b_1
XFILLER_127_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21265__A2 _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22462__A1 _13470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16166_ _19381_/B vssd1 vssd1 vccd1 vccd1 _20062_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13378_ _13785_/C vssd1 vssd1 vccd1 vccd1 _13602_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_155_984 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15117_ _15233_/A _15233_/B _15118_/A _15257_/B vssd1 vssd1 vccd1 vccd1 _15120_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17845__A _19534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12329_ _12346_/A _18755_/A _18755_/B _19512_/D _12327_/A vssd1 vssd1 vccd1 vccd1
+ _12329_/X sky130_fd_sc_hd__a32o_1
XFILLER_173_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16097_ _16020_/X _16073_/Y _16335_/A _16063_/X vssd1 vssd1 vccd1 vccd1 _16097_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18418__B1 _18154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19925_ _19925_/A _19925_/B vssd1 vssd1 vccd1 vccd1 _20032_/A sky130_fd_sc_hd__nand2_2
X_15048_ _15045_/A _15045_/B _15050_/A _15050_/B vssd1 vssd1 vccd1 vccd1 _15049_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16692__A2 _16055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12989__A _23456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11893__A _15718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19856_ _19480_/X _19659_/Y _19667_/B _19943_/A _19943_/B vssd1 vssd1 vccd1 vccd1
+ _19856_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_69_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18807_ _12130_/X _19184_/A _18796_/X _18790_/X _18792_/Y vssd1 vssd1 vccd1 vccd1
+ _18808_/C sky130_fd_sc_hd__o221ai_4
X_19787_ _23547_/Q _19787_/B _19787_/C vssd1 vssd1 vccd1 vccd1 _19788_/C sky130_fd_sc_hd__nand3b_1
X_16999_ _16998_/B _16998_/C _17022_/A _16777_/Y vssd1 vssd1 vccd1 vccd1 _17017_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__14455__B2 _15094_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18738_ _23541_/Q _18738_/B _18738_/C vssd1 vssd1 vccd1 vccd1 _18747_/B sky130_fd_sc_hd__nand3b_1
XFILLER_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18669_ _18669_/A _18669_/B _18669_/C _18669_/D vssd1 vssd1 vccd1 vccd1 _18868_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA__14207__A1 _14031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20700_ _20715_/C _20718_/A _20718_/B vssd1 vssd1 vccd1 vccd1 _20700_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21680_ _21665_/Y _21679_/X _21704_/C _21694_/A vssd1 vssd1 vccd1 vccd1 _21691_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21830__A _23481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20631_ _20631_/A vssd1 vssd1 vccd1 vccd1 _20631_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17157__B1 _17152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19697__A2 _19800_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22150__B1 _13486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23350_ _23352_/CLK _23350_/D vssd1 vssd1 vccd1 vccd1 _23350_/Q sky130_fd_sc_hd__dfxtp_1
X_20562_ _20562_/A _20562_/B vssd1 vssd1 vccd1 vccd1 _20566_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13051__C _13051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13981__A3 _13985_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22301_ _22644_/A _13599_/X _22122_/Y _22362_/A _22297_/Y vssd1 vssd1 vccd1 vccd1
+ _22301_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_149_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22364__C _22637_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14915__C1 _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23281_ _23510_/CLK _23281_/D vssd1 vssd1 vccd1 vccd1 _23281_/Q sky130_fd_sc_hd__dfxtp_1
X_20493_ _23289_/Q _20493_/B _23287_/Q _20493_/D vssd1 vssd1 vccd1 vccd1 _20798_/A
+ sky130_fd_sc_hd__nor4_2
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_567 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1162 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22232_ _21988_/A _22226_/B _21988_/B _22670_/D _22223_/X vssd1 vssd1 vccd1 vccd1
+ _22232_/X sky130_fd_sc_hd__a41o_1
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22163_ _22035_/X _22025_/Y _22040_/Y vssd1 vssd1 vccd1 vccd1 _22166_/B sky130_fd_sc_hd__o21ai_2
XFILLER_132_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21114_ _21134_/A vssd1 vssd1 vccd1 vccd1 _21236_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22094_ _22094_/A _22094_/B _22094_/C vssd1 vssd1 vccd1 vccd1 _22240_/A sky130_fd_sc_hd__nand3_1
XFILLER_132_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12899__A _12899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19970__A _20142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21045_ _21045_/A _21045_/B _21045_/C vssd1 vssd1 vccd1 vccd1 _21084_/A sky130_fd_sc_hd__nand3_2
XFILLER_87_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19621__A2 _20368_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11901__C1 _19548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17093__C1 _17712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_787 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22996_ _22996_/A vssd1 vssd1 vccd1 vccd1 _23329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21947_ _21947_/A vssd1 vssd1 vccd1 vccd1 _22089_/A sky130_fd_sc_hd__buf_2
XFILLER_131_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11700_ _15699_/A vssd1 vssd1 vccd1 vccd1 _16674_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13523__A _13523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12680_/A vssd1 vssd1 vccd1 vccd1 _12704_/A sky130_fd_sc_hd__clkbuf_4
X_21878_ _21878_/A _22263_/B _22226_/C vssd1 vssd1 vccd1 vccd1 _21878_/X sky130_fd_sc_hd__and3_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _18947_/B vssd1 vssd1 vccd1 vccd1 _11915_/A sky130_fd_sc_hd__clkinv_2
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ _12957_/Y _12815_/B _12714_/X _20961_/A _12936_/A vssd1 vssd1 vccd1 vccd1
+ _20829_/X sky130_fd_sc_hd__o32a_1
XFILLER_39_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19210__A _19210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14350_ _14403_/A _14350_/B _14350_/C _14350_/D vssd1 vssd1 vccd1 vccd1 _14414_/A
+ sky130_fd_sc_hd__nand4_2
X_23548_ _23578_/CLK _23548_/D vssd1 vssd1 vccd1 vccd1 _23548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13301_ _13585_/A _21891_/A _22558_/A _13736_/B vssd1 vssd1 vccd1 vccd1 _13303_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14281_ _13942_/X _13969_/Y _14245_/A vssd1 vssd1 vccd1 vccd1 _14361_/C sky130_fd_sc_hd__o21ai_1
X_23479_ _23510_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 _23479_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13232_ _13339_/A vssd1 vssd1 vccd1 vccd1 _22022_/A sky130_fd_sc_hd__clkbuf_4
X_16020_ _16020_/A _16020_/B _16020_/C vssd1 vssd1 vccd1 vccd1 _16020_/X sky130_fd_sc_hd__and3_2
XFILLER_196_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19845__C1 _17406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13163_ _21054_/C vssd1 vssd1 vccd1 vccd1 _21172_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12114_ _11684_/A _11828_/B _12113_/X vssd1 vssd1 vccd1 vccd1 _12114_/Y sky130_fd_sc_hd__a21oi_1
X_17971_ _19534_/B vssd1 vssd1 vccd1 vccd1 _19967_/C sky130_fd_sc_hd__buf_2
X_13094_ _20769_/A vssd1 vssd1 vccd1 vccd1 _21490_/B sky130_fd_sc_hd__buf_2
XFILLER_124_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19710_ _19710_/A _19819_/B vssd1 vssd1 vccd1 vccd1 _19713_/A sky130_fd_sc_hd__nand2_1
X_16922_ _16923_/C _16917_/X _16923_/A vssd1 vssd1 vccd1 vccd1 _16922_/Y sky130_fd_sc_hd__a21oi_1
X_12045_ _12002_/Y _12007_/Y _19512_/C _19381_/D _12166_/A vssd1 vssd1 vccd1 vccd1
+ _12046_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_78_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19612__A2 _20371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12602__A _13052_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19641_ _19588_/Y _19587_/C _19596_/X _19583_/Y vssd1 vssd1 vccd1 vccd1 _19641_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_66_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16853_ _16853_/A _16853_/B _16853_/C vssd1 vssd1 vccd1 vccd1 _16894_/B sky130_fd_sc_hd__nand3_1
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15804_ _15644_/X _16668_/C _15639_/C vssd1 vssd1 vccd1 vccd1 _15804_/Y sky130_fd_sc_hd__a21oi_1
X_19572_ _19572_/A vssd1 vssd1 vccd1 vccd1 _19572_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14988__A2 _15422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16784_ _16784_/A vssd1 vssd1 vccd1 vccd1 _16784_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13996_ _15353_/A _15353_/B _14252_/D _14791_/C _14867_/C vssd1 vssd1 vccd1 vccd1
+ _13996_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_74_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18523_ _18523_/A _18529_/A _18529_/B vssd1 vssd1 vccd1 vccd1 _18523_/Y sky130_fd_sc_hd__nand3_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735_ _15662_/B _15735_/B _15735_/C vssd1 vssd1 vccd1 vccd1 _15736_/A sky130_fd_sc_hd__and3b_4
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12947_ _20663_/D vssd1 vssd1 vccd1 vccd1 _20905_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__21183__A1 _12571_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _18461_/B vssd1 vssd1 vccd1 vccd1 _18455_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_179_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15666_ _16684_/A vssd1 vssd1 vccd1 vccd1 _15918_/C sky130_fd_sc_hd__clkbuf_4
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20930__A1 _12709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ _12674_/A _12935_/A _12877_/Y vssd1 vssd1 vccd1 vccd1 _12894_/B sky130_fd_sc_hd__o21ai_2
XFILLER_33_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17405_ _17493_/A _17493_/B _17405_/C vssd1 vssd1 vccd1 vccd1 _17663_/B sky130_fd_sc_hd__nand3_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14617_ _23582_/Q _14551_/A _14587_/X _14879_/C vssd1 vssd1 vccd1 vccd1 _14617_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18385_ _18345_/A _18388_/B _18344_/B vssd1 vssd1 vccd1 vccd1 _18385_/X sky130_fd_sc_hd__o21ba_1
X_11829_ _12118_/C vssd1 vssd1 vccd1 vccd1 _11849_/C sky130_fd_sc_hd__buf_2
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15597_ _23418_/Q _23419_/Q vssd1 vssd1 vccd1 vccd1 _15614_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22465__B _22554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17336_ _17336_/A _17336_/B _17336_/C vssd1 vssd1 vccd1 vccd1 _17350_/C sky130_fd_sc_hd__nand3_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14548_ _13945_/X _14545_/X _14547_/X _12788_/B vssd1 vssd1 vccd1 vccd1 _14548_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17267_ _17267_/A _17267_/B _17267_/C vssd1 vssd1 vccd1 vccd1 _17268_/C sky130_fd_sc_hd__nand3_2
XANTENNA__16362__A1 _16360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14479_ _14445_/Y _14441_/Y _14468_/A _14453_/Y vssd1 vssd1 vccd1 vccd1 _14483_/A
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__12286__A1_N _12297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19006_ _19210_/A _19191_/A _19013_/A _19703_/A _19180_/D vssd1 vssd1 vccd1 vccd1
+ _19007_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_134_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14373__B1 _14097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16218_ _16215_/Y _16201_/X _16216_/Y _16217_/Y vssd1 vssd1 vccd1 vccd1 _16710_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_174_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17198_ _16946_/X _16942_/X _17187_/A _17187_/B vssd1 vssd1 vccd1 vccd1 _17198_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__23264__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16149_ _16447_/A _15766_/X _16612_/B _16612_/C vssd1 vssd1 vccd1 vccd1 _16614_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_142_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19908_ _19900_/X _19903_/X _19899_/Y _19894_/Y vssd1 vssd1 vccd1 vccd1 _19909_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__12512__A _16807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_862 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14430__C _15238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19839_ _20081_/D vssd1 vssd1 vccd1 vccd1 _20263_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16968__A3 _16749_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14979__A2 _14097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22850_ _22848_/Y _22849_/X _23283_/Q vssd1 vssd1 vccd1 vccd1 _22850_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__19367__A1 _19040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23462__D _23474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21801_ _21801_/A _21801_/B _21801_/C vssd1 vssd1 vccd1 vccd1 _21804_/A sky130_fd_sc_hd__and3_1
X_22781_ _22529_/A _22777_/Y _22780_/Y vssd1 vssd1 vccd1 vccd1 _22783_/B sky130_fd_sc_hd__o21a_1
XFILLER_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21732_ _21732_/A vssd1 vssd1 vccd1 vccd1 _22107_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_334 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19949__B _20217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19119__A1 _17591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19119__B2 _12282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18853__B _18959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16050__B1 _16046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21663_ _23573_/Q vssd1 vssd1 vccd1 vccd1 _21691_/A sky130_fd_sc_hd__inv_2
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14600__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14600__B2 _14599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20614_ _20614_/A _20614_/B vssd1 vssd1 vccd1 vccd1 _20614_/Y sky130_fd_sc_hd__nand2_1
X_23402_ _23402_/CLK _23402_/D vssd1 vssd1 vccd1 vccd1 _23402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21594_ _21594_/A _21594_/B vssd1 vssd1 vccd1 vccd1 _21595_/B sky130_fd_sc_hd__nor2_1
XFILLER_177_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23333_ _23429_/CLK _23333_/D vssd1 vssd1 vccd1 vccd1 _23333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20545_ _20534_/X _20540_/X _20552_/A vssd1 vssd1 vccd1 vccd1 _20713_/B sky130_fd_sc_hd__o21ai_2
XFILLER_192_342 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23264_ _23584_/CLK _23264_/D vssd1 vssd1 vccd1 vccd1 _23264_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_165_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20476_ _20625_/A _20621_/A _20634_/A vssd1 vssd1 vccd1 vccd1 _20490_/A sky130_fd_sc_hd__o21ai_1
XFILLER_180_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20904__A _21054_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22215_ _22215_/A _22215_/B vssd1 vssd1 vccd1 vccd1 _22215_/X sky130_fd_sc_hd__or2_1
XFILLER_193_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23195_ _14569_/X input33/X _23195_/S vssd1 vssd1 vccd1 vccd1 _23196_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19842__A2 _19504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22146_ _22562_/A vssd1 vssd1 vccd1 vccd1 _22569_/A sky130_fd_sc_hd__buf_2
XFILLER_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22077_ _22218_/A _22220_/D _22218_/B vssd1 vssd1 vccd1 vccd1 _22077_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12422__A _19512_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21028_ _21028_/A _21028_/B vssd1 vssd1 vccd1 vccd1 _23543_/D sky130_fd_sc_hd__xnor2_1
XFILLER_102_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15733__A _15860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ _13686_/A _21987_/B _13848_/Y _13849_/Y vssd1 vssd1 vccd1 vccd1 _13857_/A
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__19358__A1 _17742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19358__B2 _12184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22269__C _22269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ _13119_/A _13119_/B _20962_/B _20669_/C vssd1 vssd1 vccd1 vccd1 _12801_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13781_ _13453_/A _13444_/A _13610_/Y _13609_/X vssd1 vssd1 vccd1 vccd1 _13781_/X
+ sky130_fd_sc_hd__o22a_1
X_22979_ _13264_/C input33/X _22979_/S vssd1 vssd1 vccd1 vccd1 _22980_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13253__A _13253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15520_ _15521_/B _15520_/B vssd1 vssd1 vccd1 vccd1 _15522_/A sky130_fd_sc_hd__and2b_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12677_/X _12704_/X _13003_/B _12705_/X vssd1 vssd1 vccd1 vccd1 _12733_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15171__C _15233_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22566__A _22566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15451_ _15427_/A _15451_/B _15451_/C _15451_/D vssd1 vssd1 vccd1 vccd1 _15462_/A
+ sky130_fd_sc_hd__and4b_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12663_ _12776_/A vssd1 vssd1 vccd1 vccd1 _13138_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _14439_/C _14410_/B vssd1 vssd1 vccd1 vccd1 _14405_/A sky130_fd_sc_hd__nand2_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18170_ _18170_/A _18217_/A _18272_/A _18170_/D vssd1 vssd1 vccd1 vccd1 _18170_/Y
+ sky130_fd_sc_hd__nand4_2
X_11614_ _11610_/C _11773_/C _11604_/X vssd1 vssd1 vccd1 vccd1 _12167_/A sky130_fd_sc_hd__a21boi_4
X_15382_ _15382_/A _15382_/B _15382_/C vssd1 vssd1 vccd1 vccd1 _15383_/C sky130_fd_sc_hd__and3_1
XFILLER_196_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12688_/B vssd1 vssd1 vccd1 vccd1 _12601_/C sky130_fd_sc_hd__buf_2
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ _17121_/A vssd1 vssd1 vccd1 vccd1 _17334_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14333_ _13994_/A _13994_/B _14135_/A vssd1 vssd1 vccd1 vccd1 _14333_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17052_ _16447_/Y _17975_/A _17744_/A _16523_/C vssd1 vssd1 vccd1 vccd1 _17052_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_100_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14264_ _14340_/B _14260_/Y _13914_/A _14263_/Y vssd1 vssd1 vccd1 vccd1 _14290_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_167_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16003_ _16003_/A vssd1 vssd1 vccd1 vccd1 _16268_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13215_ _13224_/B vssd1 vssd1 vccd1 vccd1 _13523_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14195_ _23360_/Q vssd1 vssd1 vccd1 vccd1 _14878_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ _13196_/C _13146_/B vssd1 vssd1 vccd1 vccd1 _13147_/C sky130_fd_sc_hd__nand2_1
XFILLER_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14658__A1 _21852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14658__B2 _20902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15855__B1 _14569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17954_ _18149_/D _18144_/B _17954_/C vssd1 vssd1 vccd1 vccd1 _17955_/B sky130_fd_sc_hd__and3_1
X_13077_ _13077_/A _13077_/B _13078_/A _13078_/B vssd1 vssd1 vccd1 vccd1 _13077_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21928__B1 _22548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16905_ _16902_/Y _17140_/A _16904_/Y vssd1 vssd1 vccd1 vccd1 _16913_/A sky130_fd_sc_hd__o21ai_1
X_12028_ _12022_/A _12025_/X _12011_/A vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__o21ai_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22050__C1 _22479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17885_ _17885_/A vssd1 vssd1 vccd1 vccd1 _18079_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19624_ _19638_/A _19627_/B _19638_/B _19638_/C vssd1 vssd1 vccd1 vccd1 _19625_/D
+ sky130_fd_sc_hd__nand4_2
X_16836_ _16836_/A _16836_/B vssd1 vssd1 vccd1 vccd1 _16845_/A sky130_fd_sc_hd__nand2_1
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15083__A1 _15356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15083__B2 _15017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19555_ _19534_/D _19532_/X _19554_/X vssd1 vssd1 vccd1 vccd1 _19555_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11890__B _19363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18376__D _18376_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ _16763_/X _16764_/Y _16766_/Y vssd1 vssd1 vccd1 vccd1 _17011_/A sky130_fd_sc_hd__o21ai_2
XFILLER_20_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13979_ _13984_/A vssd1 vssd1 vccd1 vccd1 _14246_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13633__A2 _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18506_ _18506_/A vssd1 vssd1 vccd1 vccd1 _19847_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__13163__A _21054_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15718_ _15718_/A _15798_/A _15799_/A vssd1 vssd1 vccd1 vccd1 _15719_/B sky130_fd_sc_hd__and3_1
X_19486_ _19486_/A _19486_/B vssd1 vssd1 vccd1 vccd1 _19486_/Y sky130_fd_sc_hd__nand2_1
X_16698_ _16939_/A _16939_/B _16706_/A _16706_/B vssd1 vssd1 vccd1 vccd1 _16699_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_55_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22476__A _22476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18437_ _12542_/Y _18571_/A _18571_/B _18437_/D vssd1 vssd1 vccd1 vccd1 _18576_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ _15639_/A _16668_/C _15639_/C _16044_/A vssd1 vssd1 vccd1 vccd1 _15928_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22105__B1 _22102_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_484 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19506__D1 _19502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18368_ _18264_/B _18319_/Y _18370_/B _18405_/A _18367_/Y vssd1 vssd1 vccd1 vccd1
+ _18371_/A sky130_fd_sc_hd__o221a_1
X_17319_ _17314_/X _17315_/X _17316_/Y _17318_/Y vssd1 vssd1 vccd1 vccd1 _17326_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__15138__A2 _13972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18299_ _18295_/X _18296_/X _18298_/X _18245_/C vssd1 vssd1 vccd1 vccd1 _18301_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_175_854 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20330_ _20330_/A _20330_/B _20376_/B vssd1 vssd1 vccd1 vccd1 _20331_/B sky130_fd_sc_hd__or3_2
XFILLER_135_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20261_ _20261_/A _20261_/B vssd1 vssd1 vccd1 vccd1 _23532_/D sky130_fd_sc_hd__xnor2_1
XFILLER_143_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14722__A _23595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22000_ _21884_/B _21996_/Y _21998_/Y vssd1 vssd1 vccd1 vccd1 _22000_/Y sky130_fd_sc_hd__o21ai_1
X_20192_ _20247_/B vssd1 vssd1 vccd1 vccd1 _20252_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15846__B1 _15991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13338__A _13377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14113__A3 _15231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__C _11784_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22902_ _22902_/A vssd1 vssd1 vccd1 vccd1 _23287_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22833_ _22830_/B _22759_/A _22861_/B _22861_/C _22861_/A vssd1 vssd1 vccd1 vccd1
+ _22834_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_112_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11635__A1 _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22764_ _22764_/A _22764_/B _22764_/C vssd1 vssd1 vccd1 vccd1 _22829_/A sky130_fd_sc_hd__nand3_2
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21715_ _21715_/A _21715_/B vssd1 vssd1 vccd1 vccd1 _21723_/C sky130_fd_sc_hd__nor2_1
XFILLER_13_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22695_ _22695_/A _22695_/B vssd1 vssd1 vccd1 vccd1 _23568_/D sky130_fd_sc_hd__nor2_4
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21646_ _21646_/A _21646_/B vssd1 vssd1 vccd1 vccd1 _21649_/C sky130_fd_sc_hd__or2_1
XFILLER_36_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21577_ _21577_/A _21577_/B _21577_/C vssd1 vssd1 vccd1 vccd1 _21614_/B sky130_fd_sc_hd__nand3_1
XFILLER_177_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14337__B1 _15075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23316_ _23381_/CLK _23316_/D vssd1 vssd1 vccd1 vccd1 _23316_/Q sky130_fd_sc_hd__dfxtp_1
X_20528_ _20528_/A _20528_/B _20528_/C vssd1 vssd1 vccd1 vccd1 _20529_/B sky130_fd_sc_hd__nand3_2
XFILLER_181_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20459_ _20464_/B _20464_/C vssd1 vssd1 vccd1 vccd1 _20459_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23247_ _23247_/A vssd1 vssd1 vccd1 vccd1 _23441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13000_ _12864_/A _12864_/B _12851_/Y vssd1 vssd1 vccd1 vccd1 _13001_/A sky130_fd_sc_hd__a21oi_2
XFILLER_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23178_ _23411_/Q input28/X _23178_/S vssd1 vssd1 vccd1 vccd1 _23179_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22129_ _22123_/Y _22126_/X _22264_/B _22647_/A _22128_/Y vssd1 vssd1 vccd1 vccd1
+ _22130_/D sky130_fd_sc_hd__o2111ai_1
XANTENNA__17943__A _17943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input35_A wb_dat_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14951_ _14855_/A _14855_/B _14822_/A vssd1 vssd1 vccd1 vccd1 _14951_/X sky130_fd_sc_hd__o21a_1
XFILLER_153_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13902_ _14068_/A vssd1 vssd1 vccd1 vccd1 _14795_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17670_ _17670_/A _17670_/B _17670_/C vssd1 vssd1 vccd1 vccd1 _17670_/Y sky130_fd_sc_hd__nand3_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14882_ _14883_/A _14883_/B _14883_/C vssd1 vssd1 vccd1 vccd1 _15459_/B sky130_fd_sc_hd__a21oi_2
XFILLER_48_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16621_ _16621_/A _23595_/Q _16808_/A vssd1 vssd1 vccd1 vccd1 _17250_/A sky130_fd_sc_hd__nor3_4
XFILLER_75_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13833_ _13819_/A _13819_/B _13799_/X _13813_/X vssd1 vssd1 vccd1 vccd1 _13834_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13076__B1 _12902_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19340_ _19340_/A vssd1 vssd1 vccd1 vccd1 _19345_/A sky130_fd_sc_hd__clkbuf_1
X_16552_ _16054_/X _16055_/X _16544_/B _16510_/C _16529_/A vssd1 vssd1 vccd1 vccd1
+ _16552_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13764_ _13766_/A _13766_/B _23477_/Q _21882_/B vssd1 vssd1 vccd1 vccd1 _13765_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_188_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22296__A _22476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15503_ _15503_/A _15503_/B vssd1 vssd1 vccd1 vccd1 _15527_/B sky130_fd_sc_hd__xor2_4
XFILLER_31_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19271_ _19263_/X _19261_/X _19297_/B _19297_/A vssd1 vssd1 vccd1 vccd1 _19272_/C
+ sky130_fd_sc_hd__o211ai_1
X_12715_ _12644_/X _12711_/Y _12714_/X vssd1 vssd1 vccd1 vccd1 _12980_/A sky130_fd_sc_hd__a21oi_4
X_16483_ _16483_/A _16483_/B vssd1 vssd1 vccd1 vccd1 _16483_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16294__A _16294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13695_ _13550_/Y _13594_/Y _13694_/Y vssd1 vssd1 vccd1 vccd1 _13763_/A sky130_fd_sc_hd__a21oi_2
XFILLER_31_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18222_ _18279_/D _18279_/A _20265_/C _18330_/A vssd1 vssd1 vccd1 vccd1 _18222_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15434_ _15432_/Y _15434_/B vssd1 vssd1 vccd1 vccd1 _15438_/A sky130_fd_sc_hd__and2b_1
XANTENNA__22638__A1 _13547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12646_ _20675_/A vssd1 vssd1 vccd1 vccd1 _12724_/A sky130_fd_sc_hd__buf_2
XFILLER_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18153_ _23531_/Q _18141_/C _18141_/A _18262_/A _18262_/C vssd1 vssd1 vccd1 vccd1
+ _18206_/A sky130_fd_sc_hd__a32o_1
X_15365_ _14097_/X _14999_/Y _15366_/C _15366_/D _15366_/B vssd1 vssd1 vccd1 vccd1
+ _15365_/X sky130_fd_sc_hd__o32a_1
XFILLER_184_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12577_ _12577_/A vssd1 vssd1 vccd1 vccd1 _13019_/C sky130_fd_sc_hd__buf_2
XFILLER_141_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17104_ _17104_/A _17104_/B vssd1 vssd1 vccd1 vccd1 _17106_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14316_ _23500_/Q vssd1 vssd1 vccd1 vccd1 _14407_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18084_ _18084_/A _18084_/B vssd1 vssd1 vccd1 vccd1 _18110_/B sky130_fd_sc_hd__xor2_1
XFILLER_117_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15296_ _15260_/X _15261_/X _15259_/Y vssd1 vssd1 vccd1 vccd1 _15298_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__20664__A3 _12640_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17035_ _17326_/D _18277_/D _17035_/C _18157_/C vssd1 vssd1 vccd1 vccd1 _17035_/X
+ sky130_fd_sc_hd__and4_2
X_14247_ _14282_/C vssd1 vssd1 vccd1 vccd1 _14347_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_879 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14178_ _14178_/A _14178_/B vssd1 vssd1 vccd1 vccd1 _14178_/Y sky130_fd_sc_hd__nand2_2
XFILLER_113_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13129_ _13136_/B _13136_/C _13136_/A vssd1 vssd1 vccd1 vccd1 _13129_/X sky130_fd_sc_hd__a21o_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _12051_/A _18980_/A _18984_/Y _18985_/X vssd1 vssd1 vccd1 vccd1 _19186_/A
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__12106__A2 _11875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater103 _23481_/Q vssd1 vssd1 vccd1 vccd1 _21987_/B sky130_fd_sc_hd__buf_2
X_17937_ _18256_/A vssd1 vssd1 vccd1 vccd1 _18140_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater114 _23424_/CLK vssd1 vssd1 vccd1 vccd1 _23427_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16469__A _16469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater125 _23444_/CLK vssd1 vssd1 vccd1 vccd1 _23349_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater136 _23402_/CLK vssd1 vssd1 vccd1 vccd1 _23352_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater147 _23307_/CLK vssd1 vssd1 vccd1 vccd1 _23339_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17868_ _17880_/C _17999_/A _17867_/Y vssd1 vssd1 vccd1 vccd1 _17868_/Y sky130_fd_sc_hd__a21oi_2
Xrepeater158 input5/X vssd1 vssd1 vccd1 vccd1 _23321_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15056__A1 _15408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19607_ _19601_/A _19601_/B _19755_/A _19600_/Y vssd1 vssd1 vccd1 vccd1 _19607_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__23452__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16819_ _16819_/A vssd1 vssd1 vccd1 vccd1 _16819_/X sky130_fd_sc_hd__buf_2
X_17799_ _17919_/A _17798_/C _17798_/A vssd1 vssd1 vccd1 vccd1 _17799_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_198_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19538_ _12282_/X _12283_/Y _19709_/B _19709_/C vssd1 vssd1 vccd1 vccd1 _19538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22637__C _22637_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19469_ _19389_/A _19389_/B _19389_/C _19601_/B _19601_/A vssd1 vssd1 vccd1 vccd1
+ _19755_/B sky130_fd_sc_hd__a32o_1
XANTENNA__12290__A1 _12090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21500_ _21500_/A _21548_/B _21546_/A _21548_/D vssd1 vssd1 vccd1 vccd1 _21502_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22480_ _22477_/Y _22479_/Y _22476_/X vssd1 vssd1 vccd1 vccd1 _22480_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_107_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19011__C _19700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21431_ _21431_/A _21431_/B _21431_/C vssd1 vssd1 vccd1 vccd1 _21431_/X sky130_fd_sc_hd__and3_1
XANTENNA__12042__A1 _18481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12237__A _12237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16859__A2 _17465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21362_ _21292_/Y _21433_/A _21314_/A _21359_/Y _21455_/A vssd1 vssd1 vccd1 vccd1
+ _21453_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20313_ _20313_/A _20313_/B vssd1 vssd1 vccd1 vccd1 _23533_/D sky130_fd_sc_hd__xor2_1
X_23101_ _23101_/A vssd1 vssd1 vccd1 vccd1 _23376_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__23054__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21293_ _21545_/A _20471_/Y _21292_/Y vssd1 vssd1 vccd1 vccd1 _21293_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_174_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14452__A _15208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23032_ _23346_/Q input27/X _23034_/S vssd1 vssd1 vccd1 vccd1 _23033_/A sky130_fd_sc_hd__mux2_1
X_20244_ _20244_/A _20243_/Y vssd1 vssd1 vccd1 vccd1 _20252_/C sky130_fd_sc_hd__or2b_1
XANTENNA__18859__A _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16087__A3 _17414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20175_ _20175_/A _20283_/B _20175_/C vssd1 vssd1 vccd1 vccd1 _20176_/C sky130_fd_sc_hd__nand3_2
XANTENNA__21080__A3 _20953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14098__A2 _14184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15295__A1 _14588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11856__A1 _12378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11856__B2 _14729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22816_ _23282_/Q _22817_/B vssd1 vssd1 vccd1 vccd1 _22856_/C sky130_fd_sc_hd__nand2_1
XFILLER_60_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18536__A2 _11611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22747_ _22747_/A _22747_/B vssd1 vssd1 vccd1 vccd1 _23569_/D sky130_fd_sc_hd__xor2_4
XFILLER_73_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12500_ _23593_/Q vssd1 vssd1 vccd1 vccd1 _16620_/C sky130_fd_sc_hd__inv_2
XFILLER_198_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13480_ _13600_/C vssd1 vssd1 vccd1 vccd1 _22159_/C sky130_fd_sc_hd__buf_2
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22678_ _22756_/C _22548_/A _22548_/C _22677_/Y vssd1 vssd1 vccd1 vccd1 _22678_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12431_ _12052_/A _19190_/A _12441_/A vssd1 vssd1 vccd1 vccd1 _12438_/A sky130_fd_sc_hd__o21ai_1
X_21629_ _21660_/C _21660_/A vssd1 vssd1 vccd1 vccd1 _23551_/D sky130_fd_sc_hd__xor2_1
XFILLER_138_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15770__A2 _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13781__A1 _13453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15150_ _15140_/B _15138_/X _15140_/C vssd1 vssd1 vccd1 vccd1 _15214_/B sky130_fd_sc_hd__a21bo_1
X_12362_ _12186_/Y _12327_/Y _12336_/A _12360_/Y _12329_/X vssd1 vssd1 vccd1 vccd1
+ _12363_/D sky130_fd_sc_hd__o2111ai_2
XFILLER_193_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_846 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14101_ _14791_/C _14777_/B vssd1 vssd1 vccd1 vccd1 _14101_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23045__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12293_ _12297_/A vssd1 vssd1 vccd1 vccd1 _12293_/Y sky130_fd_sc_hd__inv_2
X_15081_ _15081_/A _15081_/B vssd1 vssd1 vccd1 vccd1 _15093_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14032_ _14017_/X _13946_/A _14031_/X vssd1 vssd1 vccd1 vccd1 _14312_/B sky130_fd_sc_hd__a21o_2
XFILLER_134_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_890 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18472__A1 _11848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18840_ _18830_/Y _18833_/Y _18839_/Y vssd1 vssd1 vccd1 vccd1 _18840_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_80_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18472__B2 _18490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18771_ _18771_/A vssd1 vssd1 vccd1 vccd1 _18969_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15983_ _15983_/A vssd1 vssd1 vccd1 vccd1 _16840_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16289__A _17226_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17722_ _17722_/A vssd1 vssd1 vccd1 vccd1 _17723_/B sky130_fd_sc_hd__buf_2
XANTENNA__13706__A _22159_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14934_ _14934_/A _14934_/B _14934_/C _14934_/D vssd1 vssd1 vccd1 vccd1 _14934_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__15038__A1 _15208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18775__A2 _18966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17653_ _17653_/A _17653_/B _17653_/C vssd1 vssd1 vccd1 vccd1 _17666_/A sky130_fd_sc_hd__nand3_2
XANTENNA__16924__A1_N _16935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14865_ _14865_/A vssd1 vssd1 vccd1 vccd1 _14970_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__13425__B _13810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16604_ _16604_/A vssd1 vssd1 vccd1 vccd1 _16604_/X sky130_fd_sc_hd__clkbuf_4
X_13816_ _13816_/A _21764_/B _23475_/Q _21919_/C vssd1 vssd1 vccd1 vccd1 _13818_/B
+ sky130_fd_sc_hd__nand4_4
X_17584_ _16356_/A _17565_/X _17566_/X _17575_/X _17571_/Y vssd1 vssd1 vccd1 vccd1
+ _17585_/C sky130_fd_sc_hd__o221ai_4
XFILLER_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14796_ _14796_/A _14796_/B _15195_/C vssd1 vssd1 vccd1 vccd1 _14796_/Y sky130_fd_sc_hd__nand3_1
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ _19323_/A _20046_/A _20047_/A vssd1 vssd1 vccd1 vccd1 _19491_/B sky130_fd_sc_hd__nand3_4
X_16535_ _16519_/Y _16522_/Y _16564_/A _16534_/Y vssd1 vssd1 vccd1 vccd1 _16562_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13747_ _13748_/C _13748_/B _13715_/X vssd1 vssd1 vccd1 vccd1 _13747_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__17735__B1 _17567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19254_ _19254_/A vssd1 vssd1 vccd1 vccd1 _19254_/Y sky130_fd_sc_hd__inv_2
X_16466_ _16463_/Y _16465_/Y _16507_/A _16441_/Y vssd1 vssd1 vccd1 vccd1 _16467_/C
+ sky130_fd_sc_hd__a22oi_2
X_13678_ _13672_/X _13674_/X _13671_/A _13671_/B vssd1 vssd1 vccd1 vccd1 _13682_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__22754__A _22754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18205_ _18199_/Y _18200_/X _18263_/A vssd1 vssd1 vccd1 vccd1 _18262_/B sky130_fd_sc_hd__o21a_1
X_15417_ _15446_/D _15446_/C _15485_/D _15511_/D _15366_/D vssd1 vssd1 vccd1 vccd1
+ _15424_/A sky130_fd_sc_hd__a41o_1
X_19185_ _16360_/X _18971_/X _19858_/A _18975_/X _18978_/B vssd1 vssd1 vccd1 vccd1
+ _19185_/X sky130_fd_sc_hd__o311a_1
X_12629_ _13052_/A _21035_/C _13052_/C vssd1 vssd1 vccd1 vccd1 _12654_/A sky130_fd_sc_hd__nand3_4
X_16397_ _16397_/A _16397_/B vssd1 vssd1 vccd1 vccd1 _16407_/A sky130_fd_sc_hd__nand2_1
XFILLER_191_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18136_ _18136_/A _18136_/B vssd1 vssd1 vccd1 vccd1 _18252_/A sky130_fd_sc_hd__nand2_1
X_15348_ _15348_/A vssd1 vssd1 vccd1 vccd1 _15348_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18067_ _18067_/A _18067_/B vssd1 vssd1 vccd1 vccd1 _18068_/A sky130_fd_sc_hd__or2_1
XFILLER_145_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23036__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15279_ _15279_/A _15279_/B vssd1 vssd1 vccd1 vccd1 _15292_/B sky130_fd_sc_hd__nand2_2
XFILLER_160_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17018_ _17018_/A _17018_/B vssd1 vssd1 vccd1 vccd1 _17019_/C sky130_fd_sc_hd__nand2_1
XFILLER_171_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18463__A1 _12052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21062__A3 _12640_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20270__A1 _18211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _18969_/A _18969_/B _18969_/C _18969_/D vssd1 vssd1 vccd1 vccd1 _19059_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21980_ _21980_/A vssd1 vssd1 vccd1 vccd1 _22617_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20931_ _20919_/Y _20926_/Y _20941_/B _20941_/A vssd1 vssd1 vccd1 vccd1 _20947_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20862_ _20862_/A _20862_/B vssd1 vssd1 vccd1 vccd1 _20885_/B sky130_fd_sc_hd__nor2_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23470__D _23482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22601_ _22830_/B _22126_/X _22506_/X vssd1 vssd1 vccd1 vccd1 _22601_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23581_ _23582_/CLK _23581_/D vssd1 vssd1 vccd1 vccd1 _23581_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12263__B2 _11898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20793_ _20793_/A _20793_/B vssd1 vssd1 vccd1 vccd1 _20794_/C sky130_fd_sc_hd__nand2_1
XFILLER_195_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16365__C _18481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22532_ _22532_/A _23277_/Q vssd1 vssd1 vccd1 vccd1 _22532_/Y sky130_fd_sc_hd__nand2_1
XFILLER_195_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_774 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19479__B1 _18503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22463_ _22463_/A _22463_/B _22463_/C vssd1 vssd1 vccd1 vccd1 _22475_/B sky130_fd_sc_hd__nand3_1
XFILLER_176_960 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21414_ _21414_/A vssd1 vssd1 vccd1 vccd1 _21616_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1024 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22394_ _22463_/C _22394_/B _22394_/C vssd1 vssd1 vccd1 vccd1 _22394_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_185_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21345_ _21345_/A _21345_/B _21345_/C vssd1 vssd1 vccd1 vccd1 _21346_/A sky130_fd_sc_hd__nand3_1
XFILLER_68_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12117__D _18849_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15504__A2 _15527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21276_ _21276_/A vssd1 vssd1 vccd1 vccd1 _21448_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__20912__A _21174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20227_ _20156_/Y _20153_/Y _20224_/Y _20225_/X _20158_/B vssd1 vssd1 vccd1 vccd1
+ _20283_/A sky130_fd_sc_hd__o221a_1
X_23015_ _23338_/Q input19/X _23023_/S vssd1 vssd1 vccd1 vccd1 _23016_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16465__B1 _12238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20158_ _20158_/A _20158_/B _20158_/C _20158_/D vssd1 vssd1 vccd1 vccd1 _20159_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20089_ _20070_/Y _20172_/A _20074_/X vssd1 vssd1 vccd1 vccd1 _20090_/B sky130_fd_sc_hd__a21oi_1
XFILLER_76_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12980_ _12980_/A vssd1 vssd1 vccd1 vccd1 _12981_/C sky130_fd_sc_hd__buf_2
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14491__A2 _15446_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _11931_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_855 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18755__C _18755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _15645_/A vssd1 vssd1 vccd1 vccd1 _16657_/B sky130_fd_sc_hd__clkbuf_4
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11862_ _11861_/A _11608_/A _12245_/A vssd1 vssd1 vccd1 vccd1 _11887_/A sky130_fd_sc_hd__a21o_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18509__A2 _11926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19706__B2 _18003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13601_ _13783_/B _13783_/C vssd1 vssd1 vccd1 vccd1 _13602_/A sky130_fd_sc_hd__nand2_2
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14581_ _23420_/Q vssd1 vssd1 vccd1 vccd1 _15664_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11793_ _11886_/A vssd1 vssd1 vccd1 vccd1 _18973_/C sky130_fd_sc_hd__buf_2
X_16320_ _16355_/A _16384_/A _16458_/A _16382_/A _16316_/Y vssd1 vssd1 vccd1 vccd1
+ _16321_/B sky130_fd_sc_hd__o221ai_1
XANTENNA__13261__A _23333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13532_ _13502_/X _13736_/B _13527_/X _13531_/X vssd1 vssd1 vccd1 vccd1 _13545_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_595 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16251_ _16251_/A _16251_/B _16281_/B _16251_/D vssd1 vssd1 vccd1 vccd1 _16251_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13463_ _13463_/A vssd1 vssd1 vccd1 vccd1 _13517_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15202_ _15277_/A _15203_/B _15203_/A vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__a21o_1
XFILLER_51_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12414_ _12241_/A _18461_/B _18460_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _12455_/C
+ sky130_fd_sc_hd__o31ai_2
X_16182_ _19161_/A _15936_/A _17137_/C _16113_/A _12306_/A vssd1 vssd1 vccd1 vccd1
+ _16183_/A sky130_fd_sc_hd__a32oi_4
XFILLER_139_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13394_ _13394_/A _13394_/B vssd1 vssd1 vccd1 vccd1 _13394_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18142__B1 _23531_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15133_ _15132_/A _15132_/B _15132_/C vssd1 vssd1 vccd1 vccd1 _15134_/C sky130_fd_sc_hd__a21o_1
X_12345_ _18778_/C vssd1 vssd1 vccd1 vccd1 _19261_/C sky130_fd_sc_hd__buf_4
XFILLER_5_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12309__A2 _16364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13506__A1 _22553_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19941_ _19655_/X _19855_/C _19871_/X _19688_/B _19867_/A vssd1 vssd1 vccd1 vccd1
+ _19941_/X sky130_fd_sc_hd__o311a_1
X_15064_ _15064_/A _15064_/B vssd1 vssd1 vccd1 vccd1 _15064_/X sky130_fd_sc_hd__xor2_2
X_12276_ _11766_/C _11760_/A _11885_/Y _11880_/X _11803_/X vssd1 vssd1 vccd1 vccd1
+ _12276_/X sky130_fd_sc_hd__o311a_1
XFILLER_175_94 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14015_ _14588_/A _14015_/B _14015_/C vssd1 vssd1 vccd1 vccd1 _14120_/A sky130_fd_sc_hd__nand3b_2
XFILLER_49_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19872_ _19870_/X _19871_/X _19688_/B vssd1 vssd1 vccd1 vccd1 _19873_/A sky130_fd_sc_hd__o21ai_1
XFILLER_150_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18823_ _19019_/C vssd1 vssd1 vccd1 vccd1 _19539_/B sky130_fd_sc_hd__buf_2
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18754_ _18537_/Y _18932_/A _18602_/Y vssd1 vssd1 vccd1 vccd1 _18754_/Y sky130_fd_sc_hd__a21oi_1
X_15966_ _16119_/A _16153_/A _16132_/A vssd1 vssd1 vccd1 vccd1 _15998_/B sky130_fd_sc_hd__o21ai_4
XFILLER_95_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17705_ _17705_/A _17705_/B vssd1 vssd1 vccd1 vccd1 _17705_/Y sky130_fd_sc_hd__nand2_1
X_14917_ _14918_/C _14918_/B _14918_/A vssd1 vssd1 vccd1 vccd1 _14926_/B sky130_fd_sc_hd__a21o_1
XFILLER_64_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18685_ _18677_/Y _18678_/Y _18684_/X vssd1 vssd1 vccd1 vccd1 _18687_/B sky130_fd_sc_hd__a21o_1
XFILLER_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15897_ _16078_/A _16078_/B _16078_/C _15896_/X vssd1 vssd1 vccd1 vccd1 _16008_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19123__A _19703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17636_ _16408_/X _18002_/A _17410_/Y _17625_/Y _17629_/Y vssd1 vssd1 vccd1 vccd1
+ _17637_/C sky130_fd_sc_hd__o221ai_1
XFILLER_1_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14848_ _14846_/Y _14847_/Y _15065_/A _14853_/B vssd1 vssd1 vccd1 vccd1 _14848_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17567_ _18947_/A vssd1 vssd1 vccd1 vccd1 _17567_/X sky130_fd_sc_hd__buf_2
XFILLER_1_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14779_ _15085_/B _15085_/C _14246_/B vssd1 vssd1 vccd1 vccd1 _14779_/X sky130_fd_sc_hd__or3b_1
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19306_ _19158_/A _19304_/A _19305_/Y vssd1 vssd1 vccd1 vccd1 _19306_/X sky130_fd_sc_hd__a21o_1
X_16518_ _16518_/A _16518_/B _16518_/C vssd1 vssd1 vccd1 vccd1 _16518_/Y sky130_fd_sc_hd__nand3_1
XFILLER_56_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19173__A2 _11713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_584 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ _17498_/A _17498_/B _17498_/C vssd1 vssd1 vccd1 vccd1 _17502_/B sky130_fd_sc_hd__nand3_1
XFILLER_108_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22484__A _22484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19237_ _19147_/A _19147_/B _19256_/B _19226_/A vssd1 vssd1 vccd1 vccd1 _19244_/A
+ sky130_fd_sc_hd__a22o_1
X_16449_ _16389_/X _16523_/D _16364_/X _16438_/Y vssd1 vssd1 vccd1 vccd1 _16449_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16931__A1 _16066_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19168_ _19168_/A vssd1 vssd1 vccd1 vccd1 _19325_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18119_ _18119_/A _18245_/A vssd1 vssd1 vccd1 vccd1 _18123_/C sky130_fd_sc_hd__nand2_1
XANTENNA__17728__D _19957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19099_ _19101_/B _19101_/C _23543_/Q vssd1 vssd1 vccd1 vccd1 _19100_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__21283__A3 _21432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18684__B2 _11961_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21130_ _21130_/A vssd1 vssd1 vccd1 vccd1 _21131_/A sky130_fd_sc_hd__inv_2
XANTENNA__16695__B1 _16706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14433__C _14867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21828__A _22420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21061_ _21061_/A vssd1 vssd1 vccd1 vccd1 _21061_/X sky130_fd_sc_hd__buf_2
XFILLER_87_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20012_ _20012_/A _20012_/B _20012_/C vssd1 vssd1 vccd1 vccd1 _20108_/A sky130_fd_sc_hd__nand3_1
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23465__D _23477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19017__B _19703_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21991__A1 _21829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13346__A _23325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23193__A0 _15762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14473__A2 _14933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15670__A1 _12373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23254__S _23254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21963_ _21964_/A _21964_/B _21964_/C vssd1 vssd1 vccd1 vccd1 _21965_/B sky130_fd_sc_hd__a21o_1
XFILLER_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ _21370_/A _21172_/A _21369_/A vssd1 vssd1 vccd1 vccd1 _20914_/Y sky130_fd_sc_hd__nand3_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21894_ _21891_/Y _13553_/X _21892_/X _21798_/C _21893_/Y vssd1 vssd1 vccd1 vccd1
+ _21894_/X sky130_fd_sc_hd__o311a_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16376__B _17062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ _20845_/A vssd1 vssd1 vccd1 vccd1 _20847_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15973__A2 _15856_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23564_ _23566_/CLK _23564_/D vssd1 vssd1 vccd1 vccd1 _23564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20776_ _20776_/A vssd1 vssd1 vccd1 vccd1 _21000_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23248__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22515_ _22516_/A _22516_/B _22516_/C _22516_/D vssd1 vssd1 vccd1 vccd1 _22609_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23495_ _23499_/CLK _23507_/Q vssd1 vssd1 vccd1 vccd1 _23495_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_195_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22446_ _22445_/Y _22617_/A _22443_/Y vssd1 vssd1 vccd1 vccd1 _22447_/B sky130_fd_sc_hd__a21oi_1
XFILLER_148_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22377_ _22377_/A vssd1 vssd1 vccd1 vccd1 _22461_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__22471__A2 _22754_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ _12130_/A vssd1 vssd1 vccd1 vccd1 _12130_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_150_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21328_ _21319_/A _21319_/B _21308_/Y _21309_/X vssd1 vssd1 vccd1 vccd1 _21328_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_123_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21259_ _23564_/Q _21144_/B _21258_/Y vssd1 vssd1 vccd1 vccd1 _21259_/X sky130_fd_sc_hd__o21a_1
XANTENNA__15736__A _15736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ _11906_/Y _11914_/X _12064_/B _12064_/C vssd1 vssd1 vccd1 vccd1 _12061_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__22223__A2 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14640__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15820_ _15813_/A _15709_/A _15785_/A _17259_/A _16462_/B vssd1 vssd1 vccd1 vccd1
+ _16020_/B sky130_fd_sc_hd__o2111ai_4
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _11853_/A _11921_/Y _15736_/A _15738_/A _15841_/B vssd1 vssd1 vccd1 vccd1
+ _15753_/A sky130_fd_sc_hd__o221ai_2
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12963_ _13119_/A vssd1 vssd1 vccd1 vccd1 _20563_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _23407_/Q _14693_/X _14698_/X _23439_/Q _14701_/X vssd1 vssd1 vccd1 vccd1
+ _14702_/X sky130_fd_sc_hd__a221o_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _12391_/B _12251_/B _12253_/A vssd1 vssd1 vccd1 vccd1 _11914_/X sky130_fd_sc_hd__o21a_1
XANTENNA__21192__B _21493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18470_ _18470_/A _18997_/B _18470_/C vssd1 vssd1 vccd1 vccd1 _18478_/A sky130_fd_sc_hd__nand3_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15682_ _15682_/A _15682_/B _15974_/C _15682_/D vssd1 vssd1 vccd1 vccd1 _15682_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12894_ _12899_/A _12894_/B _12894_/C vssd1 vssd1 vccd1 vccd1 _12894_/X sky130_fd_sc_hd__and3_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17421_ _12237_/A _16741_/A _17411_/Y _17420_/Y vssd1 vssd1 vccd1 vccd1 _17426_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _14633_/A _14633_/B _14633_/C _14519_/D vssd1 vssd1 vccd1 vccd1 _14688_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_61_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11845_ _12353_/A _11822_/X _11837_/Y _11844_/Y vssd1 vssd1 vccd1 vccd1 _11912_/A
+ sky130_fd_sc_hd__o22ai_4
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_730 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17352_ _17358_/B vssd1 vssd1 vccd1 vccd1 _17514_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ input46/X _14518_/X _14563_/X vssd1 vssd1 vccd1 vccd1 _14564_/X sky130_fd_sc_hd__a21o_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _11738_/X _11740_/X _11741_/Y _11747_/X _11749_/X vssd1 vssd1 vccd1 vccd1
+ _11788_/A sky130_fd_sc_hd__o2111a_2
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _15862_/A _15862_/B _15682_/A vssd1 vssd1 vccd1 vccd1 _16303_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13515_ _13519_/A _13515_/B _13515_/C vssd1 vssd1 vccd1 vccd1 _13537_/A sky130_fd_sc_hd__nand3b_1
X_17283_ _20049_/A vssd1 vssd1 vccd1 vccd1 _17960_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23239__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14495_ _14495_/A _14495_/B _14495_/C _14495_/D vssd1 vssd1 vccd1 vccd1 _14497_/B
+ sky130_fd_sc_hd__nand4_1
X_19022_ _19018_/X _19020_/Y _19021_/X vssd1 vssd1 vccd1 vccd1 _19026_/A sky130_fd_sc_hd__a21o_1
X_16234_ _16234_/A _16234_/B _16234_/C vssd1 vssd1 vccd1 vccd1 _16242_/B sky130_fd_sc_hd__nand3_2
X_13446_ _13446_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13447_/C sky130_fd_sc_hd__nand2_1
XFILLER_70_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1030 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16165_ _16165_/A vssd1 vssd1 vccd1 vccd1 _19381_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_86_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13377_ _13377_/A _13377_/B _13377_/C _13377_/D vssd1 vssd1 vccd1 vccd1 _13785_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_155_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15116_ _15254_/A _15116_/B _15254_/C vssd1 vssd1 vccd1 vccd1 _15257_/B sky130_fd_sc_hd__and3_1
XFILLER_170_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12328_ _19180_/C vssd1 vssd1 vccd1 vccd1 _19512_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_114_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17845__B _19799_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16096_ _16096_/A vssd1 vssd1 vccd1 vccd1 _16096_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19924_ _19924_/A vssd1 vssd1 vccd1 vccd1 _20205_/A sky130_fd_sc_hd__clkbuf_2
X_15047_ _14945_/B _14945_/C _14931_/Y vssd1 vssd1 vccd1 vccd1 _15049_/B sky130_fd_sc_hd__a21o_1
X_12259_ _18500_/A vssd1 vssd1 vccd1 vccd1 _18673_/A sky130_fd_sc_hd__buf_2
XFILLER_69_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20225__A1 _18001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12989__B _13181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19855_ _19855_/A _19855_/B _19855_/C vssd1 vssd1 vccd1 vccd1 _19943_/B sky130_fd_sc_hd__nand3_2
XFILLER_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18957__A _19123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__B1 _11717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15101__B1 _14632_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13166__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18806_ _18806_/A _18806_/B vssd1 vssd1 vccd1 vccd1 _18808_/B sky130_fd_sc_hd__nand2_2
XFILLER_96_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19786_ _19785_/X _19924_/A _19776_/X _19783_/X vssd1 vssd1 vccd1 vccd1 _19787_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_95_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16998_ _16777_/Y _16998_/B _16998_/C _17376_/A vssd1 vssd1 vccd1 vccd1 _17017_/A
+ sky130_fd_sc_hd__nand4b_1
XFILLER_110_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14455__A2 _15238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18737_ _18738_/B _18738_/C _23541_/Q vssd1 vssd1 vccd1 vccd1 _19288_/A sky130_fd_sc_hd__a21bo_1
X_15949_ _15949_/A vssd1 vssd1 vccd1 vccd1 _15949_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18668_ _18669_/A _18669_/B _18669_/C _18669_/D vssd1 vssd1 vccd1 vccd1 _18868_/A
+ sky130_fd_sc_hd__a22o_2
XANTENNA__14207__A2 _14061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17619_ _17958_/A _16478_/X _17605_/Y _17598_/Y _17607_/X vssd1 vssd1 vccd1 vccd1
+ _17619_/X sky130_fd_sc_hd__o311a_1
XFILLER_24_549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18599_ _18599_/A _18599_/B vssd1 vssd1 vccd1 vccd1 _18599_/Y sky130_fd_sc_hd__nor2_2
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20630_ _20625_/Y _20626_/Y _20627_/Y _20632_/A vssd1 vssd1 vccd1 vccd1 _20631_/A
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__17157__A1 _17154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20561_ _13066_/X _20565_/D _13065_/Y vssd1 vssd1 vccd1 vccd1 _20562_/B sky130_fd_sc_hd__a21oi_2
XFILLER_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22300_ _22300_/A _22300_/B vssd1 vssd1 vccd1 vccd1 _22300_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13718__A1 _21892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23280_ _23518_/CLK _23280_/D vssd1 vssd1 vccd1 vccd1 _23280_/Q sky130_fd_sc_hd__dfxtp_1
X_20492_ _20518_/A _20492_/B vssd1 vssd1 vccd1 vccd1 _20512_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22231_ _22231_/A _22231_/B vssd1 vssd1 vccd1 vccd1 _22234_/B sky130_fd_sc_hd__nand2_1
XFILLER_192_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19854__B1 _19649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22162_ _22162_/A _22162_/B vssd1 vssd1 vccd1 vccd1 _22166_/A sky130_fd_sc_hd__nand2_2
XFILLER_105_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20462__A _20902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21113_ _21113_/A _21113_/B _21113_/C vssd1 vssd1 vccd1 vccd1 _21134_/A sky130_fd_sc_hd__nand3_1
XANTENNA__22380__C _22380_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22093_ _22093_/A _22093_/B _22093_/C _22093_/D vssd1 vssd1 vccd1 vccd1 _22094_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_182_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20216__A1 _18211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15891__A1 _15985_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21044_ _20934_/B _21176_/C _12634_/X _21635_/B _21184_/A vssd1 vssd1 vccd1 vccd1
+ _21045_/C sky130_fd_sc_hd__o221ai_1
XFILLER_160_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19621__A3 _19358_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17093__B1 _17712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23536__CLK _23558_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22995_ _14614_/X input9/X _23001_/S vssd1 vssd1 vccd1 vccd1 _22996_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21946_ _21946_/A _21946_/B _21946_/C vssd1 vssd1 vccd1 vccd1 _21947_/A sky130_fd_sc_hd__nand3_1
XFILLER_55_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12209__A1 _16066_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13523__B _22637_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19698__A _19698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21877_ _21877_/A vssd1 vssd1 vccd1 vccd1 _22263_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11935_/A vssd1 vssd1 vccd1 vccd1 _18675_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20828_ _20828_/A _20828_/B _20828_/C vssd1 vssd1 vccd1 vccd1 _20887_/A sky130_fd_sc_hd__nand3_1
XFILLER_11_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20637__A _23298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23547_ _23578_/CLK _23547_/D vssd1 vssd1 vccd1 vccd1 _23547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19210__B _19649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20759_ _20755_/X _20606_/A _20607_/B _20607_/C vssd1 vssd1 vccd1 vccd1 _20759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_196_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_896 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ _13497_/A vssd1 vssd1 vccd1 vccd1 _13736_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14280_ _14251_/Y _14245_/Y _14282_/C vssd1 vssd1 vccd1 vccd1 _14349_/C sky130_fd_sc_hd__o21bai_1
X_23478_ _23499_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _23478_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13231_ _23333_/Q vssd1 vssd1 vccd1 vccd1 _13339_/A sky130_fd_sc_hd__inv_2
X_22429_ _22428_/A _22428_/B _22402_/A _22428_/D vssd1 vssd1 vccd1 vccd1 _22430_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19845__B1 _17406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17305__D1 _17712_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13162_ _13162_/A _13162_/B vssd1 vssd1 vccd1 vccd1 _13169_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17320__A1 _18211_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12113_ _12403_/A vssd1 vssd1 vccd1 vccd1 _12113_/X sky130_fd_sc_hd__buf_2
X_17970_ _18157_/D _18157_/B _17960_/X vssd1 vssd1 vccd1 vccd1 _17970_/Y sky130_fd_sc_hd__a21oi_1
X_13093_ _23456_/Q vssd1 vssd1 vccd1 vccd1 _20769_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12044_ _18941_/B vssd1 vssd1 vccd1 vccd1 _19381_/D sky130_fd_sc_hd__buf_2
X_16921_ _17133_/A _17133_/B _16921_/C vssd1 vssd1 vccd1 vccd1 _16923_/A sky130_fd_sc_hd__and3_2
XFILLER_120_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1075 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19640_ _19637_/Y _19444_/X _19772_/A vssd1 vssd1 vccd1 vccd1 _19640_/Y sky130_fd_sc_hd__a21oi_2
X_16852_ _16823_/Y _16825_/Y _17073_/B _17073_/A _16836_/B vssd1 vssd1 vccd1 vccd1
+ _16853_/C sky130_fd_sc_hd__o221ai_1
XANTENNA__18820__A1 _19505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15803_ _17465_/A _15800_/Y _15802_/Y vssd1 vssd1 vccd1 vccd1 _15808_/A sky130_fd_sc_hd__o21ai_1
XFILLER_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19571_ _19587_/A _19588_/B _19570_/X vssd1 vssd1 vccd1 vccd1 _19571_/Y sky130_fd_sc_hd__a21oi_1
X_16783_ _16998_/C _16777_/Y _16998_/B _17022_/A vssd1 vssd1 vccd1 vccd1 _16987_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12448__A1 _11822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13995_ _14312_/D vssd1 vssd1 vccd1 vccd1 _14867_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18522_ _18522_/A _18522_/B vssd1 vssd1 vccd1 vccd1 _18529_/B sky130_fd_sc_hd__nand2_1
X_15734_ _16860_/A _17098_/C _16526_/B _15964_/B vssd1 vssd1 vccd1 vccd1 _16070_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12946_ _12933_/X _12943_/X _12944_/Y _12945_/Y vssd1 vssd1 vccd1 vccd1 _13109_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21183__A2 _21592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _23424_/Q _15665_/B vssd1 vssd1 vccd1 vccd1 _16684_/A sky130_fd_sc_hd__nand2_1
X_18453_ _18453_/A vssd1 vssd1 vccd1 vccd1 _18453_/X sky130_fd_sc_hd__buf_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _20906_/A _20907_/A _12696_/A _20908_/A vssd1 vssd1 vccd1 vccd1 _12877_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20930__A2 _21592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _17493_/A _17493_/B _17405_/C vssd1 vssd1 vccd1 vccd1 _17663_/A sky130_fd_sc_hd__a21o_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _23361_/Q vssd1 vssd1 vccd1 vccd1 _14879_/C sky130_fd_sc_hd__buf_4
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18384_ _18384_/A _18384_/B _18343_/B vssd1 vssd1 vccd1 vccd1 _18413_/A sky130_fd_sc_hd__nor3b_1
X_11828_ _11841_/A _11828_/B _12403_/A vssd1 vssd1 vccd1 vccd1 _12118_/C sky130_fd_sc_hd__nand3_1
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15596_ _23416_/Q _23417_/Q vssd1 vssd1 vccd1 vccd1 _15685_/A sky130_fd_sc_hd__nor2_1
XANTENNA__17139__A1 _12004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17335_ _17335_/A _17335_/B vssd1 vssd1 vccd1 vccd1 _17336_/C sky130_fd_sc_hd__nand2_1
XFILLER_14_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14547_ _14547_/A vssd1 vssd1 vccd1 vccd1 _14547_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11759_ _18812_/A _18814_/A _11977_/B vssd1 vssd1 vccd1 vccd1 _11760_/B sky130_fd_sc_hd__a21oi_4
XFILLER_92_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18017__A _18163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17266_ _17260_/A _17260_/B _17265_/Y _17243_/D _20049_/A vssd1 vssd1 vccd1 vccd1
+ _17275_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14478_ _14476_/X _14478_/B _14478_/C vssd1 vssd1 vccd1 vccd1 _14478_/X sky130_fd_sc_hd__and3b_1
XANTENNA__16362__A2 _15884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19005_ _11654_/A _18442_/A _19000_/Y vssd1 vssd1 vccd1 vccd1 _19013_/A sky130_fd_sc_hd__o21ai_1
X_16217_ _16217_/A _16217_/B vssd1 vssd1 vccd1 vccd1 _16217_/Y sky130_fd_sc_hd__nand2_1
X_13429_ _13430_/A _13466_/A _13425_/Y _13444_/A vssd1 vssd1 vccd1 vccd1 _13443_/A
+ sky130_fd_sc_hd__o22a_1
X_17197_ _17035_/X _16923_/A _16917_/X vssd1 vssd1 vccd1 vccd1 _17200_/B sky130_fd_sc_hd__o21ai_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16148_ _17431_/A vssd1 vssd1 vccd1 vccd1 _17565_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_127_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17311__A1 _17140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079_ _15878_/X _15879_/Y _15888_/Y vssd1 vssd1 vccd1 vccd1 _16081_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__23559__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14676__A2 _14672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19907_ _19894_/Y _19899_/Y _19901_/X vssd1 vssd1 vccd1 vccd1 _19909_/B sky130_fd_sc_hd__a21o_1
XFILLER_190_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17591__A _17591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17614__A2 _17285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19838_ _19838_/A vssd1 vssd1 vccd1 vccd1 _20081_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_874 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23148__A0 _18434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16822__B1 _16638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
X_19769_ _19771_/B _19771_/C vssd1 vssd1 vccd1 vccd1 _19769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21800_ _13826_/X _21795_/X _21794_/Y _21799_/X _13818_/B vssd1 vssd1 vccd1 vccd1
+ _21801_/C sky130_fd_sc_hd__o221ai_2
XFILLER_65_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22780_ _22780_/A _22780_/B vssd1 vssd1 vccd1 vccd1 _22780_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21731_ _23578_/Q _21729_/X _21730_/X _21728_/Y vssd1 vssd1 vccd1 vccd1 _23558_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19119__A2 _17593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16935__A _16935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16050__A1 _16372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16050__B2 _16757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21858__A_N _13867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21662_ _21657_/X _21660_/D _21661_/Y vssd1 vssd1 vccd1 vccd1 _21688_/B sky130_fd_sc_hd__a21o_1
X_23401_ _23401_/CLK _23401_/D vssd1 vssd1 vccd1 vccd1 _23401_/Q sky130_fd_sc_hd__dfxtp_1
X_20613_ _20613_/A vssd1 vssd1 vccd1 vccd1 _21415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12611__A1 _12601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21593_ _21428_/X _21637_/C _21592_/B vssd1 vssd1 vccd1 vccd1 _21594_/B sky130_fd_sc_hd__a21boi_1
XFILLER_193_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23332_ _23332_/CLK _23332_/D vssd1 vssd1 vccd1 vccd1 _23332_/Q sky130_fd_sc_hd__dfxtp_1
X_20544_ _20548_/A _20553_/B _20553_/C vssd1 vssd1 vccd1 vccd1 _20552_/A sky130_fd_sc_hd__a21o_1
Xclkbuf_3_1_0_bq_clk_i clkbuf_3_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_165_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17550__A1 _12323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23263_ _23584_/CLK _23263_/D vssd1 vssd1 vccd1 vccd1 _23263_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20475_ _20475_/A _20475_/B vssd1 vssd1 vccd1 vccd1 _20634_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22214_ _22214_/A _22214_/B _22214_/C vssd1 vssd1 vccd1 vccd1 _22214_/Y sky130_fd_sc_hd__nand3_1
XFILLER_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23194_ _23194_/A vssd1 vssd1 vccd1 vccd1 _23417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15286__A _15286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22145_ _22267_/A _22268_/A _22145_/C vssd1 vssd1 vccd1 vccd1 _22160_/B sky130_fd_sc_hd__nand3_2
XFILLER_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22076_ _22218_/B _22076_/B _22218_/A vssd1 vssd1 vccd1 vccd1 _22076_/X sky130_fd_sc_hd__and3b_1
XANTENNA__12422__B _19530_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21027_ _23562_/Q _20878_/A _20878_/B _20880_/A _21031_/A vssd1 vssd1 vccd1 vccd1
+ _21028_/B sky130_fd_sc_hd__a32o_1
XFILLER_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23139__A0 _18997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19358__A2 _17741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12800_ _20528_/C vssd1 vssd1 vccd1 vccd1 _20962_/B sky130_fd_sc_hd__clkbuf_2
X_13780_ _13842_/B vssd1 vssd1 vccd1 vccd1 _13836_/A sky130_fd_sc_hd__inv_2
X_22978_ _22978_/A vssd1 vssd1 vccd1 vccd1 _23321_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18566__B1 _12522_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21165__A2 _20966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12731_ _23448_/Q vssd1 vssd1 vccd1 vccd1 _13003_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21929_ _13469_/A _13599_/A _21922_/A _21922_/B _21928_/X vssd1 vssd1 vccd1 vccd1
+ _21938_/B sky130_fd_sc_hd__o221ai_4
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16041__A1 _12040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22566__B _22566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15450_ _15447_/Y _15448_/X _15420_/D _15420_/Y vssd1 vssd1 vccd1 vccd1 _15451_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12718_/C _12662_/B _12662_/C vssd1 vssd1 vccd1 vccd1 _12776_/A sky130_fd_sc_hd__nand3b_1
XFILLER_187_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14401_ _14438_/A _14438_/B _14442_/B vssd1 vssd1 vccd1 vccd1 _14410_/B sky130_fd_sc_hd__o21ai_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _19662_/C _15991_/A _12066_/A _12308_/A vssd1 vssd1 vccd1 vccd1 _11969_/B
+ sky130_fd_sc_hd__and4_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15382_/A _15382_/B _15382_/C vssd1 vssd1 vccd1 vccd1 _15383_/B sky130_fd_sc_hd__a21oi_1
XFILLER_168_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12593_ _23301_/Q vssd1 vssd1 vccd1 vccd1 _12688_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_716 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17120_ _17120_/A _17120_/B _17120_/C vssd1 vssd1 vccd1 vccd1 _17121_/A sky130_fd_sc_hd__nand3_1
XFILLER_128_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14332_ _14395_/A vssd1 vssd1 vccd1 vccd1 _14381_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17098__D _17108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17051_ _17050_/X _16794_/B _17434_/A _17435_/A vssd1 vssd1 vccd1 vccd1 _17744_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14263_ _13965_/X _13966_/X _14751_/B _14886_/B _14797_/A vssd1 vssd1 vccd1 vccd1
+ _14263_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16002_ _16268_/B _16002_/B _16248_/A _16249_/B vssd1 vssd1 vccd1 vccd1 _16008_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_7_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13214_ _23318_/Q vssd1 vssd1 vccd1 vccd1 _13224_/B sky130_fd_sc_hd__buf_2
XFILLER_87_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14194_ _14194_/A vssd1 vssd1 vccd1 vccd1 _15111_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15304__B1 _15301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _13196_/A _13196_/B vssd1 vssd1 vccd1 vccd1 _13146_/B sky130_fd_sc_hd__nand2_1
XFILLER_100_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _18149_/D _18144_/B _17954_/C vssd1 vssd1 vccd1 vccd1 _17955_/A sky130_fd_sc_hd__a21oi_1
X_13076_ _12903_/Y _12904_/X _12902_/C vssd1 vssd1 vccd1 vccd1 _13076_/X sky130_fd_sc_hd__o21a_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21928__B2 _21921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22050__B1 _22270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16904_ _16904_/A _16908_/A vssd1 vssd1 vccd1 vccd1 _16904_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12027_ _12016_/Y _12023_/Y _12026_/Y vssd1 vssd1 vccd1 vccd1 _12027_/Y sky130_fd_sc_hd__o21ai_4
X_17884_ _19951_/D vssd1 vssd1 vccd1 vccd1 _20164_/C sky130_fd_sc_hd__buf_2
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19623_ _19381_/X _19614_/X _19620_/X _19932_/A vssd1 vssd1 vccd1 vccd1 _19638_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16835_ _16828_/Y _16831_/X _16834_/Y vssd1 vssd1 vccd1 vccd1 _16836_/B sky130_fd_sc_hd__o21ai_1
XFILLER_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13618__B1 _22269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18006__C1 _18211_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19554_ _17050_/X _16794_/B _16816_/Y _16796_/X _18673_/A vssd1 vssd1 vccd1 vccd1
+ _19554_/X sky130_fd_sc_hd__a221o_2
XANTENNA__11890__C _16049_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16766_ _17010_/A _17009_/A vssd1 vssd1 vccd1 vccd1 _16766_/Y sky130_fd_sc_hd__nand2_1
X_13978_ _13978_/A _13978_/B vssd1 vssd1 vccd1 vccd1 _13984_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18505_ _12214_/X _16604_/X _18504_/Y vssd1 vssd1 vccd1 vccd1 _18505_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_94_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12929_ _12929_/A vssd1 vssd1 vccd1 vccd1 _20773_/C sky130_fd_sc_hd__buf_2
X_15717_ _16856_/D vssd1 vssd1 vccd1 vccd1 _15799_/A sky130_fd_sc_hd__buf_2
X_19485_ _19485_/A _19700_/A _19700_/B vssd1 vssd1 vccd1 vccd1 _19486_/B sky130_fd_sc_hd__and3_1
X_16697_ _16136_/A _16168_/C _16696_/Y vssd1 vssd1 vccd1 vccd1 _16699_/B sky130_fd_sc_hd__a21o_1
XANTENNA__22476__B _22476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_666 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18436_ _19279_/A _19280_/A vssd1 vssd1 vccd1 vccd1 _18749_/A sky130_fd_sc_hd__nor2_2
X_15648_ _15648_/A vssd1 vssd1 vccd1 vccd1 _16668_/C sky130_fd_sc_hd__buf_2
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19506__C1 _18481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14594__A1 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18367_ _23534_/Q _18362_/Y _18365_/Y _18366_/Y vssd1 vssd1 vccd1 vccd1 _18367_/Y
+ sky130_fd_sc_hd__o22ai_4
X_15579_ _15585_/D _15569_/B _23511_/Q vssd1 vssd1 vccd1 vccd1 _15580_/B sky130_fd_sc_hd__a21oi_1
XFILLER_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14275__A _14911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17318_ _17318_/A _17318_/B vssd1 vssd1 vccd1 vccd1 _17318_/Y sky130_fd_sc_hd__nand2_1
X_18298_ _18298_/A _18298_/B _18298_/C vssd1 vssd1 vccd1 vccd1 _18298_/X sky130_fd_sc_hd__or3_1
XFILLER_174_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17532__A1 _23524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17586__A _17586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19809__B1 _17613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17249_ _17249_/A vssd1 vssd1 vccd1 vccd1 _17249_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20260_ _20200_/B _20203_/B _20311_/A vssd1 vssd1 vccd1 vccd1 _20261_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__16921__C _16921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14722__B _23596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20191_ _20188_/A _20190_/Y _20189_/A vssd1 vssd1 vccd1 vccd1 _20247_/B sky130_fd_sc_hd__o21bai_2
XFILLER_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19951__D _19951_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22901_ _12788_/B input18/X _22907_/S vssd1 vssd1 vccd1 vccd1 _22902_/A sky130_fd_sc_hd__mux2_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_408 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22832_ _22861_/C _22637_/A _22637_/B _22830_/X _22861_/A vssd1 vssd1 vccd1 vccd1
+ _22834_/B sky130_fd_sc_hd__a32o_1
XFILLER_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18012__A2 _17032_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22763_ _22792_/C _22763_/B vssd1 vssd1 vccd1 vccd1 _22764_/C sky130_fd_sc_hd__and2b_1
XFILLER_198_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16665__A _16665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21714_ _21616_/X _21617_/X _21705_/A _21712_/Y vssd1 vssd1 vccd1 vccd1 _21715_/B
+ sky130_fd_sc_hd__o211a_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22694_ _22818_/A _22694_/B _22694_/C vssd1 vssd1 vccd1 vccd1 _22695_/B sky130_fd_sc_hd__and3_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14585__A1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21645_ _21645_/A _21645_/B _21645_/C vssd1 vssd1 vccd1 vccd1 _21646_/B sky130_fd_sc_hd__nor3_1
XANTENNA__12045__C1 _19381_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14585__B2 _12675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21855__B1 _13870_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21576_ _21576_/A vssd1 vssd1 vccd1 vccd1 _21694_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12417__B _19804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23315_ _23347_/CLK _23315_/D vssd1 vssd1 vccd1 vccd1 _23315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20527_ _20528_/A _20527_/B _23454_/Q vssd1 vssd1 vccd1 vccd1 _20676_/A sky130_fd_sc_hd__nand3_2
XFILLER_197_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22186__A_N _22142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23246_ _23441_/Q input26/X _23250_/S vssd1 vssd1 vccd1 vccd1 _23247_/A sky130_fd_sc_hd__mux2_1
X_20458_ _23560_/Q vssd1 vssd1 vccd1 vccd1 _20608_/A sky130_fd_sc_hd__inv_2
XFILLER_134_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23177_ _23177_/A vssd1 vssd1 vccd1 vccd1 _23410_/D sky130_fd_sc_hd__clkbuf_1
X_20389_ _20341_/X _20340_/Y _20361_/Y _20415_/B _20415_/A vssd1 vssd1 vccd1 vccd1
+ _20392_/B sky130_fd_sc_hd__a32o_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19028__A1 _11948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22128_ _13547_/A _13599_/X _22122_/Y vssd1 vssd1 vccd1 vccd1 _22128_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14950_ _14932_/X _14947_/Y _14948_/Y _14949_/Y vssd1 vssd1 vccd1 vccd1 _14953_/C
+ sky130_fd_sc_hd__o211ai_2
X_22059_ _22377_/A vssd1 vssd1 vccd1 vccd1 _22059_/X sky130_fd_sc_hd__buf_2
XANTENNA__11859__C1 _16796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13901_ _23354_/Q _13901_/B _13966_/A vssd1 vssd1 vccd1 vccd1 _14068_/A sky130_fd_sc_hd__nand3b_1
X_14881_ _14756_/B _15000_/A _14893_/A vssd1 vssd1 vccd1 vccd1 _15004_/B sky130_fd_sc_hd__o21ai_4
XANTENNA_input28_A wb_dat_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16620_ _16795_/A _17963_/C _16620_/C vssd1 vssd1 vccd1 vccd1 _16621_/A sky130_fd_sc_hd__nand3_1
X_13832_ _13645_/B _13645_/C _13822_/Y vssd1 vssd1 vccd1 vccd1 _13834_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16551_ _16549_/A _16364_/A _16364_/B _16529_/A _16544_/B vssd1 vssd1 vccd1 vccd1
+ _16551_/X sky130_fd_sc_hd__a32o_1
XANTENNA__19200__A1 _11936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13763_ _13763_/A _13763_/B _13763_/C vssd1 vssd1 vccd1 vccd1 _21857_/A sky130_fd_sc_hd__nand3_1
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22296__B _22476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15502_ _15502_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _15503_/B sky130_fd_sc_hd__nor2_2
X_12714_ _12714_/A vssd1 vssd1 vccd1 vccd1 _12714_/X sky130_fd_sc_hd__buf_2
X_19270_ _19075_/C _19075_/B _19075_/A _19087_/A _19082_/X vssd1 vssd1 vccd1 vccd1
+ _19298_/B sky130_fd_sc_hd__a32oi_4
X_16482_ _16478_/X _16458_/X _16481_/X _16384_/X _16356_/X vssd1 vssd1 vccd1 vccd1
+ _16482_/X sky130_fd_sc_hd__o32a_1
XFILLER_16_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13694_ _13595_/Y _13596_/Y _13760_/A _13760_/B vssd1 vssd1 vccd1 vccd1 _13694_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_188_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18221_ _20210_/D vssd1 vssd1 vccd1 vccd1 _20265_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15433_ _15433_/A _15433_/B vssd1 vssd1 vccd1 vccd1 _15434_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14576__A1 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12645_ _12644_/X _12688_/B _12712_/A vssd1 vssd1 vccd1 vccd1 _20675_/A sky130_fd_sc_hd__a21o_1
XFILLER_188_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14576__B2 _14863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22638__A2 _22164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18152_ _18262_/C _18262_/A vssd1 vssd1 vccd1 vccd1 _23591_/D sky130_fd_sc_hd__xor2_2
XFILLER_157_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15364_ _15420_/C _15363_/A _15363_/B _15363_/C vssd1 vssd1 vccd1 vccd1 _15366_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_196_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12576_ _12874_/D vssd1 vssd1 vccd1 vccd1 _12577_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12327__B _12346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14315_ _14355_/C vssd1 vssd1 vccd1 vccd1 _14407_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_17103_ _14599_/X _16203_/Y _15791_/X _16213_/A _19659_/C vssd1 vssd1 vccd1 vccd1
+ _17104_/B sky130_fd_sc_hd__o311a_2
XFILLER_184_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18083_ _20269_/D _18219_/D _18272_/A _20271_/A _17962_/X vssd1 vssd1 vccd1 vccd1
+ _18084_/B sky130_fd_sc_hd__a41o_1
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15919__A _15937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15295_ _14588_/X _14050_/X _14061_/X _14901_/X _15353_/C vssd1 vssd1 vccd1 vccd1
+ _15300_/A sky130_fd_sc_hd__o311a_1
XFILLER_184_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17034_ _18163_/B vssd1 vssd1 vccd1 vccd1 _18335_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_output96_A _23579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19267__A1 _19265_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14246_ _14246_/A _14246_/B vssd1 vssd1 vccd1 vccd1 _14282_/C sky130_fd_sc_hd__nand2_1
XFILLER_171_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14177_ _14177_/A _14177_/B vssd1 vssd1 vccd1 vccd1 _14180_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12343__A _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13172_/B _13128_/B vssd1 vssd1 vccd1 vccd1 _13136_/A sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_2_3_0_bq_clk_i_A clkbuf_2_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13158__B _21182_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20560__A _23456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _11764_/A _18490_/A _18984_/B vssd1 vssd1 vccd1 vccd1 _18985_/X sky130_fd_sc_hd__o21a_1
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _18207_/A _18208_/A _17933_/X _18198_/C vssd1 vssd1 vccd1 vccd1 _17936_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13059_ _12827_/A _12766_/A _13058_/B vssd1 vssd1 vccd1 vccd1 _13059_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_714 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater104 _23479_/Q vssd1 vssd1 vccd1 vccd1 _13769_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater115 _23425_/CLK vssd1 vssd1 vccd1 vccd1 _23424_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16469__B _16469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater126 _23445_/CLK vssd1 vssd1 vccd1 vccd1 _23444_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater137 _23402_/CLK vssd1 vssd1 vccd1 vccd1 _23365_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17867_ _17880_/A _17880_/B vssd1 vssd1 vccd1 vccd1 _17867_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater148 _23309_/CLK vssd1 vssd1 vccd1 vccd1 _23307_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater159 input39/X vssd1 vssd1 vccd1 vccd1 _23184_/B sky130_fd_sc_hd__clkbuf_1
X_19606_ _19609_/B _19598_/Y _19601_/X _19600_/Y vssd1 vssd1 vccd1 vccd1 _19606_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_16818_ _16816_/Y _16796_/X _16794_/B _17050_/A vssd1 vssd1 vccd1 vccd1 _17449_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17798_ _17798_/A _17919_/A _17798_/C vssd1 vssd1 vccd1 vccd1 _17798_/X sky130_fd_sc_hd__and3_1
XFILLER_4_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22487__A _22487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19537_ _19701_/A vssd1 vssd1 vccd1 vccd1 _19537_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16749_ _16749_/A _18157_/C _16749_/C vssd1 vssd1 vccd1 vccd1 _16749_/X sky130_fd_sc_hd__and3_1
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19468_ _19468_/A vssd1 vssd1 vccd1 vccd1 _19755_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12290__A2 _12279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18419_ _18420_/B _18420_/C _23537_/Q vssd1 vssd1 vccd1 vccd1 _18430_/A sky130_fd_sc_hd__a21boi_2
XFILLER_179_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14567__A1 _15762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19399_ _19399_/A _19399_/B _19399_/C vssd1 vssd1 vccd1 vccd1 _19406_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12518__A _17456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21430_ _21432_/A _21432_/B _21430_/C vssd1 vssd1 vccd1 vccd1 _21635_/C sky130_fd_sc_hd__nand3_2
XANTENNA__12042__A2 _12040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20104__A3 _18335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18850__D _19334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21361_ _21635_/A _20471_/Y _21360_/Y vssd1 vssd1 vccd1 vccd1 _21453_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__14319__B2 _15082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14733__A _23260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23100_ _23376_/Q input25/X _23106_/S vssd1 vssd1 vccd1 vccd1 _23101_/A sky130_fd_sc_hd__mux2_1
XANTENNA__23468__D _23480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20312_ _20312_/A _20312_/B _20312_/C vssd1 vssd1 vccd1 vccd1 _20313_/B sky130_fd_sc_hd__and3_1
XFILLER_135_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21292_ _20502_/X _20504_/X _21193_/C _21431_/A vssd1 vssd1 vccd1 vccd1 _21292_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_190_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17269__B1 _16311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23031_ _23031_/A vssd1 vssd1 vccd1 vccd1 _23345_/D sky130_fd_sc_hd__clkbuf_1
X_20243_ _20243_/A _20243_/B vssd1 vssd1 vccd1 vccd1 _20243_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20174_ _20095_/C _20095_/A _20172_/B _20175_/A _20283_/B vssd1 vssd1 vccd1 vccd1
+ _20176_/B sky130_fd_sc_hd__a32o_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15295__A2 _14050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17036__A3 _18335_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11856__A2 _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18875__A _18875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12700__B _21271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_706 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22815_ _22859_/A _22815_/B vssd1 vssd1 vccd1 vccd1 _22817_/B sky130_fd_sc_hd__xor2_1
XFILLER_16_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22746_ _22694_/B _22694_/C _22821_/C _22821_/A vssd1 vssd1 vccd1 vccd1 _22747_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_243 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13531__B _22380_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22677_ _22677_/A vssd1 vssd1 vccd1 vccd1 _22677_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12430_ _12425_/X _12427_/X _12429_/Y vssd1 vssd1 vccd1 vccd1 _12441_/A sky130_fd_sc_hd__o21ai_1
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21628_ _21625_/X _21626_/Y _21540_/C _21627_/Y vssd1 vssd1 vccd1 vccd1 _21660_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_40_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12361_ _12336_/A _12360_/Y _12330_/X vssd1 vssd1 vccd1 vccd1 _12363_/C sky130_fd_sc_hd__a21o_1
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21559_ _21559_/A _21559_/B _21559_/C vssd1 vssd1 vccd1 vccd1 _21559_/X sky130_fd_sc_hd__or3_1
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14100_ _14178_/B _14374_/D _14178_/A vssd1 vssd1 vccd1 vccd1 _14976_/A sky130_fd_sc_hd__nand3_4
XFILLER_181_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15080_ _15076_/Y _15078_/X _15079_/Y vssd1 vssd1 vccd1 vccd1 _15080_/X sky130_fd_sc_hd__o21a_1
X_12292_ _11717_/B _11717_/C _12238_/X _12374_/A vssd1 vssd1 vccd1 vccd1 _12292_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16180__B1 _15985_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14031_ _14077_/C vssd1 vssd1 vccd1 vccd1 _14031_/X sky130_fd_sc_hd__clkbuf_4
X_23229_ _23229_/A vssd1 vssd1 vccd1 vccd1 _23433_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18457__C1 _16526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20264__C1 _20368_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18770_ _18771_/A _18966_/A _18966_/B vssd1 vssd1 vccd1 vccd1 _18773_/C sky130_fd_sc_hd__a21o_1
XFILLER_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15982_ _15982_/A _15982_/B vssd1 vssd1 vccd1 vccd1 _15985_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17721_ _16683_/X _16667_/C _16667_/D _17029_/X vssd1 vssd1 vccd1 vccd1 _17723_/A
+ sky130_fd_sc_hd__a31o_2
X_14933_ _14933_/A _23505_/Q vssd1 vssd1 vccd1 vccd1 _14944_/A sky130_fd_sc_hd__nand2_1
XFILLER_76_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15038__A2 _15075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17652_ _17656_/A _17656_/B _17657_/B _17657_/C vssd1 vssd1 vccd1 vccd1 _17653_/C
+ sky130_fd_sc_hd__nand4_1
X_14864_ _14868_/D _14864_/B _14864_/C _15112_/C vssd1 vssd1 vccd1 vccd1 _14864_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _16647_/A _16608_/A vssd1 vssd1 vccd1 vccd1 _16607_/A sky130_fd_sc_hd__nand2_1
X_13815_ _13279_/A _13418_/A _13814_/Y vssd1 vssd1 vccd1 vccd1 _13818_/A sky130_fd_sc_hd__o21ai_2
X_17583_ _17583_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17585_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14795_ _14795_/A _14795_/B _14795_/C vssd1 vssd1 vccd1 vccd1 _14795_/Y sky130_fd_sc_hd__nand3_1
XFILLER_63_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19322_ _19525_/A _19524_/A _19517_/B vssd1 vssd1 vccd1 vccd1 _19477_/A sky130_fd_sc_hd__a21o_1
XFILLER_188_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16534_ _16533_/Y _16519_/Y _16522_/B vssd1 vssd1 vccd1 vccd1 _16534_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_32_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13746_ _13711_/A _13711_/B _13711_/C vssd1 vssd1 vccd1 vccd1 _13748_/B sky130_fd_sc_hd__a21o_1
XFILLER_91_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19253_ _19069_/A _19069_/B _19069_/C _19071_/X _19249_/X vssd1 vssd1 vccd1 vccd1
+ _19259_/A sky130_fd_sc_hd__a32o_1
XFILLER_149_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13441__B _13810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16465_ _16464_/X _16447_/Y _12238_/X _16398_/X _16399_/X vssd1 vssd1 vccd1 vccd1
+ _16465_/Y sky130_fd_sc_hd__o221ai_4
X_13677_ _13538_/X _13477_/A _13462_/A vssd1 vssd1 vccd1 vccd1 _13682_/A sky130_fd_sc_hd__a21boi_1
XFILLER_189_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18204_ _23532_/Q _18204_/B _18204_/C vssd1 vssd1 vccd1 vccd1 _18263_/A sky130_fd_sc_hd__nand3b_1
XFILLER_148_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22754__B _22754_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15416_ _15416_/A vssd1 vssd1 vccd1 vccd1 _15485_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_12628_ _20628_/C vssd1 vssd1 vccd1 vccd1 _21035_/C sky130_fd_sc_hd__clkbuf_4
X_16396_ _16396_/A _16396_/B vssd1 vssd1 vccd1 vccd1 _16397_/A sky130_fd_sc_hd__nand2_1
X_19184_ _19184_/A vssd1 vssd1 vccd1 vccd1 _19858_/A sky130_fd_sc_hd__buf_2
XFILLER_157_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18135_ _17957_/Y _18129_/Y _18132_/X _18155_/B vssd1 vssd1 vccd1 vccd1 _18136_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__17499__B1 _17152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15347_ _15293_/A _15293_/B _15332_/B vssd1 vssd1 vccd1 vccd1 _15391_/B sky130_fd_sc_hd__o21a_1
X_12559_ _19089_/A _12545_/Y _12558_/X vssd1 vssd1 vccd1 vccd1 _18733_/A sky130_fd_sc_hd__o21ai_2
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18066_ _18144_/C _18149_/B _18066_/C vssd1 vssd1 vccd1 vccd1 _18067_/B sky130_fd_sc_hd__and3_1
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15278_ _15277_/A _15277_/B _15277_/C vssd1 vssd1 vccd1 vccd1 _15279_/B sky130_fd_sc_hd__a21o_1
XFILLER_176_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17017_ _17017_/A _17017_/B _23522_/Q vssd1 vssd1 vccd1 vccd1 _17018_/B sky130_fd_sc_hd__nand3_1
X_14229_ _14230_/A _14302_/B _14229_/C _14229_/D vssd1 vssd1 vccd1 vccd1 _14235_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_172_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19660__A1 _11936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18968_ _18968_/A _19246_/A vssd1 vssd1 vccd1 vccd1 _19059_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22547__B2 _22126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17919_ _17919_/A _17919_/B _17919_/C _17919_/D vssd1 vssd1 vccd1 vccd1 _17920_/C
+ sky130_fd_sc_hd__nand4_2
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18899_ _18899_/A _18899_/B _18899_/C vssd1 vssd1 vccd1 vccd1 _19091_/B sky130_fd_sc_hd__nand3_1
XFILLER_113_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20930_ _12709_/X _21592_/A _20919_/Y _20929_/Y vssd1 vssd1 vccd1 vccd1 _20941_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_187_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20861_ _20885_/A _20869_/B vssd1 vssd1 vccd1 vccd1 _20863_/A sky130_fd_sc_hd__nand2_1
XANTENNA__22010__A _22064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22600_ _22541_/X _22596_/Y _22597_/Y _22599_/Y vssd1 vssd1 vccd1 vccd1 _22633_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_23_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23580_ _23588_/CLK _23580_/D vssd1 vssd1 vccd1 vccd1 _23580_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20792_ _20625_/B _20778_/A _20627_/Y vssd1 vssd1 vccd1 vccd1 _20793_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__22180__C1 _21853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15042__A1_N _15044_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22531_ _22529_/A _22629_/A _22528_/A _22528_/B vssd1 vssd1 vccd1 vccd1 _22532_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15737__B1 _14553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12248__A _16198_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19479__A1 _18476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22462_ _13470_/X _22461_/X _22393_/A vssd1 vssd1 vccd1 vccd1 _22463_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12015__A2 _12013_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16662__B _16662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21413_ _21410_/Y _21411_/Y _21418_/A vssd1 vssd1 vccd1 vccd1 _21413_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15559__A _15559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22393_ _22393_/A _22393_/B vssd1 vssd1 vccd1 vccd1 _22394_/C sky130_fd_sc_hd__nand2_1
XFILLER_148_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21344_ _21344_/A _21344_/B vssd1 vssd1 vccd1 vccd1 _21345_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21275_ _21327_/A _21327_/B vssd1 vssd1 vccd1 vccd1 _21311_/A sky130_fd_sc_hd__nand2_2
XFILLER_190_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23014_ _23025_/A vssd1 vssd1 vccd1 vccd1 _23023_/S sky130_fd_sc_hd__clkbuf_2
X_20226_ _20158_/B _20159_/B _20224_/Y _20225_/X vssd1 vssd1 vccd1 vccd1 _20283_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_103_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16465__A1 _16464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20157_ _20135_/X _20136_/X _20156_/Y vssd1 vssd1 vccd1 vccd1 _20159_/A sky130_fd_sc_hd__o21ai_1
XFILLER_104_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12711__A _20799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20088_ _20095_/C vssd1 vssd1 vccd1 vccd1 _20090_/A sky130_fd_sc_hd__inv_2
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _11686_/B _11676_/X _11677_/X vssd1 vssd1 vccd1 vccd1 _11931_/B sky130_fd_sc_hd__o21ai_4
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17965__A1 _14729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20564__A3 _13061_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18755__D _18755_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _11861_/A _18470_/C _12245_/A vssd1 vssd1 vccd1 vccd1 _11887_/C sky130_fd_sc_hd__nand3_2
XFILLER_73_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _21766_/A _21767_/A _13600_/C vssd1 vssd1 vccd1 vccd1 _13616_/A sky130_fd_sc_hd__nand3_2
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _23268_/Q _14520_/X _14547_/X _12712_/X vssd1 vssd1 vccd1 vccd1 _14580_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17717__A1 _16408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ _11792_/A _11792_/B vssd1 vssd1 vccd1 vccd1 _11886_/A sky130_fd_sc_hd__nand2_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13531_ _13561_/A _22380_/C _13709_/C _22278_/B vssd1 vssd1 vccd1 vccd1 _13531_/X
+ sky130_fd_sc_hd__and4_1
X_22729_ _22729_/A _22729_/B _22729_/C vssd1 vssd1 vccd1 vccd1 _22730_/A sky130_fd_sc_hd__nor3_1
XFILLER_159_939 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16250_ _16005_/Y _16249_/Y _16248_/A vssd1 vssd1 vccd1 vccd1 _16258_/A sky130_fd_sc_hd__o21ai_1
XFILLER_159_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _13462_/A vssd1 vssd1 vccd1 vccd1 _13598_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15201_ _15201_/A _15201_/B vssd1 vssd1 vccd1 vccd1 _15203_/A sky130_fd_sc_hd__xor2_1
XFILLER_139_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12413_ _12413_/A vssd1 vssd1 vccd1 vccd1 _18460_/A sky130_fd_sc_hd__buf_2
XFILLER_127_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16181_ _16181_/A _16181_/B vssd1 vssd1 vccd1 vccd1 _16181_/X sky130_fd_sc_hd__and2_1
XFILLER_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13393_ _21764_/B vssd1 vssd1 vccd1 vccd1 _22264_/B sky130_fd_sc_hd__buf_2
XFILLER_167_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15132_ _15132_/A _15132_/B _15132_/C vssd1 vssd1 vccd1 vccd1 _15134_/B sky130_fd_sc_hd__nand3_1
XFILLER_166_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12344_ _19530_/A vssd1 vssd1 vccd1 vccd1 _19903_/C sky130_fd_sc_hd__buf_2
XFILLER_182_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_964 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12605__B _12678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19940_ _19835_/Y _19836_/Y _19833_/X vssd1 vssd1 vccd1 vccd1 _19940_/X sky130_fd_sc_hd__o21a_1
XFILLER_181_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_62 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12309__A3 _16364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15063_ _15063_/A vssd1 vssd1 vccd1 vccd1 _15063_/Y sky130_fd_sc_hd__inv_2
X_12275_ _11788_/Y _11803_/X _11880_/X vssd1 vssd1 vccd1 vccd1 _12275_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_880 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18499__B _18499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ _14017_/A _14024_/B vssd1 vssd1 vccd1 vccd1 _14015_/C sky130_fd_sc_hd__nand2_1
X_19871_ _16464_/X _20081_/D _19304_/X _19525_/D vssd1 vssd1 vccd1 vccd1 _19871_/X
+ sky130_fd_sc_hd__o31a_1
X_18822_ _12105_/Y _18835_/A _19029_/A vssd1 vssd1 vccd1 vccd1 _18825_/A sky130_fd_sc_hd__o21ai_1
XFILLER_68_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23592__CLK _23598_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18753_ _18784_/A _18753_/B vssd1 vssd1 vccd1 vccd1 _18773_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15965_ _16523_/C _17456_/A _15964_/Y vssd1 vssd1 vccd1 vccd1 _16132_/A sky130_fd_sc_hd__o21ai_2
XFILLER_49_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17704_ _18059_/B vssd1 vssd1 vccd1 vccd1 _18256_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15932__A _15932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18602__C1 _17761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14916_ _14975_/C _14915_/X _14890_/A _14775_/Y _14778_/B vssd1 vssd1 vccd1 vccd1
+ _14918_/A sky130_fd_sc_hd__a32oi_4
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18684_ _12184_/X _12185_/X _12464_/Y _11961_/Y vssd1 vssd1 vccd1 vccd1 _18684_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_15896_ _15985_/C _15866_/B _15879_/Y _15888_/Y vssd1 vssd1 vccd1 vccd1 _15896_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_63_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17635_ _17635_/A vssd1 vssd1 vccd1 vccd1 _18002_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14847_ _14847_/A _14847_/B vssd1 vssd1 vccd1 vccd1 _14847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17566_ _17566_/A vssd1 vssd1 vccd1 vccd1 _17566_/X sky130_fd_sc_hd__buf_2
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14778_ _14778_/A _14778_/B vssd1 vssd1 vccd1 vccd1 _14781_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19305_ _11799_/X _11801_/X _19651_/A _19652_/A vssd1 vssd1 vccd1 vccd1 _19305_/Y
+ sky130_fd_sc_hd__o211ai_1
X_16517_ _16415_/B _16517_/B _16517_/C vssd1 vssd1 vccd1 vccd1 _16518_/B sky130_fd_sc_hd__nand3b_1
XFILLER_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13729_ _13728_/X _13723_/Y _13727_/A vssd1 vssd1 vccd1 vccd1 _13729_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17497_ _17497_/A _17497_/B _17497_/C _17497_/D vssd1 vssd1 vccd1 vccd1 _17498_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_189_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19236_ _19227_/Y _19233_/Y _19257_/A _19257_/B vssd1 vssd1 vccd1 vccd1 _19236_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16448_ _16360_/X _16447_/Y _16398_/X _12279_/A _16399_/X vssd1 vssd1 vccd1 vccd1
+ _16448_/X sky130_fd_sc_hd__o221a_1
XANTENNA__16931__A2 _16377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19167_ _19167_/A _19167_/B _19167_/C vssd1 vssd1 vccd1 vccd1 _19168_/A sky130_fd_sc_hd__nand3_4
X_16379_ _16379_/A _16379_/B vssd1 vssd1 vccd1 vccd1 _16404_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11700__A _15699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18118_ _18118_/A _18298_/B _18156_/B vssd1 vssd1 vccd1 vccd1 _18245_/A sky130_fd_sc_hd__or3b_1
XFILLER_173_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19098_ _18919_/X _19443_/B _19106_/A _19108_/A _19095_/Y vssd1 vssd1 vccd1 vccd1
+ _19101_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_172_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17892__B1 _16408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18049_ _18053_/A _18049_/B vssd1 vssd1 vccd1 vccd1 _18059_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16695__B2 _16706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14433__D _14433_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21060_ _21097_/B vssd1 vssd1 vccd1 vccd1 _21095_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22005__A _22076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22232__A3 _21988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20011_ _20011_/A _20011_/B _20011_/C vssd1 vssd1 vccd1 vccd1 _20012_/C sky130_fd_sc_hd__nand3_1
XFILLER_115_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19017__C _19364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21991__A2 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23193__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15842__A _16591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21962_ _22118_/A vssd1 vssd1 vccd1 vccd1 _22117_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22940__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20913_ _21174_/C vssd1 vssd1 vccd1 vccd1 _21369_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_344 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21893_ _21893_/A _21893_/B vssd1 vssd1 vccd1 vccd1 _21893_/Y sky130_fd_sc_hd__nor2_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20844_ _20719_/X _20731_/Y _20841_/Y _20843_/Y vssd1 vssd1 vccd1 vccd1 _20845_/A
+ sky130_fd_sc_hd__o211ai_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23563_ _23571_/CLK _23563_/D vssd1 vssd1 vccd1 vccd1 _23563_/Q sky130_fd_sc_hd__dfxtp_2
X_20775_ _20775_/A _21000_/A _20775_/C _20775_/D vssd1 vssd1 vccd1 vccd1 _20776_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_74_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22514_ _22513_/A _22513_/B _22513_/C vssd1 vssd1 vccd1 vccd1 _22516_/D sky130_fd_sc_hd__a21o_1
XFILLER_167_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23494_ _23510_/CLK _23506_/Q vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23465__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22445_ _22247_/Y _22445_/B _22445_/C _22445_/D vssd1 vssd1 vccd1 vccd1 _22445_/Y
+ sky130_fd_sc_hd__nand4b_1
XFILLER_183_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_780 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22376_ _22409_/A _22504_/A _22504_/B vssd1 vssd1 vccd1 vccd1 _22400_/B sky130_fd_sc_hd__nand3_1
XFILLER_159_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_88 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21327_ _21327_/A _21327_/B _21327_/C _21327_/D vssd1 vssd1 vccd1 vccd1 _21330_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_190_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ _12059_/A _12200_/B _12205_/A _12059_/D vssd1 vssd1 vccd1 vccd1 _12064_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21258_ _21025_/A _21029_/X _21031_/Y _21146_/B vssd1 vssd1 vccd1 vccd1 _21258_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_132_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16438__A1 _16437_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20209_ _20209_/A vssd1 vssd1 vccd1 vccd1 _20265_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21189_ _21212_/A _21212_/B _21185_/X _21188_/Y vssd1 vssd1 vccd1 vccd1 _21217_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_78_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21176__D _21182_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _16593_/A _16860_/C _15860_/C _15968_/A vssd1 vssd1 vccd1 vccd1 _15750_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12962_ _12962_/A _12962_/B _12962_/C vssd1 vssd1 vccd1 vccd1 _13141_/B sky130_fd_sc_hd__nand3_1
XFILLER_79_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A wb_dat_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _11913_/A _11913_/B _11913_/C vssd1 vssd1 vccd1 vccd1 _12253_/A sky130_fd_sc_hd__nand3_1
X_14701_ _23375_/Q _14688_/X _14700_/X vssd1 vssd1 vccd1 vccd1 _14701_/X sky130_fd_sc_hd__o21a_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21192__C _21295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ _12899_/B _12899_/C _12899_/A vssd1 vssd1 vccd1 vccd1 _12893_/Y sky130_fd_sc_hd__a21oi_2
X_15681_ _15974_/D vssd1 vssd1 vccd1 vccd1 _15682_/D sky130_fd_sc_hd__clkbuf_4
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _19949_/A _17420_/B _19674_/B _17860_/A vssd1 vssd1 vccd1 vccd1 _17420_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13272__A _13498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _11844_/A _11844_/B _12053_/A vssd1 vssd1 vccd1 vccd1 _11844_/Y sky130_fd_sc_hd__nor3_2
X_14632_ _23363_/Q vssd1 vssd1 vccd1 vccd1 _14632_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23180__S _23182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _17351_/A _17351_/B _17351_/C vssd1 vssd1 vccd1 vccd1 _17358_/B sky130_fd_sc_hd__nand3_1
X_14563_ _23265_/Q _14520_/X _14526_/X _12678_/C vssd1 vssd1 vccd1 vccd1 _14563_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _12419_/A vssd1 vssd1 vccd1 vccd1 _18859_/C sky130_fd_sc_hd__buf_2
XANTENNA__13975__A2 _13945_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _11649_/X _16140_/A _12036_/B _11695_/X vssd1 vssd1 vccd1 vccd1 _16302_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_198_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13514_ _13448_/A _13517_/C _13513_/A vssd1 vssd1 vccd1 vccd1 _13515_/C sky130_fd_sc_hd__a21o_1
X_17282_ _17270_/Y _17273_/Y _17268_/C _17276_/B vssd1 vssd1 vccd1 vccd1 _17282_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14494_ _14454_/Y _14488_/Y _14496_/B _14496_/A vssd1 vssd1 vccd1 vccd1 _14497_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19021_ _12282_/B _11686_/Y _12464_/Y _11961_/Y _11689_/Y vssd1 vssd1 vccd1 vccd1
+ _19021_/X sky130_fd_sc_hd__a221o_2
X_13445_ _13599_/A _13425_/Y _13443_/B vssd1 vssd1 vccd1 vccd1 _13446_/A sky130_fd_sc_hd__o21ai_1
X_16233_ _16233_/A _16233_/B _16710_/A vssd1 vssd1 vccd1 vccd1 _16234_/C sky130_fd_sc_hd__nand3_1
XANTENNA__12616__A _13121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16164_ _16638_/A _16639_/A vssd1 vssd1 vccd1 vccd1 _16165_/A sky130_fd_sc_hd__nand2_1
X_13376_ _13376_/A _13376_/B _21766_/A vssd1 vssd1 vccd1 vccd1 _13433_/B sky130_fd_sc_hd__nand3_2
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12327_ _12327_/A _12346_/A vssd1 vssd1 vccd1 vccd1 _12327_/Y sky130_fd_sc_hd__nand2_2
XFILLER_115_828 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15115_ _23364_/Q _15115_/B _15115_/C _15115_/D vssd1 vssd1 vccd1 vccd1 _15233_/B
+ sky130_fd_sc_hd__nand4b_4
XFILLER_127_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16095_ _16331_/B _16326_/B vssd1 vssd1 vccd1 vccd1 _16096_/A sky130_fd_sc_hd__nand2_2
XFILLER_5_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17845__C _17845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23566__D _23566_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19923_ _19923_/A _19923_/B vssd1 vssd1 vccd1 vccd1 _19923_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15046_ _15050_/A _15050_/B _15050_/C vssd1 vssd1 vccd1 vccd1 _15049_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__19615__A1 _19381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12258_ _12308_/A _16364_/A _16364_/B _12260_/D _19503_/C vssd1 vssd1 vccd1 vccd1
+ _12273_/B sky130_fd_sc_hd__a32o_2
X_19854_ _19855_/A _19855_/B _19649_/A _19649_/B vssd1 vssd1 vccd1 vccd1 _19943_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189_ _12189_/A vssd1 vssd1 vccd1 vccd1 _17098_/C sky130_fd_sc_hd__buf_2
XFILLER_95_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11910__A1 _11969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18805_ _18805_/A _18972_/B _18972_/C vssd1 vssd1 vccd1 vccd1 _18806_/B sky130_fd_sc_hd__and3_1
Xclkbuf_4_3_0_bq_clk_i clkbuf_4_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _23518_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13166__B _13177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19785_ _20120_/A vssd1 vssd1 vccd1 vccd1 _19785_/X sky130_fd_sc_hd__buf_2
X_16997_ _23523_/Q _16997_/B _16997_/C vssd1 vssd1 vccd1 vccd1 _17019_/A sky130_fd_sc_hd__nand3b_1
XFILLER_95_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22479__B _22479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18736_ _18731_/X _18732_/Y _18733_/Y _18922_/A vssd1 vssd1 vccd1 vccd1 _18738_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15948_ _15948_/A _15948_/B _15948_/C vssd1 vssd1 vccd1 vccd1 _15949_/A sky130_fd_sc_hd__and3_1
XANTENNA__12466__A2 _12463_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12320__D1 _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18667_ _18627_/Y _18628_/X _18665_/Y _18666_/X vssd1 vssd1 vccd1 vccd1 _18667_/Y
+ sky130_fd_sc_hd__o211ai_2
X_15879_ _15879_/A _15879_/B vssd1 vssd1 vccd1 vccd1 _15879_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17618_ _17589_/Y _17597_/Y _17606_/X vssd1 vssd1 vccd1 vccd1 _17618_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18598_ _18598_/A vssd1 vssd1 vccd1 vccd1 _18599_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23488__CLK _23492_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17549_ _17549_/A _17810_/D _17549_/C vssd1 vssd1 vccd1 vccd1 _17553_/A sky130_fd_sc_hd__nand3_1
XFILLER_51_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17157__A2 _17155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20560_ _23456_/Q _20704_/B vssd1 vssd1 vccd1 vccd1 _20562_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19219_ _19218_/X _18000_/A _19194_/X _19196_/Y vssd1 vssd1 vccd1 vccd1 _19219_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_192_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14915__A1 _14588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20491_ _20634_/B _20487_/X _20488_/Y _20490_/Y vssd1 vssd1 vccd1 vccd1 _20492_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_164_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22230_ _22207_/A _22207_/B _22207_/C _22225_/C vssd1 vssd1 vccd1 vccd1 _22231_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_30_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16117__B1 _15926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19854__B2 _19649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_997 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22161_ _22040_/B _22271_/A _22160_/Y vssd1 vssd1 vccd1 vccd1 _22162_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__15837__A _16062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20462__B _23458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21112_ _20980_/A _21111_/Y _20981_/Y vssd1 vssd1 vccd1 vccd1 _21113_/C sky130_fd_sc_hd__o21a_1
XFILLER_132_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22092_ _22093_/A _22093_/B _22093_/C _22084_/A vssd1 vssd1 vccd1 vccd1 _22094_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15891__A2 _15866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21043_ _21043_/A vssd1 vssd1 vccd1 vccd1 _21635_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19970__C _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17093__A1 _15621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input2_A wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22994_ _22994_/A vssd1 vssd1 vccd1 vccd1 _23328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13804__B _13804_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21945_ _21936_/Y _21941_/Y _21943_/X _21944_/X vssd1 vssd1 vccd1 vccd1 _21946_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14188__A _14188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19698__B _19903_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12209__A2 _11815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13406__A1 _21778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21876_ _21875_/Y _21782_/C _21806_/A vssd1 vssd1 vccd1 vccd1 _21946_/A sky130_fd_sc_hd__o21ai_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ _20828_/B _20828_/C _20828_/A vssd1 vssd1 vccd1 vccd1 _21121_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23546_ _23578_/CLK _23546_/D vssd1 vssd1 vccd1 vccd1 _23546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20152__A1 _19539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20758_ _21414_/A _21415_/A vssd1 vssd1 vccd1 vccd1 _21542_/A sky130_fd_sc_hd__nor2_2
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23477_ _23499_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 _23477_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_149_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20689_ _20715_/A _20715_/B vssd1 vssd1 vccd1 vccd1 _20690_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13230_ _13659_/A vssd1 vssd1 vccd1 vccd1 _13563_/C sky130_fd_sc_hd__clkbuf_2
X_22428_ _22428_/A _22428_/B _22516_/A _22428_/D vssd1 vssd1 vccd1 vccd1 _22430_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19845__A1 _19504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17305__C1 _17631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17939__B1_N _23529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16659__A1 _15932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13161_ _13157_/Y _13158_/Y _13168_/B vssd1 vssd1 vccd1 vccd1 _13162_/B sky130_fd_sc_hd__o21ai_1
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22359_ _22324_/B _22324_/C _22324_/A vssd1 vssd1 vccd1 vccd1 _22359_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_136_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17320__A2 _16480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12112_ _19157_/C vssd1 vssd1 vccd1 vccd1 _17133_/C sky130_fd_sc_hd__buf_2
X_13092_ _13083_/Y _13088_/X _13090_/Y _13091_/Y vssd1 vssd1 vccd1 vccd1 _13205_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_151_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17608__B1 _17606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ _19323_/A vssd1 vssd1 vccd1 vccd1 _19512_/C sky130_fd_sc_hd__clkbuf_4
X_16920_ _14631_/X _16668_/B _16780_/B _23428_/Q vssd1 vssd1 vccd1 vccd1 _17133_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_172_1040 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1024 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16851_ _16849_/X _16850_/X _16836_/A vssd1 vssd1 vccd1 vccd1 _16853_/B sky130_fd_sc_hd__o21ai_1
XFILLER_120_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18820__A2 _19504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22299__B _22476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15802_ _15802_/A _15802_/B vssd1 vssd1 vccd1 vccd1 _15802_/Y sky130_fd_sc_hd__nand2_2
X_19570_ _19573_/A _19573_/B _19573_/C _19572_/A vssd1 vssd1 vccd1 vccd1 _19570_/X
+ sky130_fd_sc_hd__a31o_1
X_16782_ _17217_/A _17218_/A vssd1 vssd1 vccd1 vccd1 _17022_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12448__A2 _19040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13994_ _13994_/A _13994_/B vssd1 vssd1 vccd1 vccd1 _14791_/C sky130_fd_sc_hd__nand2_2
XFILLER_46_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18521_ _12465_/X _18501_/X _12463_/Y _18518_/A _18518_/B vssd1 vssd1 vccd1 vccd1
+ _18522_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_19_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _15860_/C vssd1 vssd1 vccd1 vccd1 _16526_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_92_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_61 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12945_ _12945_/A _12945_/B vssd1 vssd1 vccd1 vccd1 _12945_/Y sky130_fd_sc_hd__nand2_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _18452_/A vssd1 vssd1 vccd1 vccd1 _19803_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16595__B1 _16319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _15664_/A _23421_/Q _15664_/C _23423_/Q vssd1 vssd1 vccd1 vccd1 _16667_/B
+ sky130_fd_sc_hd__nor4_4
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12876_ _12876_/A vssd1 vssd1 vccd1 vccd1 _20908_/A sky130_fd_sc_hd__buf_2
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _17493_/C vssd1 vssd1 vccd1 vccd1 _17405_/C sky130_fd_sc_hd__inv_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _23297_/Q vssd1 vssd1 vccd1 vccd1 _14615_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_92_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18383_ _18383_/A _18383_/B vssd1 vssd1 vccd1 vccd1 _18384_/A sky130_fd_sc_hd__and2_1
XFILLER_159_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11827_ _18657_/C vssd1 vssd1 vccd1 vccd1 _16921_/C sky130_fd_sc_hd__clkbuf_4
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_820 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18336__A1 _18335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _23414_/Q _23415_/Q vssd1 vssd1 vccd1 vccd1 _15628_/A sky130_fd_sc_hd__nor2_1
XANTENNA__17139__A2 _12006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19533__B1 _18673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17334_ _17334_/A _17334_/B _17350_/B vssd1 vssd1 vccd1 vccd1 _17335_/B sky130_fd_sc_hd__nand3_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14546_ _14546_/A vssd1 vssd1 vccd1 vccd1 _14547_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11758_ _11758_/A vssd1 vssd1 vccd1 vccd1 _18814_/A sky130_fd_sc_hd__buf_2
XFILLER_187_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17265_ _16355_/A _12518_/X _17069_/A vssd1 vssd1 vccd1 vccd1 _17265_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_197_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12346__A _12346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14477_ _14472_/D _13985_/D _13972_/X _14462_/Y _14461_/X vssd1 vssd1 vccd1 vccd1
+ _14478_/B sky130_fd_sc_hd__a32o_1
X_11689_ _12282_/B _18999_/C _11665_/A vssd1 vssd1 vccd1 vccd1 _11689_/Y sky130_fd_sc_hd__a21oi_4
X_19004_ _11822_/X _19190_/A _19012_/A vssd1 vssd1 vccd1 vccd1 _19007_/A sky130_fd_sc_hd__o21ai_1
X_16216_ _15899_/X _15910_/X _15907_/B _15902_/Y vssd1 vssd1 vccd1 vccd1 _16216_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_13428_ _21924_/A _21923_/A vssd1 vssd1 vccd1 vccd1 _13444_/A sky130_fd_sc_hd__nand2_1
X_17196_ _16970_/Y _17028_/Y _17036_/X _17195_/Y vssd1 vssd1 vccd1 vccd1 _17196_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_115_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16147_ _16147_/A vssd1 vssd1 vccd1 vccd1 _17431_/A sky130_fd_sc_hd__buf_2
X_13359_ _23325_/Q _13358_/X _13264_/B _23326_/Q vssd1 vssd1 vccd1 vccd1 _13796_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_114_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17311__A2 _17305_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16078_ _16078_/A _16078_/B _16078_/C vssd1 vssd1 vccd1 vccd1 _16297_/A sky130_fd_sc_hd__nand3_2
XFILLER_142_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13177__A _13177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19906_ _19902_/Y _19904_/X _19909_/A vssd1 vssd1 vccd1 vccd1 _19928_/C sky130_fd_sc_hd__o21bai_2
XFILLER_102_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15029_ _15035_/A _15035_/B _15028_/Y vssd1 vssd1 vccd1 vccd1 _15033_/B sky130_fd_sc_hd__a21o_1
XFILLER_190_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17075__A1 _17565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19837_ _19835_/Y _19836_/Y _19833_/X _19939_/A vssd1 vssd1 vccd1 vccd1 _19874_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_111_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23148__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16822__A1 _15749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16822__B2 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19768_ _19768_/A _19928_/A _19928_/B vssd1 vssd1 vccd1 vccd1 _19768_/Y sky130_fd_sc_hd__nand3_2
Xinput2 wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13636__A1 _21921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_620 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18719_ _18902_/B vssd1 vssd1 vccd1 vccd1 _18914_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__19799__A _19966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19699_ _19547_/X _19537_/X _19538_/X _19542_/X vssd1 vssd1 vccd1 vccd1 _19831_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21730_ _21722_/B _21728_/A _23578_/Q vssd1 vssd1 vccd1 vccd1 _21730_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17783__C1 _17771_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19949__D _19949_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16050__A2 _17226_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23114__A _23182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21661_ _21654_/A _21654_/B _23572_/Q vssd1 vssd1 vccd1 vccd1 _21661_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14736__A _23595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18208__A _18208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23400_ _23433_/CLK _23400_/D vssd1 vssd1 vccd1 vccd1 _23400_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17112__A _17112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20612_ _20612_/A vssd1 vssd1 vccd1 vccd1 _21414_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21592_ _21592_/A _21592_/B _21554_/D vssd1 vssd1 vccd1 vccd1 _21594_/A sky130_fd_sc_hd__nor3b_1
XFILLER_32_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23331_ _23332_/CLK _23331_/D vssd1 vssd1 vccd1 vccd1 _23331_/Q sky130_fd_sc_hd__dfxtp_2
X_20543_ _13054_/Y _13184_/A _20966_/C _13058_/Y vssd1 vssd1 vccd1 vccd1 _20553_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17550__A2 _17303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23262_ _23584_/CLK _23262_/D vssd1 vssd1 vccd1 vccd1 _23262_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17766__B _17766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20474_ _12871_/A _12872_/A _20620_/C _12876_/A vssd1 vssd1 vccd1 vccd1 _20475_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_193_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12375__A1 _19082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12375__B2 _19082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22213_ _22290_/B _22166_/Y _22290_/A vssd1 vssd1 vccd1 vccd1 _22214_/B sky130_fd_sc_hd__a21o_1
XFILLER_192_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1040 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23193_ _15762_/A input32/X _23195_/S vssd1 vssd1 vccd1 vccd1 _23194_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22144_ _22144_/A _22168_/A _22144_/C _22144_/D vssd1 vssd1 vccd1 vccd1 _22268_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_161_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13324__B1 _13253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22075_ _22203_/A _22203_/B _22069_/Y _22074_/X vssd1 vssd1 vccd1 vccd1 _22075_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20407__A_N _20408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__C _18511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21026_ _21026_/A _21031_/B vssd1 vssd1 vccd1 vccd1 _21028_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23139__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22977_ _13253_/A input32/X _22979_/S vssd1 vssd1 vccd1 vccd1 _22978_/A sky130_fd_sc_hd__mux2_1
XANTENNA__21165__A3 _20966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19502__A _19502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _12723_/X _12725_/X _12728_/Y vssd1 vssd1 vccd1 vccd1 _12733_/A sky130_fd_sc_hd__o21ai_1
XFILLER_128_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21928_ _22172_/C _22292_/A _22293_/A _22548_/A _21921_/C vssd1 vssd1 vccd1 vccd1
+ _21928_/X sky130_fd_sc_hd__a32o_2
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12661_/A _12661_/B vssd1 vssd1 vccd1 vccd1 _12662_/C sky130_fd_sc_hd__nand2_1
XFILLER_188_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _21859_/A _21859_/B vssd1 vssd1 vccd1 vccd1 _22107_/A sky130_fd_sc_hd__nand2_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _12260_/C vssd1 vssd1 vccd1 vccd1 _12308_/A sky130_fd_sc_hd__buf_2
X_14400_ _14400_/A _14400_/B _14400_/C vssd1 vssd1 vccd1 vccd1 _14442_/B sky130_fd_sc_hd__nand3_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _15380_/A _15380_/B vssd1 vssd1 vccd1 vccd1 _15382_/C sky130_fd_sc_hd__nand2_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12592_ _12606_/A _12606_/C _13011_/C vssd1 vssd1 vccd1 vccd1 _12601_/A sky130_fd_sc_hd__nand3_4
XFILLER_168_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18869__A2 _18627_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14331_ _14331_/A _14384_/A _14331_/C vssd1 vssd1 vccd1 vccd1 _14395_/A sky130_fd_sc_hd__nand3_1
X_23529_ _23558_/CLK _23529_/D vssd1 vssd1 vccd1 vccd1 _23529_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17050_ _17050_/A vssd1 vssd1 vccd1 vccd1 _17050_/X sky130_fd_sc_hd__clkbuf_2
X_14262_ _14262_/A vssd1 vssd1 vccd1 vccd1 _14886_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_184_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20383__A _20411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13213_ _13213_/A vssd1 vssd1 vccd1 vccd1 _23539_/D sky130_fd_sc_hd__clkbuf_1
X_16001_ _16010_/A _16000_/Y _15878_/X _15879_/Y vssd1 vssd1 vccd1 vccd1 _16249_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_183_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14193_ _14193_/A _14193_/B _14193_/C _14193_/D vssd1 vssd1 vccd1 vccd1 _14194_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_48_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15304__A1 _15358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13144_ _13143_/C _13143_/B _13143_/A vssd1 vssd1 vccd1 vccd1 _13196_/A sky130_fd_sc_hd__a21o_1
XFILLER_151_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16501__B1 _16536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15304__B2 _15415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18788__A _18788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17952_ _18148_/A _18148_/B _17952_/C vssd1 vssd1 vccd1 vccd1 _17954_/C sky130_fd_sc_hd__and3_1
X_13075_ _13089_/B _13089_/C vssd1 vssd1 vccd1 vccd1 _13075_/Y sky130_fd_sc_hd__nand2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16903_ _15918_/C _15610_/X _16365_/A _15682_/A _15660_/A vssd1 vssd1 vccd1 vccd1
+ _17140_/A sky130_fd_sc_hd__o2111ai_4
X_12026_ _12022_/X _12025_/X _12029_/B _12011_/X vssd1 vssd1 vccd1 vccd1 _12026_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__11877__B1 _12373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17883_ _19957_/A vssd1 vssd1 vccd1 vccd1 _18016_/C sky130_fd_sc_hd__buf_2
X_19622_ _19932_/A _19620_/X _19621_/X _19380_/X vssd1 vssd1 vccd1 vccd1 _19627_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16834_ _15861_/X _16058_/A _16841_/A vssd1 vssd1 vccd1 vccd1 _16834_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_120_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18006__B1 _20081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19553_ _19533_/X _19534_/X _19546_/Y _19552_/Y vssd1 vssd1 vccd1 vccd1 _19562_/B
+ sky130_fd_sc_hd__o211ai_1
X_16765_ _16765_/A vssd1 vssd1 vccd1 vccd1 _17009_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13977_ _13977_/A _13977_/B vssd1 vssd1 vccd1 vccd1 _13978_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16754__A1_N _16988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18504_ _12173_/X _12174_/X _18503_/C _12175_/X _18503_/D vssd1 vssd1 vccd1 vccd1
+ _18504_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_0_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_612 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15716_ _15713_/C _15716_/B _15716_/C vssd1 vssd1 vccd1 vccd1 _16856_/D sky130_fd_sc_hd__nand3b_4
X_19484_ _19670_/C _19480_/A _19482_/Y vssd1 vssd1 vccd1 vccd1 _19486_/A sky130_fd_sc_hd__o21ai_1
XFILLER_20_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _13179_/A _13116_/C _13156_/A _21182_/D vssd1 vssd1 vccd1 vccd1 _13113_/A
+ sky130_fd_sc_hd__nand4_1
X_16696_ _16135_/B _16135_/C _16135_/A vssd1 vssd1 vccd1 vccd1 _16696_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18435_ _18435_/A _18435_/B vssd1 vssd1 vccd1 vccd1 _19280_/A sky130_fd_sc_hd__nor2_2
XANTENNA__22476__C _22476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_678 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15647_ _15647_/A _15647_/B vssd1 vssd1 vccd1 vccd1 _17098_/B sky130_fd_sc_hd__nor2_4
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12859_ _12859_/A _12859_/B _12859_/C vssd1 vssd1 vccd1 vccd1 _12860_/A sky130_fd_sc_hd__nand3_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19506__B1 _12040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18366_ _18363_/Y _18364_/Y _18264_/C _18264_/A vssd1 vssd1 vccd1 vccd1 _18366_/Y
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__13251__C1 _13253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15578_ _15585_/D _23511_/Q _15586_/C vssd1 vssd1 vccd1 vccd1 _15580_/A sky130_fd_sc_hd__and3_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17317_ _16054_/X _16055_/X _17029_/X _16665_/X _17722_/A vssd1 vssd1 vccd1 vccd1
+ _17318_/B sky130_fd_sc_hd__o221a_1
X_14529_ _14538_/B _14538_/C _14535_/A input2/X vssd1 vssd1 vccd1 vccd1 _22968_/D
+ sky130_fd_sc_hd__and4bb_2
XFILLER_30_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18297_ _18305_/A _18305_/B _18295_/X _18296_/X vssd1 vssd1 vccd1 vccd1 _18297_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_187_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12076__A _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15138__A4 _15408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23526__CLK _23538_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17248_ _17449_/A _17450_/B _17248_/C _20317_/C vssd1 vssd1 vccd1 vccd1 _17248_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_31_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19809__A1 _17610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16490__B _17974_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21077__C1 _21271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17179_ _17179_/A _17179_/B _17179_/C vssd1 vssd1 vccd1 vccd1 _17179_/X sky130_fd_sc_hd__and3_1
XFILLER_115_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18493__B1 _18458_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21092__A2 _20984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20190_ _20184_/A _20184_/B _20186_/B vssd1 vssd1 vccd1 vccd1 _20190_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_116_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15846__A2 _15975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17048__A1 _15884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22900_ _22900_/A vssd1 vssd1 vccd1 vccd1 _23286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21852__A _21852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22831_ _22830_/B _22830_/C _22759_/A vssd1 vssd1 vccd1 vccd1 _22861_/A sky130_fd_sc_hd__o21ai_1
XFILLER_186_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22762_ _22762_/A _22762_/B vssd1 vssd1 vccd1 vccd1 _22763_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_740 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21713_ _21705_/X _21679_/X _21712_/Y vssd1 vssd1 vccd1 vccd1 _21715_/A sky130_fd_sc_hd__a21oi_1
XFILLER_25_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22693_ _22818_/A _22694_/B _22694_/C vssd1 vssd1 vccd1 vccd1 _22695_/A sky130_fd_sc_hd__a21oi_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21644_ _21645_/A _21645_/B _21645_/C vssd1 vssd1 vccd1 vccd1 _21646_/A sky130_fd_sc_hd__o21a_2
XANTENNA__12045__B1 _19512_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21855__A1 _21842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20658__A2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21575_ _21474_/B _21574_/Y _21577_/B vssd1 vssd1 vccd1 vccd1 _21575_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_193_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_642 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23314_ _23378_/CLK _23314_/D vssd1 vssd1 vccd1 vccd1 _23314_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12417__C _18788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15534__A1 _15225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20526_ _12765_/A _12936_/A _12952_/X _13025_/X vssd1 vssd1 vccd1 vccd1 _20526_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23245_ _23245_/A vssd1 vssd1 vccd1 vccd1 _23440_/D sky130_fd_sc_hd__clkbuf_1
X_20457_ _20457_/A _20457_/B vssd1 vssd1 vccd1 vccd1 _23538_/D sky130_fd_sc_hd__nor2_1
XFILLER_106_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20815__C1 _21065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23176_ _23410_/Q input27/X _23178_/S vssd1 vssd1 vccd1 vccd1 _23177_/A sky130_fd_sc_hd__mux2_1
X_20388_ _20362_/Y _20415_/B _20415_/A vssd1 vssd1 vccd1 vccd1 _20392_/A sky130_fd_sc_hd__nand3b_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22127_ _22365_/C vssd1 vssd1 vccd1 vccd1 _22647_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__19028__A2 _11951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20830__A2 _12648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22568__C1 _22392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22058_ _22057_/X _22168_/A _22033_/A vssd1 vssd1 vccd1 vccd1 _22377_/A sky130_fd_sc_hd__o21ai_1
XFILLER_153_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21009_ _20597_/C _21007_/Y _21008_/X _21157_/C _21157_/D vssd1 vssd1 vccd1 vccd1
+ _21011_/B sky130_fd_sc_hd__o311a_1
X_13900_ _14188_/C _14011_/B vssd1 vssd1 vccd1 vccd1 _13966_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14880_ _14889_/A _14889_/B _14114_/X vssd1 vssd1 vccd1 vccd1 _14893_/A sky130_fd_sc_hd__a21o_1
XANTENNA__22858__A _22858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13831_ _13799_/X _13813_/X _21786_/A _21786_/B vssd1 vssd1 vccd1 vccd1 _13834_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_910 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16550_ _16548_/X _16528_/B _16526_/C _16549_/X vssd1 vssd1 vccd1 vccd1 _16554_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_44_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19200__A2 _19196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13762_ _21856_/D _21856_/C vssd1 vssd1 vccd1 vccd1 _13763_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12284__B1 _15699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _15501_/A _15501_/B _15501_/C vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__and3_1
X_12713_ _12644_/X _12601_/C _12712_/X vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__a21oi_1
X_16481_ _12379_/X _16451_/B _16451_/C _16479_/X _16480_/X vssd1 vssd1 vccd1 vccd1
+ _16481_/X sky130_fd_sc_hd__o32a_1
XFILLER_15_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13693_ _13692_/A _13692_/B _13691_/B _21839_/B vssd1 vssd1 vccd1 vccd1 _13760_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18220_ _18279_/A _18279_/B _20317_/A _18279_/D vssd1 vssd1 vccd1 vccd1 _18220_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_102_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13280__A _13766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15432_ _15433_/B _15433_/A vssd1 vssd1 vccd1 vccd1 _15432_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12644_ _12688_/A vssd1 vssd1 vccd1 vccd1 _12644_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18151_ _17952_/C _18144_/Y _18149_/Y _18150_/X vssd1 vssd1 vccd1 vccd1 _18262_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_156_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17499__A1_N _17154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15363_ _15363_/A _15363_/B _15363_/C _15363_/D vssd1 vssd1 vccd1 vccd1 _15366_/D
+ sky130_fd_sc_hd__and4_1
X_12575_ _20493_/B _23287_/Q _23286_/Q vssd1 vssd1 vccd1 vccd1 _12874_/D sky130_fd_sc_hd__nor3_2
XFILLER_12_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16591__A _16591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17102_ _16856_/Y _17093_/Y _17096_/A vssd1 vssd1 vccd1 vccd1 _17104_/A sky130_fd_sc_hd__o21ai_1
X_14314_ _14097_/A _13964_/Y _14207_/Y vssd1 vssd1 vccd1 vccd1 _14355_/C sky130_fd_sc_hd__o21ai_1
X_18082_ _20215_/A vssd1 vssd1 vccd1 vccd1 _20271_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15294_ _15294_/A _15294_/B vssd1 vssd1 vccd1 vccd1 _15331_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17033_ _17891_/A vssd1 vssd1 vccd1 vccd1 _18163_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_156_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14245_ _14245_/A _14245_/B vssd1 vssd1 vccd1 vccd1 _14245_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14176_ _14178_/B _14276_/A _14178_/A vssd1 vssd1 vccd1 vccd1 _14177_/B sky130_fd_sc_hd__and3_1
XANTENNA_output89_A _23263_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13127_ _13172_/C _13172_/A vssd1 vssd1 vccd1 vccd1 _13128_/B sky130_fd_sc_hd__nand2_1
XANTENNA__20821__A2 _12850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _18984_/A _18984_/B vssd1 vssd1 vccd1 vccd1 _18984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23574__D _23574_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23220__A0 _16780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22023__A1 _21902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17935_ _18058_/D _18072_/D _18072_/C _17935_/D vssd1 vssd1 vccd1 vccd1 _18198_/C
+ sky130_fd_sc_hd__nand4_4
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13058_ _13058_/A _13058_/B vssd1 vssd1 vccd1 vccd1 _13058_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater105 _23332_/CLK vssd1 vssd1 vccd1 vccd1 _23429_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13455__A _22035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater116 _23428_/CLK vssd1 vssd1 vccd1 vccd1 _23425_/CLK sky130_fd_sc_hd__clkbuf_1
X_12009_ _12024_/A _12024_/B _18973_/C vssd1 vssd1 vccd1 vccd1 _12010_/B sky130_fd_sc_hd__nand3_2
Xrepeater127 _23336_/CLK vssd1 vssd1 vccd1 vccd1 _23445_/CLK sky130_fd_sc_hd__clkbuf_1
X_17866_ _12088_/A _16742_/A _17860_/Y _17859_/Y _18013_/A vssd1 vssd1 vccd1 vccd1
+ _17880_/B sky130_fd_sc_hd__o221ai_4
Xrepeater138 _23434_/CLK vssd1 vssd1 vccd1 vccd1 _23402_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater149 _23401_/CLK vssd1 vssd1 vccd1 vccd1 _23309_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_93_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19605_ _19605_/A _19605_/B _19605_/C vssd1 vssd1 vccd1 vccd1 _19764_/A sky130_fd_sc_hd__nand3_2
X_16817_ _16817_/A vssd1 vssd1 vccd1 vccd1 _17050_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15056__A3 _14933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17797_ _17779_/Y _17786_/Y _17796_/Y vssd1 vssd1 vccd1 vccd1 _17801_/B sky130_fd_sc_hd__a21o_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19536_ _17591_/A _17593_/A _19539_/B _19539_/A _17595_/A vssd1 vssd1 vccd1 vccd1
+ _19701_/A sky130_fd_sc_hd__o2111ai_2
XFILLER_81_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16748_ _18279_/B vssd1 vssd1 vccd1 vccd1 _18157_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12814__A2 _12785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19467_ _19467_/A vssd1 vssd1 vccd1 vccd1 _19625_/A sky130_fd_sc_hd__buf_2
XFILLER_59_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16679_ _15644_/X _16657_/B _15639_/C _15791_/A vssd1 vssd1 vccd1 vccd1 _16679_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18418_ _18417_/B _18417_/C _18154_/X _18399_/Y vssd1 vssd1 vccd1 vccd1 _18420_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23599__A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19398_ _19401_/A _19398_/B _19402_/A _19402_/B vssd1 vssd1 vccd1 vccd1 _19399_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18349_ _18349_/A _18349_/B _18349_/C vssd1 vssd1 vccd1 vccd1 _18350_/A sky130_fd_sc_hd__nand3_1
XFILLER_159_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12042__A3 _18941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20104__A4 _20369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21360_ _21292_/Y _21433_/A _21359_/Y vssd1 vssd1 vccd1 vccd1 _21360_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__14319__A2 _15356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20311_ _20311_/A _20311_/B vssd1 vssd1 vccd1 vccd1 _20312_/C sky130_fd_sc_hd__nand2_1
XFILLER_147_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21291_ _20502_/X _20504_/X _21430_/C _21431_/A vssd1 vssd1 vccd1 vccd1 _21359_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17269__A1 _16638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23030_ _23345_/Q input26/X _23034_/S vssd1 vssd1 vccd1 vccd1 _23031_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14452__C _15310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20242_ _20290_/B _20242_/B vssd1 vssd1 vccd1 vccd1 _20243_/A sky130_fd_sc_hd__and2_1
XANTENNA__22262__A1 _21829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18466__B1 _18997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22801__A3 _22861_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15845__A _16634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20173_ _20170_/Y _20171_/X _20176_/A vssd1 vssd1 vccd1 vccd1 _20173_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__19317__A _19320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18859__C _18859_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18221__A _20210_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23484__D _23496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15295__A3 _14061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23211__A0 _15921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20901__D _23300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21285__C _21285_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18769__A1 _11815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17441__A1 _16479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22814_ _21850_/A _21850_/B _22828_/A _22828_/B vssd1 vssd1 vccd1 vccd1 _22815_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19194__A1 _11936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22745_ _22745_/A _22818_/C vssd1 vssd1 vccd1 vccd1 _22821_/C sky130_fd_sc_hd__nand2_1
XFILLER_53_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12709__A _12709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11613__A _19662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22676_ _22676_/A _22676_/B _22720_/B _22676_/D vssd1 vssd1 vccd1 vccd1 _22676_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21627_ _21540_/A _21627_/B _21627_/C _21627_/D vssd1 vssd1 vccd1 vccd1 _21627_/Y
+ sky130_fd_sc_hd__nand4b_1
XFILLER_194_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11777__C1 _11634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12360_ _12360_/A _12360_/B _12381_/C _12381_/B vssd1 vssd1 vccd1 vccd1 _12360_/Y
+ sky130_fd_sc_hd__nand4_1
X_21558_ _21510_/C _21507_/B _21559_/C _21509_/A _21557_/Y vssd1 vssd1 vccd1 vccd1
+ _21564_/B sky130_fd_sc_hd__o221ai_2
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20509_ _20509_/A _20509_/B vssd1 vssd1 vccd1 vccd1 _20509_/Y sky130_fd_sc_hd__nor2_1
X_12291_ _12547_/B _12291_/B vssd1 vssd1 vccd1 vccd1 _12364_/C sky130_fd_sc_hd__nor2_1
XFILLER_107_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21489_ _21407_/A _21407_/B _21488_/X _21474_/B vssd1 vssd1 vccd1 vccd1 _21524_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_5_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14030_ _23498_/Q vssd1 vssd1 vccd1 vccd1 _14429_/A sky130_fd_sc_hd__buf_2
XFILLER_180_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23228_ _23433_/Q input17/X _23228_/S vssd1 vssd1 vccd1 vccd1 _23229_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18457__B1 _19969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20264__B1 _18001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23159_ _23402_/Q input19/X _23167_/S vssd1 vssd1 vccd1 vccd1 _23160_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input40_A wb_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23202__A0 _15713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15981_ _16668_/C _15693_/Y _15694_/Y _12207_/A vssd1 vssd1 vccd1 vccd1 _15982_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17720_ _12237_/A _17506_/A _17628_/Y _17712_/Y _17899_/A vssd1 vssd1 vccd1 vccd1
+ _17720_/Y sky130_fd_sc_hd__o221ai_1
XANTENNA__13275__A _13498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14932_ _14943_/A _14943_/B _14966_/B vssd1 vssd1 vccd1 vccd1 _14932_/X sky130_fd_sc_hd__and3_1
XANTENNA__21055__A1_N _21054_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17432__A1 _16370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1012 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17651_ _17657_/A _17656_/C vssd1 vssd1 vccd1 vccd1 _17653_/B sky130_fd_sc_hd__nand2_1
X_14863_ _14863_/A _23352_/Q _14863_/C _14863_/D vssd1 vssd1 vccd1 vccd1 _14868_/D
+ sky130_fd_sc_hd__nor4_4
XFILLER_48_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20972__D1 _12980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16602_ _16598_/Y _16599_/Y _16600_/Y _16601_/Y vssd1 vssd1 vccd1 vccd1 _16608_/A
+ sky130_fd_sc_hd__o211ai_2
X_13814_ _21923_/A _13814_/B _21924_/A vssd1 vssd1 vccd1 vccd1 _13814_/Y sky130_fd_sc_hd__nand3_1
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17582_ _17845_/D _18778_/A _18778_/B vssd1 vssd1 vccd1 vccd1 _17583_/B sky130_fd_sc_hd__and3_1
XFILLER_21_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14794_ _13969_/Y _15084_/A _14791_/Y _14793_/Y vssd1 vssd1 vccd1 vccd1 _14934_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__15921__C _15921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19185__A1 _16360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15994__B2 _15969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19321_ _19321_/A vssd1 vssd1 vccd1 vccd1 _19524_/A sky130_fd_sc_hd__buf_2
X_16533_ _16483_/Y _16518_/C _16512_/Y vssd1 vssd1 vccd1 vccd1 _16533_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13745_ _13739_/A _13739_/B _13739_/C _22465_/D _13743_/A vssd1 vssd1 vccd1 vccd1
+ _13745_/Y sky130_fd_sc_hd__o311ai_1
XFILLER_31_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19252_ _19434_/A _19434_/B _19434_/C vssd1 vssd1 vccd1 vccd1 _19297_/A sky130_fd_sc_hd__nand3_2
XFILLER_43_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16464_ _16464_/A vssd1 vssd1 vccd1 vccd1 _16464_/X sky130_fd_sc_hd__clkbuf_8
X_13676_ _13676_/A _13676_/B _13676_/C vssd1 vssd1 vccd1 vccd1 _13692_/A sky130_fd_sc_hd__nand3_1
X_18203_ _18154_/X _18302_/C _18302_/A vssd1 vssd1 vccd1 vccd1 _18204_/C sky130_fd_sc_hd__o21ai_1
XFILLER_148_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15415_ _15415_/A vssd1 vssd1 vccd1 vccd1 _15446_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_19183_ _19325_/A _19183_/B _19183_/C vssd1 vssd1 vccd1 vccd1 _19188_/B sky130_fd_sc_hd__nand3_1
X_12627_ _12622_/X _12624_/X _12932_/A vssd1 vssd1 vccd1 vccd1 _12627_/X sky130_fd_sc_hd__a21o_2
X_16395_ _16395_/A _16395_/B _16395_/C vssd1 vssd1 vccd1 vccd1 _16396_/A sky130_fd_sc_hd__nand3_1
XANTENNA__14834__A _14834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23569__D _23569_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18134_ _18134_/A _18134_/B _18134_/C vssd1 vssd1 vccd1 vccd1 _18155_/B sky130_fd_sc_hd__and3_1
XFILLER_157_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15346_ _15294_/A _15294_/B _15331_/B vssd1 vssd1 vccd1 vccd1 _15391_/A sky130_fd_sc_hd__a21oi_2
X_12558_ _12565_/C _12565_/B _12561_/A _19089_/B vssd1 vssd1 vccd1 vccd1 _12558_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18065_ _18144_/C _18149_/B _18066_/C vssd1 vssd1 vccd1 vccd1 _18067_/A sky130_fd_sc_hd__a21oi_1
XFILLER_171_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15277_ _15277_/A _15277_/B _15277_/C vssd1 vssd1 vccd1 vccd1 _15279_/A sky130_fd_sc_hd__nand3_1
X_12489_ _12478_/A _12478_/B _12478_/C vssd1 vssd1 vccd1 vccd1 _18524_/A sky130_fd_sc_hd__a21o_1
XFILLER_89_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17016_ _17003_/Y _17014_/Y _17015_/Y vssd1 vssd1 vccd1 vccd1 _17018_/A sky130_fd_sc_hd__a21oi_1
XFILLER_176_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14228_ _14228_/A _14228_/B vssd1 vssd1 vccd1 vccd1 _14229_/D sky130_fd_sc_hd__nand2_1
XANTENNA__19645__C1 _19502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _14790_/B _14795_/A _14795_/B _14396_/A _14796_/B vssd1 vssd1 vccd1 vccd1
+ _14167_/A sky130_fd_sc_hd__a32o_1
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20290__B _20290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ _18969_/A _18969_/B vssd1 vssd1 vccd1 vccd1 _19246_/A sky130_fd_sc_hd__nand2_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_523 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17918_ _17919_/A _17919_/B _17919_/C _17919_/D vssd1 vssd1 vccd1 vccd1 _17920_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12496__B1 _12211_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18898_ _18717_/C _18717_/A _18717_/B _18902_/A _18914_/C vssd1 vssd1 vccd1 vccd1
+ _18899_/C sky130_fd_sc_hd__a32oi_1
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17849_ _17742_/X _17741_/X _17605_/A _17581_/A _17605_/B vssd1 vssd1 vccd1 vccd1
+ _17982_/B sky130_fd_sc_hd__o2111a_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14237__A1 _14230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20860_ _20860_/A vssd1 vssd1 vccd1 vccd1 _20885_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19519_ _19575_/A _19575_/B _19519_/C _19519_/D vssd1 vssd1 vccd1 vccd1 _19519_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17104__B _17104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20791_ _12633_/A _20786_/Y _20778_/X _20920_/A _20783_/Y vssd1 vssd1 vccd1 vccd1
+ _20794_/B sky130_fd_sc_hd__o221ai_1
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22530_ _22530_/A vssd1 vssd1 vccd1 vccd1 _22530_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_732 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15737__A1 _15864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19957__D _19957_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_607 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22461_ _22461_/A vssd1 vssd1 vccd1 vccd1 _22461_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19479__A2 _18484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21412_ _23567_/Q vssd1 vssd1 vccd1 vccd1 _21418_/A sky130_fd_sc_hd__inv_2
X_22392_ _22392_/A _22392_/B _22392_/C vssd1 vssd1 vccd1 vccd1 _22393_/B sky130_fd_sc_hd__and3_1
XANTENNA__15559__B _15559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12971__A1 _12979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21343_ _21264_/Y _21240_/A _21342_/C vssd1 vssd1 vccd1 vccd1 _21343_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_194_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12264__A _16049_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21274_ _21274_/A _21397_/A _21274_/C vssd1 vssd1 vccd1 vccd1 _21327_/B sky130_fd_sc_hd__nand3_1
XFILLER_118_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23013_ _23013_/A vssd1 vssd1 vccd1 vccd1 _23337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20225_ _18001_/X _20164_/B _20263_/A _20223_/Y _20221_/X vssd1 vssd1 vccd1 vccd1
+ _20225_/X sky130_fd_sc_hd__o311a_1
XANTENNA__16465__A2 _16447_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20156_ _20158_/A _20156_/B vssd1 vssd1 vccd1 vccd1 _20156_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14476__A1 _15044_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13095__A _21490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_67 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20087_ _20095_/A _20172_/B _20095_/C vssd1 vssd1 vccd1 vccd1 _20087_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_58_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_707 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15976__A1 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11860_ _11860_/A _11860_/B _11860_/C vssd1 vssd1 vccd1 vccd1 _12019_/A sky130_fd_sc_hd__and3_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15976__B2 _16123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11791_ _23584_/Q _11644_/C _11808_/A _11741_/A vssd1 vssd1 vccd1 vccd1 _11792_/B
+ sky130_fd_sc_hd__o211ai_4
X_20989_ _20989_/A _20989_/B vssd1 vssd1 vccd1 vccd1 _20994_/A sky130_fd_sc_hd__nor2_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22171__B1 _22381_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13530_ _21921_/C vssd1 vssd1 vccd1 vccd1 _22278_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_53_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_704 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22728_ _22750_/A _22750_/B vssd1 vssd1 vccd1 vccd1 _22731_/A sky130_fd_sc_hd__xnor2_1
XFILLER_43_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13461_ _13461_/A _13461_/B _13461_/C vssd1 vssd1 vccd1 vccd1 _13462_/A sky130_fd_sc_hd__nand3_1
XANTENNA__14654__A _21853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22659_ _22661_/B _22710_/A _22556_/X _22658_/Y vssd1 vssd1 vccd1 vccd1 _22671_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15200_ _15196_/X _15197_/X _15199_/Y vssd1 vssd1 vccd1 vccd1 _15201_/B sky130_fd_sc_hd__o21a_1
X_12412_ _12410_/Y _12100_/C _18997_/A vssd1 vssd1 vccd1 vccd1 _12413_/A sky130_fd_sc_hd__a21oi_2
XFILLER_167_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16180_ _15985_/A _15985_/B _15985_/C vssd1 vssd1 vccd1 vccd1 _16180_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_139_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13392_ _13392_/A _13392_/B vssd1 vssd1 vccd1 vccd1 _21764_/B sky130_fd_sc_hd__nand2_2
XFILLER_166_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15131_ _15035_/B _15028_/Y _15035_/A vssd1 vssd1 vccd1 vccd1 _15132_/C sky130_fd_sc_hd__a21boi_1
X_12343_ _12343_/A vssd1 vssd1 vccd1 vccd1 _19530_/A sky130_fd_sc_hd__buf_2
XFILLER_138_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12274_ _12266_/Y _12339_/C _12295_/A vssd1 vssd1 vccd1 vccd1 _12288_/A sky130_fd_sc_hd__o21a_1
X_15062_ _15067_/B _15067_/C _15067_/A vssd1 vssd1 vccd1 vccd1 _15063_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__15900__A1 _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14013_ _14193_/A _14013_/B _14027_/A _14023_/C vssd1 vssd1 vccd1 vccd1 _14017_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_153_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19870_ _20269_/C _19864_/B _17546_/C _19655_/X vssd1 vssd1 vccd1 vccd1 _19870_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_134_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18821_ _11654_/A _12424_/A _18820_/Y vssd1 vssd1 vccd1 vccd1 _19029_/A sky130_fd_sc_hd__o21ai_4
XFILLER_110_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18752_ _18714_/Y _18715_/X _18892_/A vssd1 vssd1 vccd1 vccd1 _18752_/X sky130_fd_sc_hd__o21a_1
X_15964_ _17060_/A _15964_/B _17061_/A vssd1 vssd1 vccd1 vccd1 _15964_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17703_ _17703_/A _17703_/B _17703_/C vssd1 vssd1 vccd1 vccd1 _18253_/B sky130_fd_sc_hd__nand3_2
XANTENNA__18602__B1 _17761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14915_ _14588_/X _14050_/X _14061_/X _14901_/X _14448_/A vssd1 vssd1 vccd1 vccd1
+ _14915_/X sky130_fd_sc_hd__o311a_1
X_18683_ _18474_/X _19491_/A _18481_/X _18473_/X vssd1 vssd1 vccd1 vccd1 _18687_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_49_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15895_ _15895_/A _16022_/A _15895_/C vssd1 vssd1 vccd1 vccd1 _16078_/C sky130_fd_sc_hd__nand3_1
XANTENNA__13690__A2 _22713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17634_ _17634_/A _17634_/B vssd1 vssd1 vccd1 vccd1 _17637_/B sky130_fd_sc_hd__nand2_1
X_14846_ _14846_/A _14846_/B vssd1 vssd1 vccd1 vccd1 _14846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19123__C _19123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17565_ _17565_/A vssd1 vssd1 vccd1 vccd1 _17565_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14777_ _14777_/A _14777_/B _14777_/C vssd1 vssd1 vccd1 vccd1 _14778_/B sky130_fd_sc_hd__and3_1
XFILLER_56_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11989_ _18468_/A vssd1 vssd1 vccd1 vccd1 _12121_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_182_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19304_ _19304_/A vssd1 vssd1 vccd1 vccd1 _19304_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_90_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16516_ _16394_/A _16517_/C _16415_/B vssd1 vssd1 vccd1 vccd1 _16518_/A sky130_fd_sc_hd__a21bo_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13728_ _13723_/C _13723_/B _13717_/Y vssd1 vssd1 vccd1 vccd1 _13728_/X sky130_fd_sc_hd__a21bo_1
XFILLER_147_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17496_ _17337_/C _17386_/X _17337_/B vssd1 vssd1 vccd1 vccd1 _17498_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__16916__B1 _12051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19235_ _19256_/B _19256_/C _19256_/A vssd1 vssd1 vccd1 vccd1 _19257_/B sky130_fd_sc_hd__a21o_1
XFILLER_149_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16447_ _16447_/A _16447_/B vssd1 vssd1 vccd1 vccd1 _16447_/Y sky130_fd_sc_hd__nor2_4
X_13659_ _13659_/A _13659_/B vssd1 vssd1 vccd1 vccd1 _13659_/Y sky130_fd_sc_hd__nand2_2
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19166_ _12052_/A _19838_/A _19184_/A _19165_/Y _19158_/Y vssd1 vssd1 vccd1 vccd1
+ _19167_/C sky130_fd_sc_hd__o221ai_4
X_16378_ _16374_/A _16457_/B _16377_/X _16225_/X vssd1 vssd1 vccd1 vccd1 _16379_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_9_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23267__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19330__A1 _17408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18117_ _18298_/A _18298_/B vssd1 vssd1 vccd1 vccd1 _18119_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15329_ _15329_/A _15328_/Y vssd1 vssd1 vccd1 vccd1 _15330_/B sky130_fd_sc_hd__or2b_1
X_19097_ _19088_/B _19088_/C _19091_/C vssd1 vssd1 vccd1 vccd1 _19443_/B sky130_fd_sc_hd__a21boi_4
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18048_ _18129_/A vssd1 vssd1 vccd1 vccd1 _18049_/B sky130_fd_sc_hd__inv_2
XANTENNA__17892__B2 _17303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20010_ _20011_/A _20011_/B _19940_/X _19939_/Y vssd1 vssd1 vccd1 vccd1 _20012_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13627__B _22269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19999_ _19963_/A _19963_/B _19997_/Y _19998_/X vssd1 vssd1 vccd1 vccd1 _20003_/D
+ sky130_fd_sc_hd__o22ai_2
XFILLER_115_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19017__D _19017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1019 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13130__A1 _21121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15842__B _16591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15670__A3 _15655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21961_ _21965_/A _21961_/B _21961_/C vssd1 vssd1 vccd1 vccd1 _22118_/A sky130_fd_sc_hd__nand3b_2
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20912_ _21174_/A vssd1 vssd1 vccd1 vccd1 _21370_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_21892_ _21892_/A vssd1 vssd1 vccd1 vccd1 _21892_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _20843_/A _20843_/B vssd1 vssd1 vccd1 vccd1 _20843_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16376__D _16497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23562_ _23566_/CLK _23562_/D vssd1 vssd1 vccd1 vccd1 _23562_/Q sky130_fd_sc_hd__dfxtp_1
X_20774_ _20773_/D _20773_/A _20773_/C _20773_/B vssd1 vssd1 vccd1 vccd1 _20775_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22513_ _22513_/A _22513_/B _22513_/C vssd1 vssd1 vccd1 vccd1 _22516_/C sky130_fd_sc_hd__nand3_1
XANTENNA__16383__A1 _16225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23493_ _23518_/CLK _23505_/Q vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfxtp_1
XFILLER_196_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22444_ _22247_/Y _22348_/Y _22349_/Y _22443_/Y _22617_/A vssd1 vssd1 vccd1 vccd1
+ _22447_/A sky130_fd_sc_hd__o311a_1
XFILLER_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15289__B _15402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12944__A1 _12709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22375_ _22409_/A _22504_/A _22504_/B vssd1 vssd1 vccd1 vccd1 _22400_/A sky130_fd_sc_hd__a21o_1
XFILLER_136_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21326_ _21225_/X _21221_/B _21321_/Y vssd1 vssd1 vccd1 vccd1 _21330_/A sky130_fd_sc_hd__a21o_1
XFILLER_190_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1088 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21100__A _21121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19085__B1 _18617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21257_ _21254_/Y _21255_/X _21256_/Y vssd1 vssd1 vccd1 vccd1 _21257_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12722__A _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21967__B1 _21858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20208_ _20208_/A vssd1 vssd1 vccd1 vccd1 _20307_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21188_ _21290_/C _21210_/B _21211_/B vssd1 vssd1 vccd1 vccd1 _21188_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__12441__B _12441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15646__B1 _15664_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20139_ _19504_/X _19505_/X _17414_/B _17414_/A _20369_/B vssd1 vssd1 vccd1 vccd1
+ _20139_/Y sky130_fd_sc_hd__o2111ai_4
XANTENNA__19505__A _19505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12961_ _13107_/A _13107_/B _13107_/C _13109_/B _13109_/C vssd1 vssd1 vccd1 vccd1
+ _12962_/C sky130_fd_sc_hd__a32oi_4
XFILLER_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _23343_/Q _14689_/X _14694_/X _23311_/Q _14699_/X vssd1 vssd1 vccd1 vccd1
+ _14700_/X sky130_fd_sc_hd__a221o_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _11912_/A _11912_/B _11912_/C _11912_/D vssd1 vssd1 vccd1 vccd1 _11913_/C
+ sky130_fd_sc_hd__nand4_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _15630_/Y _15713_/B _14569_/X vssd1 vssd1 vccd1 vccd1 _15974_/D sky130_fd_sc_hd__a21o_2
XFILLER_166_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12880__B1 _12608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ _20805_/C _21124_/B vssd1 vssd1 vccd1 vccd1 _12899_/A sky130_fd_sc_hd__nand2_2
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _23427_/Q vssd1 vssd1 vccd1 vccd1 _14631_/X sky130_fd_sc_hd__buf_4
XFILLER_73_676 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _11846_/A vssd1 vssd1 vccd1 vccd1 _12053_/A sky130_fd_sc_hd__buf_2
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _17350_/A _17350_/B _17350_/C _17350_/D vssd1 vssd1 vccd1 vccd1 _17351_/C
+ sky130_fd_sc_hd__nand4_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14562_ _23417_/Q vssd1 vssd1 vccd1 vccd1 _15762_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11774_/A _11774_/B vssd1 vssd1 vccd1 vccd1 _12419_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _15761_/X _15762_/Y _16054_/X _16055_/X _15763_/Y vssd1 vssd1 vccd1 vccd1
+ _16402_/B sky130_fd_sc_hd__o221a_1
X_13513_ _13513_/A _13517_/C _13517_/A vssd1 vssd1 vccd1 vccd1 _13515_/B sky130_fd_sc_hd__nand3_1
XFILLER_158_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17281_ _17047_/A _17047_/B _17047_/C _17089_/C _17089_/D vssd1 vssd1 vccd1 vccd1
+ _17281_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14493_ _14493_/A _14493_/B vssd1 vssd1 vccd1 vccd1 _14496_/A sky130_fd_sc_hd__nand2_1
X_19020_ _16604_/A _11846_/A _19019_/Y vssd1 vssd1 vccd1 vccd1 _19020_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_186_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16232_ _16180_/Y _16181_/B _16181_/A vssd1 vssd1 vccd1 vccd1 _16234_/B sky130_fd_sc_hd__o21ai_1
X_13444_ _13444_/A vssd1 vssd1 vccd1 vccd1 _13599_/A sky130_fd_sc_hd__buf_2
XFILLER_70_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16400__A1_N _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12616__B _13121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17859__D1 _20055_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16163_ _12510_/A _16142_/B _15957_/C _16144_/B vssd1 vssd1 vccd1 vccd1 _16639_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_16_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13375_ _13796_/A vssd1 vssd1 vccd1 vccd1 _21766_/A sky130_fd_sc_hd__buf_2
XFILLER_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15114_ _23363_/Q _15114_/B vssd1 vssd1 vccd1 vccd1 _15115_/D sky130_fd_sc_hd__nand2_1
XFILLER_182_773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12326_ _16318_/C vssd1 vssd1 vccd1 vccd1 _12346_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16094_ _16094_/A _16094_/B vssd1 vssd1 vccd1 vccd1 _16331_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17845__D _17845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19922_ _19922_/A _19922_/B vssd1 vssd1 vccd1 vccd1 _23528_/D sky130_fd_sc_hd__xnor2_4
X_15045_ _15045_/A _15045_/B vssd1 vssd1 vccd1 vccd1 _15050_/C sky130_fd_sc_hd__nor2_1
X_12257_ _17133_/C vssd1 vssd1 vccd1 vccd1 _19503_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output71_A _14702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19853_ _19850_/Y _19851_/X _19863_/C vssd1 vssd1 vccd1 vccd1 _19853_/Y sky130_fd_sc_hd__o21ai_1
X_12188_ _12186_/Y _12187_/Y _11997_/X vssd1 vssd1 vccd1 vccd1 _12188_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_96_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11910__A2 _11907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18804_ _18804_/A _18804_/B vssd1 vssd1 vccd1 vccd1 _18808_/A sky130_fd_sc_hd__nand2_1
XFILLER_122_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19784_ _19775_/Y _19782_/X _19783_/X _19793_/A vssd1 vssd1 vccd1 vccd1 _19787_/B
+ sky130_fd_sc_hd__a22o_1
X_16996_ _17381_/A vssd1 vssd1 vccd1 vccd1 _16996_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_bq_clk_i_A bq_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22479__C _22637_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18735_ _19279_/A _19280_/A vssd1 vssd1 vccd1 vccd1 _18922_/A sky130_fd_sc_hd__or2_1
XFILLER_23_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15947_ _15782_/Y _15785_/Y _15651_/Y _15670_/X vssd1 vssd1 vccd1 vccd1 _15947_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12320__C1 _19534_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18666_ _18669_/C _18669_/D _18665_/C vssd1 vssd1 vccd1 vccd1 _18666_/X sky130_fd_sc_hd__a21o_2
XFILLER_92_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _20142_/A _16549_/C _15887_/C _15866_/B vssd1 vssd1 vccd1 vccd1 _15878_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_97_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17617_ _17462_/Y _17473_/C _17473_/D vssd1 vssd1 vccd1 vccd1 _17622_/A sky130_fd_sc_hd__a21boi_1
X_14829_ _14825_/A _14825_/B _14825_/C vssd1 vssd1 vccd1 vccd1 _14831_/B sky130_fd_sc_hd__a21oi_1
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18597_ _18756_/A _18597_/B _19364_/B vssd1 vssd1 vccd1 vccd1 _18598_/A sky130_fd_sc_hd__nand3_1
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12079__A _20217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14612__A1 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19536__D1 _17595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14612__B2 _15921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_186 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17548_ _17838_/A _17548_/B vssd1 vssd1 vccd1 vccd1 _17549_/C sky130_fd_sc_hd__nand2_1
XANTENNA__19551__A1 _19203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17479_ _17477_/Y _17478_/X _17290_/A vssd1 vssd1 vccd1 vccd1 _17482_/B sky130_fd_sc_hd__o21ai_1
XFILLER_177_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19218_ _19218_/A vssd1 vssd1 vccd1 vccd1 _19218_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14915__A2 _14050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20490_ _20490_/A _20490_/B vssd1 vssd1 vccd1 vccd1 _20490_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_910 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19303__A1 _19172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16117__A1 _17326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19149_ _19047_/A _19047_/C _19047_/B _18872_/Y _18844_/C vssd1 vssd1 vccd1 vccd1
+ _19149_/Y sky130_fd_sc_hd__a32oi_4
XANTENNA__17314__B1 _12323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22160_ _22388_/C _22160_/B vssd1 vssd1 vccd1 vccd1 _22160_/Y sky130_fd_sc_hd__nand2_2
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15837__B _16073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22016__A _22548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21111_ _21111_/A _21111_/B vssd1 vssd1 vccd1 vccd1 _21111_/Y sky130_fd_sc_hd__nand2_1
XFILLER_105_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22091_ _22667_/D _21987_/C _21987_/A _21989_/C _21989_/A vssd1 vssd1 vccd1 vccd1
+ _22093_/B sky130_fd_sc_hd__a32o_1
XFILLER_114_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21042_ _21174_/C _21174_/A vssd1 vssd1 vccd1 vccd1 _21043_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19970__D _20142_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17093__A2 _15618_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23492__D _23504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16668__B _16668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22993_ _21744_/B input8/X _23001_/S vssd1 vssd1 vccd1 vccd1 _22994_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21944_ _21892_/X _13765_/X _21893_/A _21893_/B _21798_/C vssd1 vssd1 vccd1 vccd1
+ _21944_/X sky130_fd_sc_hd__o221a_2
XFILLER_55_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21875_ _21875_/A _21875_/B vssd1 vssd1 vccd1 vccd1 _21875_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13406__A2 _22264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14603__A1 _12100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20137__C1 _17414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20826_ _20649_/Y _20646_/Y _20663_/Y _20664_/X vssd1 vssd1 vccd1 vccd1 _20828_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_51_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23545_ _23578_/CLK _23545_/D vssd1 vssd1 vccd1 vccd1 _23545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_882 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20152__A2 _20151_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20757_ _21414_/A _21415_/A _20751_/Y _20754_/X _20756_/Y vssd1 vssd1 vccd1 vccd1
+ _20761_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_156_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23582__CLK _23582_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20688_ _20688_/A _20688_/B _20688_/C vssd1 vssd1 vccd1 vccd1 _20715_/B sky130_fd_sc_hd__nand3_1
X_23476_ _23492_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 _23476_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22427_ _22430_/A _22427_/B _22427_/C vssd1 vssd1 vccd1 vccd1 _22457_/A sky130_fd_sc_hd__nand3b_1
XFILLER_136_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17305__B1 _12040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19845__A2 _19505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17856__A1 _17980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16659__A2 _16665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13160_ _13157_/Y _13158_/Y _13159_/X _13184_/A _12941_/A vssd1 vssd1 vccd1 vccd1
+ _13168_/B sky130_fd_sc_hd__o2111ai_4
X_22358_ _22356_/Y _22357_/Y _22357_/B vssd1 vssd1 vccd1 vccd1 _22436_/A sky130_fd_sc_hd__o21a_1
XFILLER_152_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12111_ _12107_/X _12110_/Y _12104_/X vssd1 vssd1 vccd1 vccd1 _12491_/B sky130_fd_sc_hd__a21oi_2
X_21309_ _21317_/A _21317_/B _21308_/C _21308_/D vssd1 vssd1 vccd1 vccd1 _21309_/X
+ sky130_fd_sc_hd__a22o_1
X_13091_ _13091_/A _20595_/C vssd1 vssd1 vccd1 vccd1 _13091_/Y sky130_fd_sc_hd__nand2_1
X_22289_ _22289_/A _22289_/B _22289_/C _22289_/D vssd1 vssd1 vccd1 vccd1 _22289_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_46_1011 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17608__A1 _17613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ _18481_/B _12040_/X _18941_/B _12166_/A _11996_/Y vssd1 vssd1 vccd1 vccd1
+ _12046_/A sky130_fd_sc_hd__a32o_1
XANTENNA__13342__A1 _22276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22601__A1 _22830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1052 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16850_ _15861_/X _16479_/A _16828_/A _17064_/A _16832_/Y vssd1 vssd1 vccd1 vccd1
+ _16850_/X sky130_fd_sc_hd__o221a_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15801_ _11738_/X _11740_/X _11741_/Y _15798_/A _15799_/A vssd1 vssd1 vccd1 vccd1
+ _15802_/A sky130_fd_sc_hd__o2111ai_4
XANTENNA__22299__C _22510_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16781_ _18435_/B _16781_/B vssd1 vssd1 vccd1 vccd1 _17218_/A sky130_fd_sc_hd__nor2_2
X_13993_ _23495_/Q vssd1 vssd1 vccd1 vccd1 _14252_/D sky130_fd_sc_hd__buf_2
XFILLER_46_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18520_ _18520_/A _18520_/B vssd1 vssd1 vccd1 vccd1 _18522_/A sky130_fd_sc_hd__nand2_1
X_15732_ _16805_/A vssd1 vssd1 vccd1 vccd1 _15860_/C sky130_fd_sc_hd__buf_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ _12709_/X _12936_/X _12654_/A _12627_/X _12604_/Y vssd1 vssd1 vccd1 vccd1
+ _12944_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _12429_/Y _12441_/B _12425_/X _12427_/X vssd1 vssd1 vccd1 vccd1 _18458_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14529__D input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15663_ _15712_/C vssd1 vssd1 vccd1 vccd1 _15920_/B sky130_fd_sc_hd__buf_2
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16595__A1 _11971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ _12875_/A _12875_/B _12875_/C vssd1 vssd1 vccd1 vccd1 _12876_/A sky130_fd_sc_hd__nand3_2
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _17134_/A _17326_/B _17326_/C vssd1 vssd1 vccd1 vccd1 _17493_/C sky130_fd_sc_hd__a21bo_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _21745_/B vssd1 vssd1 vccd1 vccd1 _14614_/X sky130_fd_sc_hd__clkbuf_4
X_18382_ _18410_/A _18411_/A _18382_/C vssd1 vssd1 vccd1 vccd1 _18383_/B sky130_fd_sc_hd__or3_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _12118_/A vssd1 vssd1 vccd1 vccd1 _11849_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15594_ _23517_/Q _15594_/B vssd1 vssd1 vccd1 vccd1 _23505_/D sky130_fd_sc_hd__xor2_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18336__A2 _17323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19533__B2 _18096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17333_ _17331_/A _17331_/B _17337_/A _17337_/B vssd1 vssd1 vccd1 vccd1 _17336_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12081__A1 _11916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14545_ _14545_/A vssd1 vssd1 vccd1 vccd1 _14545_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _11757_/A vssd1 vssd1 vccd1 vccd1 _18812_/A sky130_fd_sc_hd__buf_2
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17264_ _17610_/A _17285_/A _17260_/Y _17263_/Y vssd1 vssd1 vccd1 vccd1 _17275_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_105_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16898__A2 _16908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14476_ _15044_/C _14462_/Y _14461_/X _14472_/D _14472_/Y vssd1 vssd1 vccd1 vccd1
+ _14476_/X sky130_fd_sc_hd__a41o_1
XFILLER_174_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11688_ _18470_/C vssd1 vssd1 vccd1 vccd1 _18999_/C sky130_fd_sc_hd__buf_4
X_19003_ _18993_/Y _19000_/Y _19191_/A _19210_/A vssd1 vssd1 vccd1 vccd1 _19012_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_174_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16215_ _15902_/B _16202_/Y _16214_/Y vssd1 vssd1 vccd1 vccd1 _16215_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_146_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13427_ _13348_/X _13355_/A _13394_/A vssd1 vssd1 vccd1 vccd1 _21923_/A sky130_fd_sc_hd__a21o_1
XANTENNA__23093__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_954 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17195_ _17182_/X _17190_/Y _17200_/A vssd1 vssd1 vccd1 vccd1 _17195_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_128_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17847__A1 _16382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16146_ _16146_/A vssd1 vssd1 vccd1 vccd1 _16147_/A sky130_fd_sc_hd__buf_2
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _13358_/A vssd1 vssd1 vccd1 vccd1 _13358_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12309_ _12327_/A _16364_/A _16364_/B _16500_/D _12508_/A vssd1 vssd1 vccd1 vccd1
+ _12310_/A sky130_fd_sc_hd__a32o_1
X_16077_ _16326_/B _16061_/Y _16072_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 _16077_/X
+ sky130_fd_sc_hd__a31o_1
X_13289_ _13249_/A _13680_/B _13288_/Y vssd1 vssd1 vccd1 vccd1 _13303_/C sky130_fd_sc_hd__a21oi_1
XFILLER_170_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_776 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19905_ _19758_/Y _19757_/Y _19752_/Y _19745_/Y vssd1 vssd1 vccd1 vccd1 _19909_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15028_ _15077_/B _15035_/D vssd1 vssd1 vccd1 vccd1 _15028_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19836_ _19836_/A _19836_/B vssd1 vssd1 vccd1 vccd1 _19836_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16822__A2 _15749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19767_ _19932_/A _19771_/B _19771_/C _19932_/B vssd1 vssd1 vccd1 vccd1 _19928_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_96_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16979_ _16979_/A _16979_/B _16979_/C vssd1 vssd1 vccd1 vccd1 _16979_/Y sky130_fd_sc_hd__nand3_1
Xinput3 wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18718_ _18903_/A vssd1 vssd1 vccd1 vccd1 _18914_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19698_ _19698_/A _19903_/C _19698_/C _19800_/C vssd1 vssd1 vccd1 vccd1 _19717_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__19799__B _20062_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16035__B1 _16308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18649_ _18649_/A _19155_/C _19155_/D vssd1 vssd1 vccd1 vccd1 _18798_/A sky130_fd_sc_hd__nand3_2
XFILLER_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21660_ _21660_/A _21660_/B _21660_/C _21660_/D vssd1 vssd1 vccd1 vccd1 _21688_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_40_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18327__A2 _18376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14736__B _23596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20611_ _20611_/A _20611_/B vssd1 vssd1 vccd1 vccd1 _23540_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__12072__A1 _23256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21591_ _21548_/D _21432_/A _21432_/B _21635_/A _21635_/B vssd1 vssd1 vccd1 vccd1
+ _21598_/A sky130_fd_sc_hd__a311o_1
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20542_ _20542_/A _20542_/B _20542_/C vssd1 vssd1 vccd1 vccd1 _20553_/B sky130_fd_sc_hd__nand3_1
X_23330_ _23332_/CLK _23330_/D vssd1 vssd1 vccd1 vccd1 _23330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23261_ _23261_/A vssd1 vssd1 vccd1 vccd1 _23581_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__23084__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20473_ _20473_/A _20628_/C _20473_/C vssd1 vssd1 vccd1 vccd1 _20475_/A sky130_fd_sc_hd__nand3_1
XANTENNA__13021__B1 _20481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17766__C _17766_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23487__D _23499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12375__A2 _16480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22212_ _22044_/Y _22036_/X _22211_/Y _22197_/A vssd1 vssd1 vccd1 vccd1 _22214_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__22831__A1 _22830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23192_ _23192_/A vssd1 vssd1 vccd1 vccd1 _23416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1052 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22143_ _22028_/B _23331_/Q _23332_/Q vssd1 vssd1 vccd1 vccd1 _22144_/D sky130_fd_sc_hd__a21oi_1
XFILLER_156_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22074_ _22074_/A vssd1 vssd1 vccd1 vccd1 _22074_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21025_ _21025_/A _21029_/A _21029_/B vssd1 vssd1 vccd1 vccd1 _21031_/B sky130_fd_sc_hd__nand3_1
XFILLER_101_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18015__A1 _18001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22976_ _22976_/A vssd1 vssd1 vccd1 vccd1 _23320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19763__A1 _19380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21927_ _21927_/A vssd1 vssd1 vccd1 vccd1 _22548_/A sky130_fd_sc_hd__buf_2
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17774__B1 _17771_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17303__A _17303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12660_ _20966_/A _20966_/B _21039_/B vssd1 vssd1 vccd1 vccd1 _12661_/B sky130_fd_sc_hd__and3_1
XFILLER_150_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21858_ _13867_/Y _21858_/B _21981_/A _21858_/D vssd1 vssd1 vccd1 vccd1 _21859_/B
+ sky130_fd_sc_hd__nand4b_1
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14052__A2 _14050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11611_ _11611_/A _11611_/B vssd1 vssd1 vccd1 vccd1 _12260_/C sky130_fd_sc_hd__nand2_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _20809_/A _20809_/B vssd1 vssd1 vccd1 vccd1 _20810_/B sky130_fd_sc_hd__nand2_1
X_12591_ _23287_/Q vssd1 vssd1 vccd1 vccd1 _12606_/C sky130_fd_sc_hd__inv_2
XFILLER_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21789_ _21875_/A _21789_/B _21875_/B vssd1 vssd1 vccd1 vccd1 _21805_/B sky130_fd_sc_hd__nand3_1
XFILLER_184_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14330_ _14330_/A vssd1 vssd1 vccd1 vccd1 _14381_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_23528_ _23538_/CLK _23528_/D vssd1 vssd1 vccd1 vccd1 _23528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23040__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15758__A _16612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14261_ _14261_/A vssd1 vssd1 vccd1 vccd1 _14751_/B sky130_fd_sc_hd__buf_2
XFILLER_7_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23459_ _23492_/CLK _23471_/Q vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_183_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16000_ _16000_/A _16000_/B _16000_/C vssd1 vssd1 vccd1 vccd1 _16000_/Y sky130_fd_sc_hd__nand3_1
XFILLER_13_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13212_ _20611_/A _13212_/B vssd1 vssd1 vccd1 vccd1 _13213_/A sky130_fd_sc_hd__or2_1
XFILLER_183_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14192_ _23358_/Q _23357_/Q vssd1 vssd1 vccd1 vccd1 _14193_/B sky130_fd_sc_hd__nor2_1
XFILLER_152_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_890 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13143_ _13143_/A _13143_/B _13143_/C vssd1 vssd1 vccd1 vccd1 _13196_/C sky130_fd_sc_hd__nand3_1
XANTENNA__12182__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16501__B2 _16526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17951_ _17951_/A _18148_/A _17951_/C _17951_/D vssd1 vssd1 vccd1 vccd1 _17952_/C
+ sky130_fd_sc_hd__nand4_2
X_13074_ _13078_/A _13078_/B _13079_/B vssd1 vssd1 vccd1 vccd1 _13089_/C sky130_fd_sc_hd__nand3_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16902_ _12004_/X _12006_/X _16677_/B _16213_/A vssd1 vssd1 vccd1 vccd1 _16902_/Y
+ sky130_fd_sc_hd__o211ai_2
X_12025_ _12131_/A vssd1 vssd1 vccd1 vccd1 _12025_/X sky130_fd_sc_hd__clkbuf_2
X_17882_ _17868_/Y _17873_/Y _17881_/Y vssd1 vssd1 vccd1 vccd1 _17902_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11877__A1 _16464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11877__B2 _19040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19621_ _18673_/X _20368_/B _19358_/Y _18373_/A _12353_/X vssd1 vssd1 vccd1 vccd1
+ _19621_/X sky130_fd_sc_hd__o32a_2
XFILLER_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16833_ _16828_/A _17064_/A _16832_/Y vssd1 vssd1 vccd1 vccd1 _16841_/A sky130_fd_sc_hd__o21ai_1
XFILLER_66_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19552_ _19560_/A _19552_/B _19552_/C vssd1 vssd1 vccd1 vccd1 _19552_/Y sky130_fd_sc_hd__nand3b_1
X_16764_ _16759_/B _16759_/C _16486_/Y _16492_/Y vssd1 vssd1 vccd1 vccd1 _16764_/Y
+ sky130_fd_sc_hd__a22oi_1
X_13976_ _14863_/C _14863_/D _13946_/A vssd1 vssd1 vccd1 vccd1 _13977_/A sky130_fd_sc_hd__o21ai_1
XFILLER_46_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18503_ _18503_/A _18503_/B _18503_/C _18503_/D vssd1 vssd1 vccd1 vccd1 _18503_/Y
+ sky130_fd_sc_hd__nand4_4
X_15715_ _15715_/A _15735_/B vssd1 vssd1 vccd1 vccd1 _15716_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12927_ _21050_/D vssd1 vssd1 vccd1 vccd1 _21182_/D sky130_fd_sc_hd__buf_2
X_19483_ _17627_/A _19190_/A _19670_/C _19480_/X _19482_/Y vssd1 vssd1 vccd1 vccd1
+ _19483_/Y sky130_fd_sc_hd__o221ai_4
X_16695_ _16939_/A _16939_/B _16706_/A _16706_/B vssd1 vssd1 vccd1 vccd1 _16699_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_624 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13741__A _22474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18434_ _18434_/A _18434_/B vssd1 vssd1 vccd1 vccd1 _19279_/A sky130_fd_sc_hd__nor2_4
XFILLER_94_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15646_ _15644_/X _15921_/B _15664_/C vssd1 vssd1 vccd1 vccd1 _15647_/B sky130_fd_sc_hd__a21oi_2
XFILLER_22_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12858_ _12858_/A _12858_/B vssd1 vssd1 vccd1 vccd1 _12859_/C sky130_fd_sc_hd__nand2_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19506__A1 _19504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18365_ _18363_/Y _18364_/Y _18319_/D vssd1 vssd1 vccd1 vccd1 _18365_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11809_ _11809_/A _16796_/A vssd1 vssd1 vccd1 vccd1 _11809_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12054__A1 _12311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15577_ _15577_/A _23508_/Q _23509_/Q _23510_/Q vssd1 vssd1 vccd1 vccd1 _15585_/D
+ sky130_fd_sc_hd__or4_2
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12824_/B vssd1 vssd1 vccd1 vccd1 _13119_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17316_ _16464_/X _17304_/A _17140_/B _17305_/Y _17307_/Y vssd1 vssd1 vccd1 vccd1
+ _17316_/Y sky130_fd_sc_hd__o221ai_4
X_14528_ input41/X _14518_/X _14527_/X vssd1 vssd1 vccd1 vccd1 _14528_/X sky130_fd_sc_hd__a21o_1
X_18296_ _18296_/A vssd1 vssd1 vccd1 vccd1 _18296_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20521__C1 _12980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17247_ _17050_/X _16819_/X _15884_/A vssd1 vssd1 vccd1 vccd1 _17450_/B sky130_fd_sc_hd__a21oi_1
XFILLER_119_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14459_ _14459_/A _14469_/C _15233_/C _14459_/D vssd1 vssd1 vccd1 vccd1 _14472_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19809__A2 _18455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13554__A1 _22474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17178_ _17179_/B _17179_/C _17179_/A vssd1 vssd1 vccd1 vccd1 _17178_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17883__A _19957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16129_ _11935_/X _16377_/A _15975_/B _16128_/X _16610_/A vssd1 vssd1 vccd1 vccd1
+ _16129_/X sky130_fd_sc_hd__o221a_1
XFILLER_116_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_916 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16499__A _16499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15059__A1 _15538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19819_ _19819_/A _19819_/B vssd1 vssd1 vccd1 vccd1 _19820_/B sky130_fd_sc_hd__nand2_1
XFILLER_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17107__B _17235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22830_ _22830_/A _22830_/B _22830_/C _22830_/D vssd1 vssd1 vccd1 vccd1 _22830_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21852__B _23482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23125__A _23182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22761_ _21997_/X _22830_/C _22830_/D _22707_/A vssd1 vssd1 vccd1 vccd1 _22762_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14747__A _15338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21712_ _23576_/Q vssd1 vssd1 vccd1 vccd1 _21712_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22692_ _22818_/C _22821_/A vssd1 vssd1 vccd1 vccd1 _22694_/C sky130_fd_sc_hd__nand2_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21643_ _21643_/A _21643_/B vssd1 vssd1 vccd1 vccd1 _21645_/C sky130_fd_sc_hd__xnor2_1
XFILLER_178_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12267__A _18947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15782__A2 _15781_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21855__A2 _21858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21574_ _21473_/A _21524_/A _21524_/C vssd1 vssd1 vccd1 vccd1 _21574_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23313_ _23345_/CLK _23313_/D vssd1 vssd1 vccd1 vccd1 _23313_/Q sky130_fd_sc_hd__dfxtp_1
X_20525_ _12674_/X _12714_/X _12957_/Y _13018_/Y _13021_/Y vssd1 vssd1 vccd1 vccd1
+ _20525_/X sky130_fd_sc_hd__o32a_1
XANTENNA__12417__D _15699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_654 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20456_ _20448_/A _20448_/B _20454_/Y _20455_/Y vssd1 vssd1 vccd1 vccd1 _20457_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_181_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23244_ _23440_/Q input25/X _23250_/S vssd1 vssd1 vccd1 vccd1 _23245_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20815__B1 _21054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20387_ _20411_/B vssd1 vssd1 vccd1 vccd1 _20415_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_23175_ _23175_/A vssd1 vssd1 vccd1 vccd1 _23409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17141__D1 _19653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22126_ _22126_/A vssd1 vssd1 vccd1 vccd1 _22126_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22057_ _22057_/A vssd1 vssd1 vccd1 vccd1 _22057_/X sky130_fd_sc_hd__buf_2
XFILLER_43_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21008_ _21008_/A _21008_/B _21008_/C vssd1 vssd1 vccd1 vccd1 _21008_/X sky130_fd_sc_hd__and3_1
XFILLER_102_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13830_ _13822_/Y _13824_/Y _13829_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13264__C _13264_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ _13540_/A _13540_/B _13540_/C _13543_/Y _13535_/A vssd1 vssd1 vccd1 vccd1
+ _21856_/C sky130_fd_sc_hd__a32o_2
XANTENNA__12284__A1 _12282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22959_ _22959_/A vssd1 vssd1 vccd1 vccd1 _23313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15500_ _15501_/A _15501_/B _15501_/C vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__a21oi_1
XFILLER_188_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12712_ _12712_/A vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__buf_4
X_16480_ _16480_/A vssd1 vssd1 vccd1 vccd1 _16480_/X sky130_fd_sc_hd__buf_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _13692_/A _13692_/B _13692_/C vssd1 vssd1 vccd1 vccd1 _13760_/A sky130_fd_sc_hd__nand3_1
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15431_ _15431_/A _15431_/B vssd1 vssd1 vccd1 vccd1 _15433_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__17968__A _18080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ _13011_/A _20639_/A _13011_/C _13011_/D vssd1 vssd1 vccd1 vccd1 _12688_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18150_ _18144_/B _18149_/B _18144_/C vssd1 vssd1 vccd1 vccd1 _18150_/X sky130_fd_sc_hd__a21bo_1
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15362_ _15096_/A _15096_/B _15358_/A _15416_/A _15415_/A vssd1 vssd1 vccd1 vccd1
+ _15363_/C sky130_fd_sc_hd__a32o_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12574_ _23288_/Q vssd1 vssd1 vccd1 vccd1 _20493_/B sky130_fd_sc_hd__buf_2
XFILLER_184_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17101_ _16832_/Y _16841_/B _16828_/Y vssd1 vssd1 vccd1 vccd1 _17106_/A sky130_fd_sc_hd__a21oi_1
XFILLER_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16591__B _16591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14313_ _14407_/B vssd1 vssd1 vccd1 vccd1 _14344_/B sky130_fd_sc_hd__clkbuf_2
X_18081_ _19705_/A vssd1 vssd1 vccd1 vccd1 _20215_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15488__A _15488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15293_ _15293_/A _15293_/B vssd1 vssd1 vccd1 vccd1 _15332_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17032_ _17032_/A _17032_/B vssd1 vssd1 vccd1 vccd1 _17891_/A sky130_fd_sc_hd__nand2_2
XFILLER_144_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14244_ _13951_/A _13951_/B _14097_/A vssd1 vssd1 vccd1 vccd1 _14245_/B sky130_fd_sc_hd__a21o_1
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14175_ _14121_/B _14756_/A _14174_/Y vssd1 vssd1 vccd1 vccd1 _14177_/A sky130_fd_sc_hd__o21ai_1
XFILLER_178_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13126_ _13117_/X _13126_/B _13126_/C vssd1 vssd1 vccd1 vccd1 _13172_/A sky130_fd_sc_hd__nand3b_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _18983_/A _18983_/B _18983_/C vssd1 vssd1 vccd1 vccd1 _19043_/A sky130_fd_sc_hd__nand3_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _17934_/A _17934_/B vssd1 vssd1 vccd1 vccd1 _18058_/D sky130_fd_sc_hd__nor2_2
XANTENNA__23220__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13115_/A _13115_/B _20669_/C vssd1 vssd1 vccd1 vccd1 _13058_/A sky130_fd_sc_hd__nand3_1
XFILLER_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16112__A _18093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater106 _23325_/CLK vssd1 vssd1 vccd1 vccd1 _23332_/CLK sky130_fd_sc_hd__clkbuf_1
X_12008_ _11822_/A _18500_/A _12002_/Y _12007_/Y _12166_/A vssd1 vssd1 vccd1 vccd1
+ _12008_/X sky130_fd_sc_hd__o221a_1
Xrepeater117 _23416_/CLK vssd1 vssd1 vccd1 vccd1 _23428_/CLK sky130_fd_sc_hd__clkbuf_1
X_17865_ _17644_/A _18003_/A _17858_/Y vssd1 vssd1 vccd1 vccd1 _18013_/A sky130_fd_sc_hd__o21ai_2
Xrepeater128 _23398_/CLK vssd1 vssd1 vccd1 vccd1 _23336_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater139 _23434_/CLK vssd1 vssd1 vccd1 vccd1 _23409_/CLK sky130_fd_sc_hd__clkbuf_1
X_19604_ _19406_/A _19420_/A _19603_/Y vssd1 vssd1 vccd1 vccd1 _19605_/C sky130_fd_sc_hd__a21oi_1
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16816_ _12510_/A _16816_/B _16816_/C vssd1 vssd1 vccd1 vccd1 _16816_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_94_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17796_ _17790_/Y _17919_/B _17795_/X vssd1 vssd1 vccd1 vccd1 _17796_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23590__D _23590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19535_ _18435_/A _11841_/Y _11849_/A _19700_/C _19700_/D vssd1 vssd1 vccd1 vccd1
+ _19547_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16747_ _18161_/B vssd1 vssd1 vccd1 vccd1 _18279_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13959_ _14795_/C vssd1 vssd1 vccd1 vccd1 _15254_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__13472__B1 _13470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19466_ _19430_/Y _19432_/Y _19464_/Y _19465_/X vssd1 vssd1 vccd1 vccd1 _19467_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_34_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16678_ _16904_/A vssd1 vssd1 vccd1 vccd1 _16911_/B sky130_fd_sc_hd__buf_2
XFILLER_179_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18417_ _18417_/A _18417_/B _18417_/C _18417_/D vssd1 vssd1 vccd1 vccd1 _18420_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_50_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15629_ _15685_/A vssd1 vssd1 vccd1 vccd1 _16187_/B sky130_fd_sc_hd__clkbuf_2
X_19397_ _19601_/A _19601_/B _19468_/A _19600_/A vssd1 vssd1 vccd1 vccd1 _19402_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12087__A _17610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16782__A _17217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18348_ _18348_/A _18348_/B vssd1 vssd1 vccd1 vccd1 _18349_/C sky130_fd_sc_hd__nor2_1
XFILLER_188_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18279_ _18279_/A _18279_/B _19900_/A _18279_/D vssd1 vssd1 vccd1 vccd1 _18279_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_163_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20310_ _20310_/A _20310_/B _20310_/C vssd1 vssd1 vccd1 vccd1 _20312_/B sky130_fd_sc_hd__nand3_1
XFILLER_162_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 x[7] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_4
X_21290_ _21380_/A _21290_/B _21290_/C vssd1 vssd1 vccd1 vccd1 _21317_/B sky130_fd_sc_hd__nand3b_2
XFILLER_128_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20241_ _20290_/B _20242_/B _20243_/B vssd1 vssd1 vccd1 vccd1 _20244_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__17269__A2 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19663__B1 _17643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22262__A2 _13431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20172_ _20172_/A _20172_/B vssd1 vssd1 vccd1 vccd1 _20176_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19317__B _19321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18859__D _18859_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23211__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16229__B1 _17420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18769__A2 _17846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13160__C1 _13184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17977__B1 _20210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12700__D _21054_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17441__A2 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19179__C1 _19178_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15452__A1 _15371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22813_ _22813_/A _22813_/B vssd1 vssd1 vccd1 vccd1 _22828_/A sky130_fd_sc_hd__nor2_2
XANTENNA__12266__A1 _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19194__A2 _19196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22744_ _22623_/B _22623_/C _22623_/A vssd1 vssd1 vccd1 vccd1 _22745_/A sky130_fd_sc_hd__a21oi_1
XFILLER_197_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11613__B _15991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22675_ _22675_/A _22675_/B vssd1 vssd1 vccd1 vccd1 _22675_/Y sky130_fd_sc_hd__nand2_1
XFILLER_197_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21626_ _23570_/Q _21579_/C _21579_/A _21540_/B vssd1 vssd1 vccd1 vccd1 _21626_/Y
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__22486__C1 _22392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21557_ _21590_/A _21590_/B vssd1 vssd1 vccd1 vccd1 _21557_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20500__A2 _21431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20508_ _20502_/X _20504_/X _20645_/C _20496_/X vssd1 vssd1 vccd1 vccd1 _20509_/B
+ sky130_fd_sc_hd__o211ai_4
X_12290_ _12090_/A _12279_/X _12244_/X _12271_/A _12289_/A vssd1 vssd1 vccd1 vccd1
+ _12291_/B sky130_fd_sc_hd__o311a_1
XFILLER_107_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21488_ _21400_/A _21400_/B _21476_/A vssd1 vssd1 vccd1 vccd1 _21488_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16180__A2 _15985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23227_ _23227_/A vssd1 vssd1 vccd1 vccd1 _23432_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18457__A1 _19803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20439_ _20449_/A _20449_/B _20438_/A vssd1 vssd1 vccd1 vccd1 _20442_/B sky130_fd_sc_hd__a21oi_1
XFILLER_106_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20661__B _20894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23158_ _23169_/A vssd1 vssd1 vccd1 vccd1 _23167_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_134_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22109_ _22348_/B _22348_/C _22249_/B _21980_/A vssd1 vssd1 vccd1 vccd1 _22109_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15980_ _15889_/X _15971_/X _15976_/Y _15979_/Y vssd1 vssd1 vccd1 vccd1 _15995_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23202__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23089_ _23371_/Q input20/X _23095_/S vssd1 vssd1 vccd1 vccd1 _23090_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A wb_dat_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14931_ _14943_/B _14966_/B _14943_/A vssd1 vssd1 vccd1 vccd1 _14931_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_121_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17650_ _17657_/B _17657_/C vssd1 vssd1 vccd1 vccd1 _17656_/C sky130_fd_sc_hd__nand2_1
XANTENNA__17432__A2 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14862_ _13937_/X _14860_/Y _15112_/B vssd1 vssd1 vccd1 vccd1 _15094_/A sky130_fd_sc_hd__o21ai_1
XFILLER_36_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1024 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_771 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16640__B1 _16064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16601_ _17108_/B _16601_/B _16601_/C _18859_/D vssd1 vssd1 vccd1 vccd1 _16601_/Y
+ sky130_fd_sc_hd__nand4_2
X_13813_ _13813_/A vssd1 vssd1 vccd1 vccd1 _13813_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17581_ _17581_/A vssd1 vssd1 vccd1 vccd1 _18778_/A sky130_fd_sc_hd__buf_2
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14793_ _14798_/A _14911_/B _14793_/C vssd1 vssd1 vccd1 vccd1 _14793_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__22174__D1 _22487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19320_ _19320_/A vssd1 vssd1 vccd1 vccd1 _19525_/A sky130_fd_sc_hd__clkbuf_2
X_16532_ _16532_/A _16532_/B _16532_/C vssd1 vssd1 vccd1 vccd1 _16564_/A sky130_fd_sc_hd__nand3_1
XFILLER_17_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13744_ _13744_/A _13744_/B _22192_/D _21832_/A vssd1 vssd1 vccd1 vccd1 _13744_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19251_ _18968_/A _19246_/Y _19236_/Y _19245_/X _18969_/D vssd1 vssd1 vccd1 vccd1
+ _19434_/C sky130_fd_sc_hd__o2111ai_4
X_16463_ _16438_/Y _16364_/X _16462_/X vssd1 vssd1 vccd1 vccd1 _16463_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_31_413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13675_ _13671_/A _13671_/B _13672_/X _13674_/X vssd1 vssd1 vccd1 vccd1 _13676_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_18202_ _18122_/Y _18192_/Y _18195_/Y vssd1 vssd1 vccd1 vccd1 _18302_/A sky130_fd_sc_hd__o21ai_2
X_15414_ _15377_/A _15377_/B _15382_/B vssd1 vssd1 vccd1 vccd1 _15463_/B sky130_fd_sc_hd__o21ai_1
X_19182_ _19332_/B _19182_/B vssd1 vssd1 vccd1 vccd1 _19183_/C sky130_fd_sc_hd__nor2_2
Xclkbuf_0_bq_clk_i bq_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_bq_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_12626_ _20620_/C vssd1 vssd1 vccd1 vccd1 _12932_/A sky130_fd_sc_hd__clkinv_2
X_16394_ _16394_/A vssd1 vssd1 vccd1 vccd1 _16517_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18133_ _18133_/A _18133_/B vssd1 vssd1 vccd1 vccd1 _18134_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19003__A1_N _18993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15345_ _15345_/A vssd1 vssd1 vccd1 vccd1 _23277_/D sky130_fd_sc_hd__clkbuf_1
X_12557_ _12557_/A _18571_/A _18571_/B vssd1 vssd1 vccd1 vccd1 _19089_/B sky130_fd_sc_hd__nand3_4
XFILLER_89_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18064_ _18062_/Y _17952_/C _18144_/B _18063_/Y vssd1 vssd1 vccd1 vccd1 _18066_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_144_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15276_ _15276_/A _15294_/B vssd1 vssd1 vccd1 vccd1 _15277_/C sky130_fd_sc_hd__nand2_1
XFILLER_184_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12488_ _12490_/A _12490_/B _12480_/A _12480_/B vssd1 vssd1 vccd1 vccd1 _12494_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_89_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17015_ _17014_/B _17014_/C _17014_/A vssd1 vssd1 vccd1 vccd1 _17015_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14182__A1 _14181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14227_ _14227_/A _14227_/B vssd1 vssd1 vccd1 vccd1 _14228_/B sky130_fd_sc_hd__nor2_1
XANTENNA__19645__B1 _19648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23585__D _23585_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16459__B1 _16356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14158_ _14150_/D _15019_/A _14407_/A _13985_/X vssd1 vssd1 vccd1 vccd1 _14818_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _13109_/A _13109_/B _13109_/C vssd1 vssd1 vccd1 vccd1 _13136_/C sky130_fd_sc_hd__nand3_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ _18966_/A _18966_/B vssd1 vssd1 vccd1 vccd1 _18969_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14089_ _23495_/Q vssd1 vssd1 vccd1 vccd1 _14089_/Y sky130_fd_sc_hd__clkinv_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _17913_/Y _17917_/B _17917_/C vssd1 vssd1 vccd1 vccd1 _17919_/D sky130_fd_sc_hd__nand3b_1
XFILLER_113_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18897_ _18904_/A _18904_/B _18897_/C _18897_/D vssd1 vssd1 vccd1 vccd1 _18899_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_39_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15681__A _15974_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17848_ _17974_/C _20133_/D _17855_/A _17853_/A vssd1 vssd1 vccd1 vccd1 _17848_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17779_ _17779_/A _17779_/B _17779_/C vssd1 vssd1 vccd1 vccd1 _17779_/Y sky130_fd_sc_hd__nand3_2
XFILLER_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18992__A _19186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__A _16677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19518_ _19524_/B _19524_/C _19524_/A vssd1 vssd1 vccd1 vccd1 _19519_/D sky130_fd_sc_hd__nand3b_1
XANTENNA__13996__A1 _15353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13996__B2 _14867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20790_ _20790_/A _20790_/B vssd1 vssd1 vccd1 vccd1 _20794_/A sky130_fd_sc_hd__nand2_1
XANTENNA__22180__A1 _14614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19449_ _19793_/A _19295_/X _19448_/Y vssd1 vssd1 vccd1 vccd1 _19449_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22460_ _22541_/A _22541_/B vssd1 vssd1 vccd1 vccd1 _22499_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_619 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22019__A _23331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21411_ _21411_/A _21411_/B vssd1 vssd1 vccd1 vccd1 _21411_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22391_ _22391_/A vssd1 vssd1 vccd1 vccd1 _22392_/A sky130_fd_sc_hd__buf_2
XFILLER_191_900 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21342_ _21354_/A _21342_/B _21342_/C vssd1 vssd1 vccd1 vccd1 _21342_/Y sky130_fd_sc_hd__nand3_1
XFILLER_136_838 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21273_ _21273_/A vssd1 vssd1 vccd1 vccd1 _21397_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20481__B _20481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23012_ _23337_/Q input17/X _23012_/S vssd1 vssd1 vccd1 vccd1 _23013_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20224_ _20221_/X _20223_/Y _20083_/A vssd1 vssd1 vccd1 vccd1 _20224_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20155_ _20083_/Y _20131_/X _20150_/Y _20154_/X vssd1 vssd1 vccd1 vccd1 _20167_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_131_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_991 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20086_ _20086_/A _20159_/C vssd1 vssd1 vccd1 vccd1 _20095_/C sky130_fd_sc_hd__nor2_2
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_719 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15976__A2 _15972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15830__D1 _18481_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11723_/A _11918_/A _11739_/B vssd1 vssd1 vccd1 vccd1 _11792_/A sky130_fd_sc_hd__o21ai_4
XFILLER_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18375__B1 _18376_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20988_ _20994_/B _20994_/C vssd1 vssd1 vccd1 vccd1 _20990_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22727_ _22678_/X _22675_/Y _22676_/Y vssd1 vssd1 vccd1 vccd1 _22750_/B sky130_fd_sc_hd__a21bo_1
XFILLER_159_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16386__C1 _17243_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_727 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1096 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13460_ _13460_/A _13474_/A _13474_/B _13460_/D vssd1 vssd1 vccd1 vccd1 _13461_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_159_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22658_ _22581_/X _22657_/Y _22584_/C vssd1 vssd1 vccd1 vccd1 _22658_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_90_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12411_ _18810_/A vssd1 vssd1 vccd1 vccd1 _18997_/A sky130_fd_sc_hd__buf_2
XFILLER_90_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21609_ _21568_/A _21589_/Y _21608_/Y vssd1 vssd1 vccd1 vccd1 _21630_/A sky130_fd_sc_hd__o21ai_2
XFILLER_159_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13391_ _13323_/X _13338_/X _13377_/C _22022_/A _13379_/X vssd1 vssd1 vccd1 vccd1
+ _13392_/B sky130_fd_sc_hd__a311o_1
XFILLER_51_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22589_ _22589_/A _22589_/B _22589_/C vssd1 vssd1 vccd1 vccd1 _22598_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12455__A _19648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15130_ _15129_/A _15130_/B _15130_/C vssd1 vssd1 vccd1 vccd1 _15132_/B sky130_fd_sc_hd__nand3b_1
X_12342_ _19512_/D vssd1 vssd1 vccd1 vccd1 _17546_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_181_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ _15060_/X _14941_/Y _14945_/Y _14953_/C _14951_/X vssd1 vssd1 vccd1 vccd1
+ _15067_/A sky130_fd_sc_hd__a32o_2
X_12273_ _12273_/A _12273_/B _12273_/C _12273_/D vssd1 vssd1 vccd1 vccd1 _12295_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_49_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15900__A2 _11807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ _14012_/A vssd1 vssd1 vccd1 vccd1 _14015_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20788__A2 _20786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11922__B1 _23591_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18820_ _19505_/A _19504_/A _19000_/B _19157_/A vssd1 vssd1 vccd1 vccd1 _18820_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15113__B1 _23364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23187__A0 _16510_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16861__B1 _11971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18751_ _18751_/A _18751_/B _18751_/C vssd1 vssd1 vccd1 vccd1 _18751_/X sky130_fd_sc_hd__and3_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15963_ _15862_/A _15862_/B _17061_/A _17060_/A vssd1 vssd1 vccd1 vccd1 _16153_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17702_ _17385_/Y _17701_/X _17537_/A vssd1 vssd1 vccd1 vccd1 _17703_/C sky130_fd_sc_hd__o21a_1
XANTENNA__18602__A1 _12167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14914_ _13933_/A _15084_/A _14911_/Y _14910_/X vssd1 vssd1 vccd1 vccd1 _14918_/B
+ sky130_fd_sc_hd__o211ai_2
X_18682_ _18784_/A vssd1 vssd1 vccd1 vccd1 _18880_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15894_ _15894_/A vssd1 vssd1 vccd1 vccd1 _15895_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22111__B _22112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16613__B1 _16612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17633_ _17723_/C _17960_/B _18016_/D vssd1 vssd1 vccd1 vccd1 _17634_/B sky130_fd_sc_hd__and3_1
XFILLER_1_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14845_ _15065_/A _14853_/B vssd1 vssd1 vccd1 vccd1 _14845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19123__D _19548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17564_ _17562_/Y _17563_/Y _17473_/D vssd1 vssd1 vccd1 vccd1 _17616_/A sky130_fd_sc_hd__o21ai_4
X_14776_ _14245_/A _14773_/Y _14775_/Y vssd1 vssd1 vccd1 vccd1 _14778_/A sky130_fd_sc_hd__o21ai_1
X_11988_ _15699_/A _12183_/A _11982_/Y _11987_/Y vssd1 vssd1 vccd1 vccd1 _12166_/A
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_44_560 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19303_ _19172_/A _19172_/B _19172_/C _19183_/C vssd1 vssd1 vccd1 vccd1 _19303_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_56_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16515_ _16356_/X _16458_/X _16514_/X _16384_/X _16370_/X vssd1 vssd1 vccd1 vccd1
+ _16522_/B sky130_fd_sc_hd__o32a_1
X_13727_ _13727_/A _13727_/B _13723_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_72_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17495_ _17497_/A _17497_/B _17497_/C _17497_/D vssd1 vssd1 vccd1 vccd1 _17498_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19234_ _19060_/B _19057_/D _19058_/A vssd1 vssd1 vccd1 vccd1 _19257_/A sky130_fd_sc_hd__a21boi_2
XFILLER_56_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16446_ _16446_/A _16446_/B vssd1 vssd1 vccd1 vccd1 _16507_/A sky130_fd_sc_hd__nand2_4
X_13658_ _13660_/A _21882_/B _13660_/C vssd1 vssd1 vccd1 vccd1 _13658_/Y sky130_fd_sc_hd__nand3_2
XFILLER_20_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12609_ _12606_/Y _20495_/C _12608_/X vssd1 vssd1 vccd1 vccd1 _20528_/A sky130_fd_sc_hd__a21o_2
XFILLER_157_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16377_ _16377_/A vssd1 vssd1 vccd1 vccd1 _16377_/X sky130_fd_sc_hd__buf_2
X_19165_ _19502_/A _19308_/B _19165_/C _20369_/C vssd1 vssd1 vccd1 vccd1 _19165_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13589_ _13554_/X _13555_/Y _13507_/Y _13494_/Y vssd1 vssd1 vccd1 vccd1 _13590_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_76_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18116_ _18033_/A _18033_/C _18033_/B vssd1 vssd1 vccd1 vccd1 _18298_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__19330__A2 _19803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15328_ _15328_/A _15380_/B _15328_/C vssd1 vssd1 vccd1 vccd1 _15328_/Y sky130_fd_sc_hd__nand3_2
XFILLER_173_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19096_ _19106_/A _19106_/B _19095_/Y _19108_/A vssd1 vssd1 vccd1 vccd1 _19101_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18047_ _17922_/X _17924_/X _17930_/Y _17957_/Y vssd1 vssd1 vccd1 vccd1 _18053_/A
+ sky130_fd_sc_hd__o22ai_2
X_15259_ _15259_/A _15259_/B _15259_/C vssd1 vssd1 vccd1 vccd1 _15259_/Y sky130_fd_sc_hd__nand3_1
XFILLER_132_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19998_ _19992_/X _19835_/Y _19987_/Y _19991_/Y vssd1 vssd1 vccd1 vccd1 _19998_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13627__C _13816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1159 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18949_ _12089_/A _18096_/A _18945_/Y _19261_/A vssd1 vssd1 vccd1 vccd1 _18950_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__22302__A _22476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22925__A0 _20894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21960_ _21964_/A _21964_/B _21964_/C vssd1 vssd1 vccd1 vccd1 _21961_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__15842__C _16612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20911_ _20494_/D _20498_/A _13018_/Y vssd1 vssd1 vccd1 vccd1 _20911_/X sky130_fd_sc_hd__a21o_1
XFILLER_54_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21891_ _21891_/A _22558_/A vssd1 vssd1 vccd1 vccd1 _21891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15812__D1 _16365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19611__A _20320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20842_ _20842_/A _20842_/B vssd1 vssd1 vccd1 vccd1 _20843_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19554__C1 _18673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23561_ _23566_/CLK _23561_/D vssd1 vssd1 vccd1 vccd1 _23561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20773_ _20773_/A _20773_/B _20773_/C _20773_/D vssd1 vssd1 vccd1 vccd1 _21000_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_161_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22512_ _22505_/X _22507_/Y _22509_/X _22511_/Y vssd1 vssd1 vccd1 vccd1 _22513_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23492_ _23492_/CLK _23504_/Q vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16383__A2 _17285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22443_ _22443_/A _22443_/B vssd1 vssd1 vccd1 vccd1 _22443_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22374_ _22122_/Y _22362_/A _22300_/B _22297_/Y vssd1 vssd1 vccd1 vccd1 _22504_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_135_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21325_ _21311_/Y _21320_/Y _21322_/Y _21324_/X vssd1 vssd1 vccd1 vccd1 _21331_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_136_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15343__B1 _15442_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14490__A _15082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21256_ _23565_/Q vssd1 vssd1 vccd1 vccd1 _21256_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19085__B2 _18928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20207_ _20207_/A _20207_/B _20207_/C _20207_/D vssd1 vssd1 vccd1 vccd1 _20208_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11619__A _12167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21187_ _21187_/A _21187_/B vssd1 vssd1 vccd1 vccd1 _21211_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20138_ _20138_/A _20138_/B _20320_/B _20320_/C vssd1 vssd1 vccd1 vccd1 _20138_/X
+ sky130_fd_sc_hd__and4_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22916__A0 _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20069_ _20071_/A _20160_/A _20071_/C vssd1 vssd1 vccd1 vccd1 _20069_/X sky130_fd_sc_hd__and3_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _12949_/Y _12955_/Y _12959_/Y vssd1 vssd1 vccd1 vccd1 _13109_/C sky130_fd_sc_hd__a21oi_4
XFILLER_180_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15752__C _15968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11911_ _11912_/A _11912_/B _11912_/C _11912_/D vssd1 vssd1 vccd1 vccd1 _11913_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _20673_/B vssd1 vssd1 vccd1 vccd1 _21124_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _23395_/Q vssd1 vssd1 vccd1 vccd1 _19156_/B sky130_fd_sc_hd__buf_2
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11842_ _11840_/X _11841_/Y _12118_/A vssd1 vssd1 vccd1 vccd1 _11846_/A sky130_fd_sc_hd__o21ai_4
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _13228_/X _14532_/X _14557_/X _14560_/X vssd1 vssd1 vccd1 vccd1 _14561_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _12245_/A _11861_/A _11773_/C vssd1 vssd1 vccd1 vccd1 _11774_/B sky130_fd_sc_hd__nand3b_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16300_ _16300_/A vssd1 vssd1 vccd1 vccd1 _16322_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_13_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13512_ _13494_/Y _13507_/Y _13511_/Y vssd1 vssd1 vccd1 vccd1 _13519_/A sky130_fd_sc_hd__a21boi_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _17297_/C vssd1 vssd1 vccd1 vccd1 _17290_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14492_ _14495_/A _14492_/B _14492_/C vssd1 vssd1 vccd1 vccd1 _14493_/B sky130_fd_sc_hd__nand3_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ _16227_/X _16230_/X _16222_/A vssd1 vssd1 vccd1 vccd1 _16234_/A sky130_fd_sc_hd__o21ai_1
XFILLER_16_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13443_ _13443_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _13447_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12185__A _12185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21104__C1 _20966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17859__C1 _17766_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16162_ _16815_/C _16817_/A vssd1 vssd1 vccd1 vccd1 _16638_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12616__C _21039_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13374_ _13783_/B _13802_/A vssd1 vssd1 vccd1 vccd1 _13796_/A sky130_fd_sc_hd__nand2_1
XFILLER_177_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_966 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15113_ _14632_/X _15112_/Y _23364_/Q _14883_/B vssd1 vssd1 vccd1 vccd1 _15233_/A
+ sky130_fd_sc_hd__o211ai_4
X_12325_ _16921_/C vssd1 vssd1 vccd1 vccd1 _16318_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16093_ _16326_/A vssd1 vssd1 vccd1 vccd1 _16093_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15885__A1 _15882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19921_ _23547_/Q _19781_/A _19781_/B _19789_/Y vssd1 vssd1 vccd1 vccd1 _19922_/B
+ sky130_fd_sc_hd__a31o_1
X_15044_ _15041_/Y _15195_/B _15044_/C _15044_/D vssd1 vssd1 vccd1 vccd1 _15045_/B
+ sky130_fd_sc_hd__and4b_1
XANTENNA__19076__A1 _18617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12256_ _12256_/A vssd1 vssd1 vccd1 vccd1 _12260_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19852_ _19480_/X _19659_/Y _19667_/B vssd1 vssd1 vccd1 vccd1 _19863_/C sky130_fd_sc_hd__o21ai_1
XFILLER_96_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22080__B1 _21995_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12187_ _12187_/A _19019_/B vssd1 vssd1 vccd1 vccd1 _12187_/Y sky130_fd_sc_hd__nand2_2
XFILLER_150_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18803_ _18803_/A vssd1 vssd1 vccd1 vccd1 _18844_/C sky130_fd_sc_hd__buf_2
XFILLER_96_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output64_A _14676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19783_ _19783_/A vssd1 vssd1 vccd1 vccd1 _19783_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16995_ _16997_/B _16997_/C _23523_/Q vssd1 vssd1 vccd1 vccd1 _17381_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__22907__A0 _12601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19379__A2 _19800_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18734_ _19279_/A _19280_/A _18731_/X _18732_/Y _18733_/Y vssd1 vssd1 vccd1 vccd1
+ _18738_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_114_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15946_ _15946_/A vssd1 vssd1 vccd1 vccd1 _15946_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15662__C _15662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22383__A1 _13470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18665_ _18669_/C _18669_/D _18665_/C vssd1 vssd1 vccd1 vccd1 _18665_/Y sky130_fd_sc_hd__nand3_4
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _19363_/C _19363_/D _16462_/D vssd1 vssd1 vccd1 vccd1 _15887_/C sky130_fd_sc_hd__and3_2
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21591__C1 _21635_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19431__A _19431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17616_ _17616_/A _17616_/B _17616_/C vssd1 vssd1 vccd1 vccd1 _17656_/A sky130_fd_sc_hd__nand3_1
X_14828_ _14824_/X _14830_/A _14831_/A vssd1 vssd1 vccd1 vccd1 _14828_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_91_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18596_ _18518_/B _18520_/B _18518_/A vssd1 vssd1 vccd1 vccd1 _18619_/A sky130_fd_sc_hd__a21boi_1
XFILLER_184_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19536__C1 _19539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17547_ _17546_/C _17391_/B _17391_/C _17888_/A _19862_/A vssd1 vssd1 vccd1 vccd1
+ _17548_/B sky130_fd_sc_hd__a32o_1
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12623__A1 _20799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14759_ _14886_/C vssd1 vssd1 vccd1 vccd1 _15254_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19551__A2 _18003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17478_ _17277_/Y _17281_/Y _17282_/Y _17287_/Y vssd1 vssd1 vccd1 vccd1 _17478_/X
+ sky130_fd_sc_hd__o211a_2
X_19217_ _19202_/Y _19212_/Y _19216_/Y vssd1 vssd1 vccd1 vccd1 _19217_/X sky130_fd_sc_hd__o21a_1
XFILLER_149_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16429_ _16517_/B _16476_/D vssd1 vssd1 vccd1 vccd1 _16472_/C sky130_fd_sc_hd__nand2_1
XFILLER_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12095__A _12100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14915__A3 _14061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19303__A2 _19172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19148_ _19148_/A _19148_/B _19148_/C vssd1 vssd1 vccd1 vccd1 _19148_/X sky130_fd_sc_hd__and3_1
XANTENNA__17314__A1 _12279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17314__B2 _16741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17865__A2 _18003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19079_ _19069_/Y _19071_/X _18931_/X _18882_/B vssd1 vssd1 vccd1 vccd1 _19079_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21110_ _21159_/A _21228_/A _21110_/C vssd1 vssd1 vccd1 vccd1 _21113_/B sky130_fd_sc_hd__nand3_1
XFILLER_160_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22090_ _22090_/A _22096_/B _22090_/C _22090_/D vssd1 vssd1 vccd1 vccd1 _22093_/A
+ sky130_fd_sc_hd__or4_1
X_21041_ _20940_/B _20929_/Y _20940_/C vssd1 vssd1 vccd1 vccd1 _21045_/B sky130_fd_sc_hd__o21ai_1
XFILLER_113_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18510__A _18511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22992_ _23038_/S vssd1 vssd1 vccd1 vccd1 _23001_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_55_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21871__A _21987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21943_ _21878_/X _21799_/X _21893_/Y vssd1 vssd1 vccd1 vccd1 _21943_/X sky130_fd_sc_hd__o21a_2
XFILLER_55_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16965__A _17388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16053__A1 _12040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14188__C _14188_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21874_ _21874_/A _21874_/B vssd1 vssd1 vccd1 vccd1 _21982_/A sky130_fd_sc_hd__xor2_2
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19698__D _19800_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20137__B1 _17414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20825_ _20676_/B _20821_/X _20955_/A _20673_/A _20955_/C vssd1 vssd1 vccd1 vccd1
+ _20828_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_42_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1011 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11902__A _11902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23544_ _23575_/CLK _23544_/D vssd1 vssd1 vccd1 vccd1 _23544_/Q sky130_fd_sc_hd__dfxtp_1
X_20756_ _20755_/X _20606_/A _20607_/B _20607_/C vssd1 vssd1 vccd1 vccd1 _20756_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_23_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20152__A3 _19539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23475_ _23499_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 _23475_/Q sky130_fd_sc_hd__dfxtp_4
X_20687_ _20533_/B _20670_/A _20676_/A _13053_/X vssd1 vssd1 vccd1 vccd1 _20688_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_195_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_538 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22426_ _22516_/A _22428_/D _22425_/C vssd1 vssd1 vccd1 vccd1 _22427_/C sky130_fd_sc_hd__a21o_1
XANTENNA__17305__A1 _14729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17856__A2 _17465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22357_ _22357_/A _22357_/B vssd1 vssd1 vccd1 vccd1 _22357_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ _12093_/A _19010_/A _19193_/C _16027_/A vssd1 vssd1 vccd1 vccd1 _12110_/Y
+ sky130_fd_sc_hd__nand4b_4
XFILLER_40_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21308_ _21317_/A _21317_/B _21308_/C _21308_/D vssd1 vssd1 vccd1 vccd1 _21308_/Y
+ sky130_fd_sc_hd__nand4_2
X_13090_ _13085_/A _13085_/B _20595_/A _20595_/B vssd1 vssd1 vccd1 vccd1 _13090_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_163_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22288_ _22288_/A _22288_/B vssd1 vssd1 vccd1 vccd1 _22288_/Y sky130_fd_sc_hd__nand2_2
XFILLER_156_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12041_ _12475_/B vssd1 vssd1 vccd1 vccd1 _18941_/B sky130_fd_sc_hd__buf_2
XANTENNA__22062__B1 _13469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13342__A2 _21987_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17608__A2 _16478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21239_ _21015_/X _21012_/X _21140_/C _21154_/Y _21237_/Y vssd1 vssd1 vccd1 vccd1
+ _21240_/B sky130_fd_sc_hd__o311a_1
XANTENNA__22601__A2 _22126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1064 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15800_ _15928_/C _17414_/C _17414_/D _19308_/B vssd1 vssd1 vccd1 vccd1 _15800_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_65_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16780_ _18434_/B _16780_/B vssd1 vssd1 vccd1 vccd1 _17217_/A sky130_fd_sc_hd__nor2_2
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13992_ _13933_/Y _13954_/Y _13991_/Y vssd1 vssd1 vccd1 vccd1 _14005_/A sky130_fd_sc_hd__o21ai_1
XFILLER_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15731_ _15731_/A _15731_/B vssd1 vssd1 vccd1 vccd1 _16805_/A sky130_fd_sc_hd__nand2_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ _12571_/X _13177_/A _12796_/X _12766_/X _13113_/C vssd1 vssd1 vccd1 vccd1
+ _12943_/X sky130_fd_sc_hd__o41a_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18450_ _12311_/A _19859_/A _18462_/A vssd1 vssd1 vccd1 vccd1 _18458_/A sky130_fd_sc_hd__o21ai_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12874_ _20897_/C _12874_/B _13011_/C _12874_/D vssd1 vssd1 vccd1 vccd1 _12875_/A
+ sky130_fd_sc_hd__nand4_1
X_15662_ _15735_/C _15662_/B _15662_/C _15762_/A vssd1 vssd1 vccd1 vccd1 _15920_/A
+ sky130_fd_sc_hd__nor4_4
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16595__A2 _11972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17401_/A _17401_/B vssd1 vssd1 vccd1 vccd1 _17493_/B sky130_fd_sc_hd__nand2_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _23329_/Q vssd1 vssd1 vccd1 vccd1 _21745_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11825_ _11841_/A _18653_/C _12403_/A vssd1 vssd1 vccd1 vccd1 _12118_/A sky130_fd_sc_hd__a21o_2
X_18381_ _18410_/A _18411_/A _18382_/C vssd1 vssd1 vccd1 vccd1 _18383_/A sky130_fd_sc_hd__o21ai_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15593_ _23514_/Q _23515_/Q _23516_/Q _15586_/A hold23/A vssd1 vssd1 vccd1 vccd1
+ _15594_/B sky130_fd_sc_hd__o41a_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18336__A3 _17324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17332_ _17332_/A _17337_/C vssd1 vssd1 vccd1 vccd1 _17336_/A sky130_fd_sc_hd__nand2_1
X_14544_ _14693_/A vssd1 vssd1 vccd1 vccd1 _14544_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_844 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _11823_/A _11823_/B vssd1 vssd1 vccd1 vccd1 _11757_/A sky130_fd_sc_hd__nand2_2
XFILLER_92_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18017__D _18017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17263_ _17586_/A _17587_/A _16056_/X _19543_/B _17454_/B vssd1 vssd1 vccd1 vccd1
+ _17263_/Y sky130_fd_sc_hd__a32oi_2
X_14475_ _14806_/C vssd1 vssd1 vccd1 vccd1 _15044_/C sky130_fd_sc_hd__buf_2
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11687_ _23397_/Q vssd1 vssd1 vccd1 vccd1 _18470_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_186_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19002_ _18439_/X _18440_/X _18657_/C _18788_/A vssd1 vssd1 vccd1 vccd1 _19210_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_186_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13426_ _13323_/X _13338_/X _13354_/C _13354_/B _13394_/Y vssd1 vssd1 vccd1 vccd1
+ _21924_/A sky130_fd_sc_hd__a41o_2
X_16214_ _12018_/X _12020_/X _17753_/A _17753_/B vssd1 vssd1 vccd1 vccd1 _16214_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_139_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17194_ _16952_/Y _17191_/Y _17182_/X _17193_/Y vssd1 vssd1 vccd1 vccd1 _17200_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_128_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16145_ _17741_/A _17742_/A _17055_/A vssd1 vssd1 vccd1 vccd1 _16146_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__20563__C _23457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17847__A2 _17846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13357_ _13354_/Y _22186_/C _13802_/B vssd1 vssd1 vccd1 vccd1 _13357_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12308_ _12308_/A vssd1 vssd1 vccd1 vccd1 _12508_/A sky130_fd_sc_hd__buf_2
XFILLER_115_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19049__A1 _19046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16076_ _16020_/X _16073_/Y _16335_/A _16063_/X vssd1 vssd1 vccd1 vccd1 _16076_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13288_ _13471_/A _13269_/X _13516_/A _13285_/X vssd1 vssd1 vccd1 vccd1 _13288_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_143_969 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19904_ _19900_/X _19903_/X _19899_/Y _19894_/Y vssd1 vssd1 vccd1 vccd1 _19904_/X
+ sky130_fd_sc_hd__o211a_1
X_15027_ _15023_/A _15030_/B _15030_/C vssd1 vssd1 vccd1 vccd1 _15035_/D sky130_fd_sc_hd__a21o_1
X_12239_ _12239_/A vssd1 vssd1 vccd1 vccd1 _16523_/A sky130_fd_sc_hd__buf_4
XFILLER_170_788 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18330__A _18330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23593__D _23593_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_980 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20064__C1 _19800_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19835_ _19835_/A vssd1 vssd1 vccd1 vccd1 _19835_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11895__A2 _17149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16283__A1 _16275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19766_ _19380_/X _19621_/X _19620_/X vssd1 vssd1 vccd1 vccd1 _19932_/B sky130_fd_sc_hd__o21ai_2
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16978_ _16744_/B _16784_/Y _16744_/A vssd1 vssd1 vccd1 vccd1 _16979_/C sky130_fd_sc_hd__a21boi_1
Xinput4 wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18717_ _18717_/A _18717_/B _18717_/C vssd1 vssd1 vccd1 vccd1 _18903_/A sky130_fd_sc_hd__nand3_1
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15929_ _16281_/A _15925_/Y _15923_/X vssd1 vssd1 vccd1 vccd1 _15929_/Y sky130_fd_sc_hd__a21oi_1
X_19697_ _19903_/C _19800_/C _19698_/C _19903_/A vssd1 vssd1 vccd1 vccd1 _19717_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19799__C _19799_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16035__A1 _16032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19161__A _19161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18648_ _23390_/Q _23391_/Q _23392_/Q _23393_/Q vssd1 vssd1 vccd1 vccd1 _19155_/D
+ sky130_fd_sc_hd__nor4_2
XFILLER_188_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17783__A1 _17747_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14597__A1 _15664_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18579_ _18576_/Y _18578_/Y _18573_/Y vssd1 vssd1 vccd1 vccd1 _18579_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20610_ _20610_/A _20765_/A vssd1 vssd1 vccd1 vccd1 _20611_/B sky130_fd_sc_hd__nor2_1
XFILLER_177_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21590_ _21590_/A _21590_/B vssd1 vssd1 vccd1 vccd1 _21602_/A sky130_fd_sc_hd__or2_1
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20541_ _20525_/X _20526_/X _20530_/Y _20533_/Y vssd1 vssd1 vccd1 vccd1 _20548_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_20_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23260_ _23260_/A _23260_/B vssd1 vssd1 vccd1 vccd1 _23261_/A sky130_fd_sc_hd__and2_1
X_20472_ _12871_/A _12872_/A _23450_/Q _12876_/A vssd1 vssd1 vccd1 vccd1 _20621_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_146_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22211_ _22211_/A _22211_/B vssd1 vssd1 vccd1 vccd1 _22211_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23191_ _15662_/C input29/X _23195_/S vssd1 vssd1 vccd1 vccd1 _23192_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_936 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22142_ _22186_/B _22142_/B _22186_/C vssd1 vssd1 vccd1 vccd1 _22267_/A sky130_fd_sc_hd__nand3_4
XFILLER_161_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15864__A _15864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_788 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_619 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22073_ _22073_/A _22073_/B _22073_/C vssd1 vssd1 vccd1 vccd1 _22074_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21024_ _21029_/A _21029_/B _21025_/A vssd1 vssd1 vccd1 vccd1 _21026_/A sky130_fd_sc_hd__a21o_1
XFILLER_99_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22347__A1 _21981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22347__B2 _21981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18015__A2 _18330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22975_ _13228_/X input29/X _22979_/S vssd1 vssd1 vccd1 vccd1 _22976_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21926_ _21920_/X _21922_/Y _21925_/X vssd1 vssd1 vccd1 vccd1 _21938_/A sky130_fd_sc_hd__o21ai_1
XFILLER_28_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11618__A_N _11604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21857_ _21857_/A _21857_/B vssd1 vssd1 vccd1 vccd1 _21858_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11632__A _23598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ _11606_/X _19156_/C _11610_/C vssd1 vssd1 vccd1 vccd1 _11611_/B sky130_fd_sc_hd__nand3b_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20808_ _20819_/A _20819_/B vssd1 vssd1 vccd1 vccd1 _20817_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12590_ _23288_/Q _23286_/Q vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21788_ _21764_/X _21769_/X _21755_/X _21760_/X vssd1 vssd1 vccd1 vccd1 _21875_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_24_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23527_ _23588_/CLK _23527_/D vssd1 vssd1 vccd1 vccd1 _23527_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20739_ _20562_/A _20562_/B _20566_/X vssd1 vssd1 vccd1 vccd1 _20867_/B sky130_fd_sc_hd__o21ba_1
XFILLER_183_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_847 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14260_ _14260_/A _14330_/A vssd1 vssd1 vccd1 vccd1 _14260_/Y sky130_fd_sc_hd__nand2_1
X_23458_ _23571_/CLK hold15/X vssd1 vssd1 vccd1 vccd1 _23458_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21592__C_N _21554_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13211_ _13210_/A _20465_/D _13210_/C vssd1 vssd1 vccd1 vccd1 _13212_/B sky130_fd_sc_hd__a21oi_1
X_22409_ _22409_/A vssd1 vssd1 vccd1 vccd1 _22509_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14191_ _14191_/A _14191_/B _14191_/C vssd1 vssd1 vccd1 vccd1 _15111_/A sky130_fd_sc_hd__nand3_4
XANTENNA__12463__A _19017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23389_ _23389_/CLK _23389_/D vssd1 vssd1 vccd1 vccd1 _23389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13142_ _13141_/A _13141_/B _13141_/C vssd1 vssd1 vccd1 vccd1 _13143_/C sky130_fd_sc_hd__a21o_1
XFILLER_125_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17950_ _17948_/X _18139_/B _17825_/Y vssd1 vssd1 vccd1 vccd1 _17951_/C sky130_fd_sc_hd__a21o_1
XANTENNA__21495__B _21495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ _12911_/Y _12906_/Y _12902_/C vssd1 vssd1 vccd1 vccd1 _13089_/B sky130_fd_sc_hd__o21ai_1
XFILLER_97_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18788__C _19804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16901_ _16911_/A _16904_/A _16900_/Y vssd1 vssd1 vccd1 vccd1 _16901_/Y sky130_fd_sc_hd__o21ai_1
X_12024_ _12024_/A _12024_/B _15718_/A vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__nand3_2
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17881_ _17881_/A _17881_/B _17881_/C vssd1 vssd1 vccd1 vccd1 _17881_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__11877__A2 _11760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19620_ _19620_/A vssd1 vssd1 vccd1 vccd1 _19620_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16832_ _16832_/A _17068_/A vssd1 vssd1 vccd1 vccd1 _16832_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19551_ _19203_/X _18003_/A _19550_/Y vssd1 vssd1 vccd1 vccd1 _19552_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__18006__A2 _17712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16763_ _16763_/A _16763_/B _16763_/C vssd1 vssd1 vccd1 vccd1 _16763_/X sky130_fd_sc_hd__and3_1
X_13975_ _14001_/A _13945_/X _13939_/A _14191_/B vssd1 vssd1 vccd1 vccd1 _13978_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21010__A1 _13202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18502_ _12238_/A _19040_/A _12422_/D vssd1 vssd1 vccd1 vccd1 _18511_/B sky130_fd_sc_hd__o21ai_2
XFILLER_19_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15714_ _16856_/C vssd1 vssd1 vccd1 vccd1 _15798_/A sky130_fd_sc_hd__buf_2
X_19482_ _19482_/A _19482_/B vssd1 vssd1 vccd1 vccd1 _19482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ _21036_/C vssd1 vssd1 vccd1 vccd1 _21050_/D sky130_fd_sc_hd__buf_2
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16694_ _16201_/X _16690_/X _16691_/Y _16693_/Y vssd1 vssd1 vccd1 vccd1 _16706_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18433_ _18433_/A _18433_/B vssd1 vssd1 vccd1 vccd1 _23598_/D sky130_fd_sc_hd__nand2_1
XANTENNA__14579__A1 _15674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15645_ _15645_/A vssd1 vssd1 vccd1 vccd1 _15921_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _20962_/A _13003_/B _20962_/C vssd1 vssd1 vccd1 vccd1 _12858_/B sky130_fd_sc_hd__and3_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19506__A2 _19505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ _18364_/A _18364_/B vssd1 vssd1 vccd1 vccd1 _18364_/Y sky130_fd_sc_hd__nand2_1
X_11808_ _11808_/A vssd1 vssd1 vccd1 vccd1 _16796_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15576_ _23510_/Q _15576_/B vssd1 vssd1 vccd1 vccd1 _23498_/D sky130_fd_sc_hd__xor2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _20894_/A _12788_/B _12915_/A vssd1 vssd1 vccd1 vccd1 _12824_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12054__A2 _12053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _16464_/X _17635_/A _16908_/X _17307_/A vssd1 vssd1 vccd1 vccd1 _17315_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_42_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11739_ _11739_/A _11739_/B vssd1 vssd1 vccd1 vccd1 _11860_/B sky130_fd_sc_hd__nand2_1
X_14527_ _23262_/Q _14520_/X _14526_/X _20583_/A vssd1 vssd1 vccd1 vccd1 _14527_/X
+ sky130_fd_sc_hd__a22o_1
X_18295_ _18295_/A vssd1 vssd1 vccd1 vccd1 _18295_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23588__D _23588_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17246_ _17397_/A _17246_/B _17397_/B vssd1 vssd1 vccd1 vccd1 _17291_/B sky130_fd_sc_hd__and3_1
X_14458_ _14458_/A vssd1 vssd1 vccd1 vccd1 _15233_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__14200__B1 _14089_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1026 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19809__A3 _18461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_903 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13409_ _13613_/A vssd1 vssd1 vccd1 vccd1 _13410_/A sky130_fd_sc_hd__buf_2
XANTENNA__13469__A _13469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13554__A2 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17177_ _17334_/A _17335_/A _17334_/B _17350_/B vssd1 vssd1 vccd1 vccd1 _17181_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_127_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14389_ _14114_/X _13914_/A _14381_/A _14381_/B _14388_/X vssd1 vssd1 vccd1 vccd1
+ _14390_/C sky130_fd_sc_hd__o221ai_1
XANTENNA__12373__A _12373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16128_ _16592_/A vssd1 vssd1 vccd1 vccd1 _16128_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_928 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16059_ _16028_/A _16028_/B _16464_/A _16479_/A vssd1 vssd1 vccd1 vccd1 _16060_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_88_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_6_0_bq_clk_i_A clkbuf_4_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15059__A2 _14933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18995__A _23396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19818_ _19701_/B _19807_/X _19975_/A _20061_/A _20146_/A vssd1 vssd1 vccd1 vccd1
+ _19992_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__11717__A _18945_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14267__B1 _14108_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17107__C _17243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19749_ _19740_/A _19880_/A _19748_/Y vssd1 vssd1 vccd1 vccd1 _19749_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13932__A _15353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22760_ _22701_/B _22707_/A _22762_/B vssd1 vssd1 vccd1 vccd1 _22792_/C sky130_fd_sc_hd__a21oi_1
XFILLER_65_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17756__A1 _12088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_49 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18219__B _19425_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21711_ _21711_/A _21711_/B vssd1 vssd1 vccd1 vccd1 _23555_/D sky130_fd_sc_hd__xnor2_1
X_22691_ _22690_/B _22690_/C _23279_/Q vssd1 vssd1 vccd1 vccd1 _22821_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__20760__B1 _21542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21642_ _21642_/A _21642_/B vssd1 vssd1 vccd1 vccd1 _21643_/B sky130_fd_sc_hd__nand2_1
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15859__A _15859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21573_ _21542_/X _21631_/C _21572_/Y vssd1 vssd1 vccd1 vccd1 _21579_/A sky130_fd_sc_hd__o21ai_1
XFILLER_36_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23312_ _23347_/CLK _23312_/D vssd1 vssd1 vccd1 vccd1 _23312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20524_ _20524_/A vssd1 vssd1 vccd1 vccd1 _20714_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23243_ _23243_/A vssd1 vssd1 vccd1 vccd1 _23439_/D sky130_fd_sc_hd__clkbuf_1
X_20455_ _20455_/A vssd1 vssd1 vccd1 vccd1 _20455_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13098__B _21554_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23174_ _23409_/Q input26/X _23178_/S vssd1 vssd1 vccd1 vccd1 _23175_/A sky130_fd_sc_hd__mux2_1
X_20386_ _20364_/A _20385_/Y _20384_/C vssd1 vssd1 vccd1 vccd1 _20411_/B sky130_fd_sc_hd__o21bai_1
XFILLER_133_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22125_ _22644_/A _13431_/X _22135_/A vssd1 vssd1 vccd1 vccd1 _22130_/C sky130_fd_sc_hd__o21ai_1
XFILLER_133_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13702__C1 _13415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22056_ _22025_/Y _22032_/Y _22035_/X vssd1 vssd1 vccd1 vccd1 _22061_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__22032__A3 _13810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21007_ _20585_/A _20598_/X _21008_/A _20593_/C vssd1 vssd1 vccd1 vccd1 _21007_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_134_1165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17017__C _23522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16856__C _16856_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13760_ _13760_/A _13760_/B vssd1 vssd1 vccd1 vccd1 _21856_/D sky130_fd_sc_hd__and2_2
XFILLER_90_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22958_ _23313_/Q input26/X _22962_/S vssd1 vssd1 vccd1 vccd1 _22959_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12284__A2 _12283_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21909_ _22064_/A _22064_/B _21909_/C vssd1 vssd1 vccd1 vccd1 _21910_/B sky130_fd_sc_hd__and3_1
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12711_ _20799_/A _20639_/D vssd1 vssd1 vccd1 vccd1 _12711_/Y sky130_fd_sc_hd__nor2_2
XFILLER_44_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13691_ _21839_/B _13691_/B vssd1 vssd1 vccd1 vccd1 _13692_/C sky130_fd_sc_hd__nor2_1
XFILLER_188_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22889_ _22895_/A _22889_/B vssd1 vssd1 vccd1 vccd1 _22891_/B sky130_fd_sc_hd__or2_1
XFILLER_102_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15430_ _15430_/A _15430_/B vssd1 vssd1 vccd1 vccd1 _15431_/B sky130_fd_sc_hd__xnor2_1
XFILLER_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12642_ _23286_/Q vssd1 vssd1 vccd1 vccd1 _13011_/D sky130_fd_sc_hd__inv_2
XFILLER_169_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15361_ _14995_/A _14995_/B _15358_/Y _15488_/B vssd1 vssd1 vccd1 vccd1 _15363_/B
+ sky130_fd_sc_hd__a211o_1
X_12573_ _13014_/A vssd1 vssd1 vccd1 vccd1 _20799_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_178_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17100_ _16828_/Y _17091_/Y _17097_/Y _17099_/Y vssd1 vssd1 vccd1 vccd1 _17118_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_15_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14312_ _14386_/A _14312_/B _14312_/C _14312_/D vssd1 vssd1 vccd1 vccd1 _14407_/B
+ sky130_fd_sc_hd__nand4_2
X_18080_ _18080_/A vssd1 vssd1 vccd1 vccd1 _19705_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15292_ _15292_/A _15292_/B vssd1 vssd1 vccd1 vccd1 _15292_/X sky130_fd_sc_hd__or2_1
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17031_ _14631_/X _16668_/B _16780_/B _16918_/Y vssd1 vssd1 vccd1 vccd1 _17032_/B
+ sky130_fd_sc_hd__o211ai_4
X_14243_ _14243_/A _14901_/A _14774_/C vssd1 vssd1 vccd1 vccd1 _14245_/A sky130_fd_sc_hd__nand3_2
XFILLER_109_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15930__B1 _15926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18799__B _18799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14174_ _14174_/A _14174_/B vssd1 vssd1 vccd1 vccd1 _14174_/Y sky130_fd_sc_hd__nand2_2
XFILLER_194_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22008__B1 _22218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13125_ _13125_/A _13125_/B vssd1 vssd1 vccd1 vccd1 _13172_/C sky130_fd_sc_hd__nor2_1
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18982_ _12130_/X _20080_/A _18971_/X _19158_/A _18975_/X vssd1 vssd1 vccd1 vccd1
+ _18983_/C sky130_fd_sc_hd__o221ai_1
XANTENNA__23595__CLK _23598_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _18139_/C vssd1 vssd1 vccd1 vccd1 _17933_/X sky130_fd_sc_hd__clkbuf_2
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13056_ _13056_/A vssd1 vssd1 vccd1 vccd1 _13056_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ _12004_/X _12006_/X _19019_/B _19019_/C vssd1 vssd1 vccd1 vccd1 _12007_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_87_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_972 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater107 _23389_/CLK vssd1 vssd1 vccd1 vccd1 _23385_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__19704__A _19708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17864_ _18604_/A vssd1 vssd1 vccd1 vccd1 _18003_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_120_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater118 _23395_/CLK vssd1 vssd1 vccd1 vccd1 _23416_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18632__C1 _19805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater129 _23378_/CLK vssd1 vssd1 vccd1 vccd1 _23443_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_0_0_bq_clk_i clkbuf_3_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_19603_ _19399_/C _19399_/B _19399_/A vssd1 vssd1 vccd1 vccd1 _19603_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_94_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16815_ _16815_/A _16815_/B _16815_/C _16815_/D vssd1 vssd1 vccd1 vccd1 _16816_/C
+ sky130_fd_sc_hd__nor4_1
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17795_ _17919_/A _17798_/C _17798_/A vssd1 vssd1 vccd1 vccd1 _17795_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19534_ _19534_/A _19534_/B _19534_/C _19534_/D vssd1 vssd1 vccd1 vccd1 _19534_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__17224__A _19662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16746_ _17898_/D vssd1 vssd1 vccd1 vccd1 _18161_/B sky130_fd_sc_hd__clkbuf_2
X_13958_ _14790_/B vssd1 vssd1 vccd1 vccd1 _14795_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13472__B2 _22096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19465_ _19428_/A _19424_/A _19427_/C vssd1 vssd1 vccd1 vccd1 _19465_/X sky130_fd_sc_hd__a21o_1
X_12909_ _12903_/Y _12904_/X _12902_/D vssd1 vssd1 vccd1 vccd1 _12909_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16677_ _16677_/A _16677_/B _16677_/C vssd1 vssd1 vccd1 vccd1 _16904_/A sky130_fd_sc_hd__nand3_2
X_13889_ _13889_/A _14863_/D vssd1 vssd1 vccd1 vccd1 _13890_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18416_ _18411_/X _18415_/Y _18414_/B vssd1 vssd1 vccd1 vccd1 _18417_/C sky130_fd_sc_hd__o21bai_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15628_ _15628_/A vssd1 vssd1 vccd1 vccd1 _15712_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19396_ _19396_/A _19468_/A vssd1 vssd1 vccd1 vccd1 _19402_/A sky130_fd_sc_hd__nand2_1
XFILLER_146_1058 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16782__B _17218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18347_ _18345_/A _18388_/A _18388_/B vssd1 vssd1 vccd1 vccd1 _18348_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15559_ _15559_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15561_/A sky130_fd_sc_hd__nor2_1
XFILLER_187_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18278_ _20317_/A vssd1 vssd1 vccd1 vccd1 _19900_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12815__B _12815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17229_ _17236_/B _17236_/C _17228_/X vssd1 vssd1 vccd1 vccd1 _17232_/B sky130_fd_sc_hd__a21o_1
Xinput40 wb_we_i vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 x[8] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_4
XFILLER_156_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20240_ _20182_/A _20181_/A _20180_/Y vssd1 vssd1 vccd1 vccd1 _20243_/B sky130_fd_sc_hd__o21ai_4
XFILLER_157_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19663__B2 _19859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20171_ _20175_/A _20171_/B _20175_/C vssd1 vssd1 vccd1 vccd1 _20171_/X sky130_fd_sc_hd__and3_1
XFILLER_170_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16229__A1 _16049_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18769__A3 _18617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16229__B2 _19503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17977__A1 _17285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17977__B2 _17465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23136__A _23182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22812_ _22812_/A _22812_/B vssd1 vssd1 vccd1 vccd1 _22859_/A sky130_fd_sc_hd__and2_2
XANTENNA__17134__A _17134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22743_ _22821_/B _22743_/B vssd1 vssd1 vccd1 vccd1 _22747_/A sky130_fd_sc_hd__nand2_2
XFILLER_198_714 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12278__A _16437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16401__A1 _16360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22674_ _22676_/A _22676_/D vssd1 vssd1 vccd1 vccd1 _22675_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21625_ _21625_/A _21625_/B _21625_/C vssd1 vssd1 vccd1 vccd1 _21625_/X sky130_fd_sc_hd__and3_1
XFILLER_166_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_994 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21556_ _21556_/A _21556_/B vssd1 vssd1 vccd1 vccd1 _21590_/B sky130_fd_sc_hd__xnor2_2
XFILLER_193_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20507_ _21169_/A _12695_/A _20663_/C _20663_/D _20506_/X vssd1 vssd1 vccd1 vccd1
+ _20507_/X sky130_fd_sc_hd__a41o_1
XFILLER_5_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21487_ _21487_/A _21487_/B vssd1 vssd1 vccd1 vccd1 _23548_/D sky130_fd_sc_hd__xor2_1
XFILLER_153_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12726__B1 _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23226_ _23432_/Q input16/X _23228_/S vssd1 vssd1 vccd1 vccd1 _23227_/A sky130_fd_sc_hd__mux2_1
X_20438_ _20438_/A _20449_/A _20449_/B vssd1 vssd1 vccd1 vccd1 _20455_/A sky130_fd_sc_hd__and3_1
XFILLER_106_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23157_ _23157_/A vssd1 vssd1 vccd1 vccd1 _23401_/D sky130_fd_sc_hd__clkbuf_1
X_20369_ _20369_/A _20369_/B _20369_/C vssd1 vssd1 vccd1 vccd1 _20369_/X sky130_fd_sc_hd__and3_1
XFILLER_164_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22108_ _22348_/B _22348_/C _22249_/B vssd1 vssd1 vccd1 vccd1 _22108_/X sky130_fd_sc_hd__and3_1
XFILLER_122_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23088_ _23088_/A vssd1 vssd1 vccd1 vccd1 _23370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22039_ _22381_/A _22039_/B _22039_/C vssd1 vssd1 vccd1 vccd1 _22040_/B sky130_fd_sc_hd__nand3_4
X_14930_ _14928_/X _14929_/Y _14814_/B vssd1 vssd1 vccd1 vccd1 _14943_/A sky130_fd_sc_hd__o21ai_1
XFILLER_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input26_A wb_dat_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ _23362_/Q vssd1 vssd1 vccd1 vccd1 _15112_/B sky130_fd_sc_hd__clkinv_2
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16640__A1 _16638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16600_ _16601_/B _16601_/C _11935_/A _16319_/A vssd1 vssd1 vccd1 vccd1 _16600_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_21_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13812_ _13812_/A _13812_/B _13812_/C vssd1 vssd1 vccd1 vccd1 _13813_/A sky130_fd_sc_hd__nand3_1
XFILLER_91_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17580_ _17580_/A _17580_/B vssd1 vssd1 vccd1 vccd1 _17585_/A sky130_fd_sc_hd__nand2_1
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13454__A1 _13552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14792_ _14795_/A _14795_/B _23502_/Q vssd1 vssd1 vccd1 vccd1 _14798_/A sky130_fd_sc_hd__nand3_1
XANTENNA__15115__A_N _23364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16531_ _16531_/A _16558_/A vssd1 vssd1 vccd1 vccd1 _16532_/A sky130_fd_sc_hd__nor2_1
XANTENNA__19185__A3 _19858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13743_ _13743_/A vssd1 vssd1 vccd1 vccd1 _21832_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_188_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19250_ _19069_/A _19069_/B _19069_/C _19071_/X _19249_/X vssd1 vssd1 vccd1 vccd1
+ _19434_/B sky130_fd_sc_hd__a32oi_4
XFILLER_44_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16462_ _19512_/D _16462_/B _16526_/B _16462_/D vssd1 vssd1 vccd1 vccd1 _16462_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13674_ _13674_/A _13680_/C _13680_/D vssd1 vssd1 vccd1 vccd1 _13674_/X sky130_fd_sc_hd__and3_1
X_18201_ _18252_/A _18140_/C _18140_/B _18196_/X vssd1 vssd1 vccd1 vccd1 _18204_/B
+ sky130_fd_sc_hd__o211ai_1
X_15413_ _15413_/A _15413_/B vssd1 vssd1 vccd1 vccd1 _15429_/A sky130_fd_sc_hd__xor2_1
XFILLER_188_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19181_ _19168_/A _19183_/B _19332_/B _19182_/B vssd1 vssd1 vccd1 vccd1 _19188_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_12625_ _23449_/Q vssd1 vssd1 vccd1 vccd1 _20620_/C sky130_fd_sc_hd__buf_2
X_16393_ _16359_/Y _16324_/Y _16381_/Y _16392_/Y vssd1 vssd1 vccd1 vccd1 _16394_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_197_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18132_ _18132_/A _18132_/B _18132_/C vssd1 vssd1 vccd1 vccd1 _18132_/X sky130_fd_sc_hd__or3_1
XFILLER_12_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12556_ _12552_/Y _12555_/X _12557_/A vssd1 vssd1 vccd1 vccd1 _12561_/A sky130_fd_sc_hd__o21bai_1
X_15344_ _15344_/A _15344_/B vssd1 vssd1 vccd1 vccd1 _15345_/A sky130_fd_sc_hd__and2_1
XFILLER_40_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18063_ _17942_/C _17942_/A _23529_/Q vssd1 vssd1 vccd1 vccd1 _18063_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12487_ _12487_/A _12487_/B _12487_/C vssd1 vssd1 vccd1 vccd1 _12536_/A sky130_fd_sc_hd__nand3_2
XFILLER_8_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15275_ _15293_/B _15275_/B _15272_/Y _15294_/A vssd1 vssd1 vccd1 vccd1 _15294_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12717__B1 _12980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17014_ _17014_/A _17014_/B _17014_/C vssd1 vssd1 vccd1 vccd1 _17014_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_output94_A _23268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14226_ _14215_/Y _14218_/Y _14816_/A vssd1 vssd1 vccd1 vccd1 _14228_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__19645__A1 _19504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16459__B2 _16458_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ _14797_/B vssd1 vssd1 vccd1 vccd1 _15019_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16123__A _16123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19137__C _19391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21386__D _21490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13108_ _13109_/A _13109_/B _13109_/C vssd1 vssd1 vccd1 vccd1 _13136_/B sky130_fd_sc_hd__a21o_1
X_18965_ _18969_/C _18969_/D vssd1 vssd1 vccd1 vccd1 _18968_/A sky130_fd_sc_hd__nand2_2
X_14088_ _13948_/X _14029_/C _14863_/A _13901_/B vssd1 vssd1 vccd1 vccd1 _14203_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21204__A1 _12785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17916_ _17916_/A _17916_/B _17916_/C vssd1 vssd1 vccd1 vccd1 _17917_/C sky130_fd_sc_hd__nand3_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _13035_/X _13036_/X _13032_/X _13038_/Y vssd1 vssd1 vccd1 vccd1 _20557_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18896_ _18897_/C _18897_/D _18895_/X vssd1 vssd1 vccd1 vccd1 _18899_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12496__A2 _12181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17847_ _16382_/A _17846_/X _17736_/A vssd1 vssd1 vccd1 vccd1 _17853_/A sky130_fd_sc_hd__o21ai_2
XFILLER_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17778_ _17781_/A _17838_/C _17782_/B _17782_/C vssd1 vssd1 vccd1 vccd1 _17779_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_187_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18992__B _18992_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19517_ _19525_/A _19517_/B vssd1 vssd1 vccd1 vccd1 _19524_/C sky130_fd_sc_hd__nand2_2
X_16729_ _16950_/B _16723_/X _16715_/Y _16720_/Y vssd1 vssd1 vccd1 vccd1 _16735_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__13996__A2 _15353_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19448_ _19778_/D vssd1 vssd1 vccd1 vccd1 _19448_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19379_ _19614_/A _19800_/C _19361_/B vssd1 vssd1 vccd1 vccd1 _19573_/A sky130_fd_sc_hd__a21o_1
XFILLER_72_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12826__A _23454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21410_ _21346_/X _21340_/Y _21247_/X vssd1 vssd1 vccd1 vccd1 _21410_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_187_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22390_ _13470_/A _22461_/A _22283_/X _22567_/A _22386_/Y vssd1 vssd1 vccd1 vccd1
+ _22394_/B sky130_fd_sc_hd__o221ai_1
XFILLER_124_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21341_ _21240_/Y _21246_/X _21340_/Y vssd1 vssd1 vccd1 vccd1 _21341_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21858__B _21858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12971__A3 _12980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21272_ _21273_/A _21274_/C _21274_/A vssd1 vssd1 vccd1 vccd1 _21327_/A sky130_fd_sc_hd__a21o_1
XANTENNA__14760__B _14760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23011_ _23011_/A vssd1 vssd1 vccd1 vccd1 _23336_/D sky130_fd_sc_hd__clkbuf_1
X_20223_ _20219_/X _20220_/Y _20287_/B _20277_/B vssd1 vssd1 vccd1 vccd1 _20223_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_131_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16855__D1 _16856_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20651__C1 _23452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20154_ _20158_/A _20156_/B _20153_/Y vssd1 vssd1 vccd1 vccd1 _20154_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16091__A2_N _16071_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15872__A _18755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20085_ _19951_/B _20043_/A _20083_/Y vssd1 vssd1 vccd1 vccd1 _20159_/C sky130_fd_sc_hd__a21oi_2
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22943__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16622__A1 _11960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15830__C1 _12149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20987_ _21111_/B _20987_/B _21111_/A vssd1 vssd1 vccd1 vccd1 _20994_/B sky130_fd_sc_hd__nand3_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18375__A1 _18376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18375__B2 _20366_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22726_ _22726_/A _22726_/B vssd1 vssd1 vccd1 vccd1 _22750_/A sky130_fd_sc_hd__xnor2_1
XFILLER_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22657_ _22559_/X _22478_/X _22663_/B vssd1 vssd1 vccd1 vccd1 _22657_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_186_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11640__A _16604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ _19155_/B _18469_/B _12410_/C _18998_/C vssd1 vssd1 vccd1 vccd1 _12410_/Y
+ sky130_fd_sc_hd__nand4_4
X_21608_ _21612_/C vssd1 vssd1 vccd1 vccd1 _21608_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13390_ _13602_/C _21902_/C _13354_/C vssd1 vssd1 vccd1 vccd1 _13392_/A sky130_fd_sc_hd__a21o_1
XFILLER_166_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22588_ _22649_/C _22556_/B _22585_/Y _22587_/Y vssd1 vssd1 vccd1 vccd1 _22589_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12455__B _19530_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16689__A1 _16674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12341_ _12337_/Y _12338_/Y _12339_/Y _12340_/X vssd1 vssd1 vccd1 vccd1 _12348_/B
+ sky130_fd_sc_hd__o211ai_1
X_21539_ _21539_/A _21540_/C vssd1 vssd1 vccd1 vccd1 _23549_/D sky130_fd_sc_hd__xnor2_1
XFILLER_194_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15060_ _14809_/Y _14810_/X _14811_/X _14855_/Y _14856_/X vssd1 vssd1 vccd1 vccd1
+ _15060_/X sky130_fd_sc_hd__o32a_1
XFILLER_181_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ _12335_/C _12335_/D vssd1 vssd1 vccd1 vccd1 _12339_/C sky130_fd_sc_hd__nand2_1
XFILLER_5_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14011_ _14077_/C _14011_/B vssd1 vssd1 vccd1 vccd1 _14012_/A sky130_fd_sc_hd__nand2_1
XFILLER_181_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23209_ _15605_/A input8/X _23217_/S vssd1 vssd1 vccd1 vccd1 _23210_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12902__C _12902_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15113__A1 _14632_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23187__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18750_ _18731_/X _18732_/Y _18733_/Y vssd1 vssd1 vccd1 vccd1 _19107_/B sky130_fd_sc_hd__a21oi_2
XFILLER_110_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15962_ _16612_/C vssd1 vssd1 vccd1 vccd1 _17060_/A sky130_fd_sc_hd__buf_2
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16861__B2 _11972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22934__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17701_ _17928_/A _17519_/B _17832_/B vssd1 vssd1 vccd1 vccd1 _17701_/X sky130_fd_sc_hd__a21o_1
XANTENNA__18063__B1 _23529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14913_ _14910_/X _14911_/Y _14912_/X vssd1 vssd1 vccd1 vccd1 _14918_/C sky130_fd_sc_hd__a21o_1
XANTENNA__18602__A2 _12168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18681_ _18681_/A _18681_/B _18681_/C vssd1 vssd1 vccd1 vccd1 _18784_/A sky130_fd_sc_hd__nand3_2
XFILLER_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15893_ _15867_/Y _15888_/Y _15892_/Y vssd1 vssd1 vccd1 vccd1 _16078_/B sky130_fd_sc_hd__a21oi_2
XFILLER_64_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17632_ _17712_/D vssd1 vssd1 vccd1 vccd1 _18016_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14844_ _14844_/A _14844_/B _14844_/C vssd1 vssd1 vccd1 vccd1 _14853_/B sky130_fd_sc_hd__nand3_1
XFILLER_84_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17563_ _17453_/B _17453_/C _17453_/A vssd1 vssd1 vccd1 vccd1 _17563_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_511 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14775_ _13942_/X _14020_/Y _14774_/Y vssd1 vssd1 vccd1 vccd1 _14775_/Y sky130_fd_sc_hd__o21ai_2
X_11987_ _19019_/C _19000_/B vssd1 vssd1 vccd1 vccd1 _11987_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19302_ _19172_/A _19172_/B _19172_/C vssd1 vssd1 vccd1 vccd1 _19302_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ _16480_/X _15698_/A _15698_/B _12379_/X _16479_/X vssd1 vssd1 vccd1 vccd1
+ _16514_/X sky130_fd_sc_hd__o32a_1
XFILLER_32_712 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_572 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13726_ _13730_/C _13730_/A _13730_/B vssd1 vssd1 vccd1 vccd1 _13754_/A sky130_fd_sc_hd__a21o_1
X_17494_ _17493_/A _17493_/B _17493_/C vssd1 vssd1 vccd1 vccd1 _17497_/B sky130_fd_sc_hd__a21o_1
XFILLER_95_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19233_ _19256_/B vssd1 vssd1 vccd1 vccd1 _19233_/Y sky130_fd_sc_hd__inv_2
X_16445_ _16445_/A _16445_/B _16457_/D _17445_/A vssd1 vssd1 vccd1 vccd1 _16446_/B
+ sky130_fd_sc_hd__nand4_1
X_13657_ _13269_/X _13313_/X _13467_/X _13320_/A vssd1 vssd1 vccd1 vccd1 _13665_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16129__B1 _15975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19164_ _19651_/A _19652_/A vssd1 vssd1 vccd1 vccd1 _19838_/A sky130_fd_sc_hd__nand2_4
X_12608_ _23291_/Q vssd1 vssd1 vccd1 vccd1 _12608_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_192_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _19503_/C _17062_/B _16443_/C _16497_/A vssd1 vssd1 vccd1 vccd1 _16457_/B
+ sky130_fd_sc_hd__nand4_2
X_13588_ _13494_/Y _13511_/Y _13507_/Y vssd1 vssd1 vccd1 vccd1 _13590_/B sky130_fd_sc_hd__a21o_1
X_18115_ _18118_/A _18156_/B vssd1 vssd1 vccd1 vccd1 _18298_/A sky130_fd_sc_hd__or2b_1
XFILLER_9_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15327_ _15380_/B _15328_/C _15328_/A vssd1 vssd1 vccd1 vccd1 _15329_/A sky130_fd_sc_hd__a21oi_2
X_19095_ _19107_/B _19107_/C vssd1 vssd1 vccd1 vccd1 _19095_/Y sky130_fd_sc_hd__nand2_1
X_12539_ _18565_/A _12540_/A _12227_/C _12080_/B vssd1 vssd1 vccd1 vccd1 _18571_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_118_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18046_ _17922_/X _17924_/X _17930_/Y _17957_/Y _18129_/A vssd1 vssd1 vccd1 vccd1
+ _18072_/B sky130_fd_sc_hd__o221ai_4
X_15258_ _15303_/A _15265_/A _15262_/A _15303_/D vssd1 vssd1 vccd1 vccd1 _15259_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19148__B _19148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14209_ _15111_/A _15111_/B _15112_/C _14094_/X vssd1 vssd1 vccd1 vccd1 _14764_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_126_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18826__C1 _19029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15189_ _15191_/A _15191_/B _15190_/A _15190_/B vssd1 vssd1 vccd1 vccd1 _15193_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_125_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16301__B1 _16054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19997_ _19987_/Y _19991_/Y _19993_/X vssd1 vssd1 vccd1 vccd1 _19997_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23178__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19164__A _19651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18948_ _18945_/Y _19261_/A _18947_/X vssd1 vssd1 vccd1 vccd1 _18950_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__22302__B _22476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22925__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13130__A3 _12979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18879_ _19073_/A _18781_/B _18882_/A vssd1 vssd1 vccd1 vccd1 _18879_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_94_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20910_ _20900_/Y _20905_/Y _20909_/X vssd1 vssd1 vccd1 vccd1 _20943_/A sky130_fd_sc_hd__a21oi_1
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21890_ _21878_/X _21799_/X _21893_/A _21893_/B vssd1 vssd1 vccd1 vccd1 _21890_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20841_ _20841_/A _20841_/B _20842_/A _20842_/B vssd1 vssd1 vccd1 vccd1 _20841_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23560_ _23571_/CLK _23560_/D vssd1 vssd1 vccd1 vccd1 _23560_/Q sky130_fd_sc_hd__dfxtp_2
X_20772_ _20773_/B _20769_/Y _20775_/A _20775_/D vssd1 vssd1 vccd1 vccd1 _20772_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__16368__B1 _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22511_ _22509_/C _22506_/X _22510_/X vssd1 vssd1 vccd1 vccd1 _22511_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23491_ _23510_/CLK _23503_/Q vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23102__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22442_ _22538_/A _22538_/B _22730_/B vssd1 vssd1 vccd1 vccd1 _22443_/B sky130_fd_sc_hd__nand3_2
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19857__A1 _12279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17317__C1 _17722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20773__A _20773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22373_ _22281_/X _22371_/X _22372_/X _22366_/Y vssd1 vssd1 vccd1 vccd1 _22504_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_136_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_945 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21324_ _21327_/C _21327_/D _21311_/A vssd1 vssd1 vccd1 vccd1 _21324_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21255_ _21255_/A _21353_/A _21345_/C vssd1 vssd1 vccd1 vccd1 _21255_/X sky130_fd_sc_hd__and3_1
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13818__C _21925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11904__A1 _11912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20206_ _20206_/A _20247_/B vssd1 vssd1 vccd1 vccd1 _20207_/C sky130_fd_sc_hd__nand2_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11619__B _12168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21186_ _21186_/A vssd1 vssd1 vccd1 vccd1 _21290_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20137_ _17591_/X _17593_/X _17414_/B _17414_/A _17595_/X vssd1 vssd1 vccd1 vccd1
+ _20137_/Y sky130_fd_sc_hd__o2111ai_1
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22916__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21109__A _21109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20068_ _20160_/A _20071_/C _20071_/A vssd1 vssd1 vccd1 vccd1 _20068_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _11969_/B _11907_/B _11717_/B _12297_/A vssd1 vssd1 vccd1 vccd1 _12251_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22129__C1 _22647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ _13052_/C _13052_/A vssd1 vssd1 vccd1 vccd1 _20673_/B sky130_fd_sc_hd__and2_1
XFILLER_173_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11841_/A _12403_/A vssd1 vssd1 vccd1 vccd1 _11841_/Y sky130_fd_sc_hd__nand2_4
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14560_ input45/X _14549_/X _14693_/A _11677_/X _14559_/X vssd1 vssd1 vccd1 vccd1
+ _14560_/X sky130_fd_sc_hd__a221o_1
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11772_ _11861_/A _18999_/C _12245_/A vssd1 vssd1 vccd1 vccd1 _11774_/A sky130_fd_sc_hd__a21bo_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13555_/A _13511_/B _13555_/B vssd1 vssd1 vccd1 vccd1 _13511_/Y sky130_fd_sc_hd__nand3_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17041__B _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22709_ _22709_/A _22800_/C vssd1 vssd1 vccd1 vccd1 _22709_/Y sky130_fd_sc_hd__nor2_1
XFILLER_198_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14491_ _14298_/C _15446_/C _14377_/C _14495_/A _14492_/B vssd1 vssd1 vccd1 vccd1
+ _14493_/A sky130_fd_sc_hd__a32o_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _16480_/A _16741_/A _16194_/C _16198_/X _16749_/A vssd1 vssd1 vccd1 vccd1
+ _16230_/X sky130_fd_sc_hd__o311a_1
XFILLER_186_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13442_ _13490_/B _13440_/Y _13400_/Y _13482_/A vssd1 vssd1 vccd1 vccd1 _13458_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__21104__B1 _21490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17859__B1 _20055_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_1072 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16161_ _15971_/X _16598_/B _16590_/A _19811_/A _16499_/A vssd1 vssd1 vccd1 vccd1
+ _16641_/B sky130_fd_sc_hd__o2111ai_2
X_13373_ _23325_/Q _13358_/X _22018_/A vssd1 vssd1 vccd1 vccd1 _13802_/A sky130_fd_sc_hd__o21ai_1
XFILLER_186_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15112_ _15112_/A _15112_/B _15112_/C _15112_/D vssd1 vssd1 vccd1 vccd1 _15112_/Y
+ sky130_fd_sc_hd__nand4_2
X_12324_ _12324_/A vssd1 vssd1 vccd1 vccd1 _12324_/X sky130_fd_sc_hd__buf_2
XFILLER_6_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16092_ _16089_/X _16090_/X _16091_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 _16424_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_142_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19920_ _19920_/A _19923_/B vssd1 vssd1 vccd1 vccd1 _19922_/A sky130_fd_sc_hd__nand2_2
XFILLER_170_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15885__A2 _15884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12255_ _12391_/B _12251_/B _12393_/B _12393_/A vssd1 vssd1 vccd1 vccd1 _12300_/B
+ sky130_fd_sc_hd__o211ai_1
X_15043_ _15208_/A _15075_/B _14926_/C _14926_/A _15037_/Y vssd1 vssd1 vccd1 vccd1
+ _15044_/D sky130_fd_sc_hd__a221o_1
XANTENNA__19076__A2 _18928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19851_ _19855_/A _19855_/B _19855_/C vssd1 vssd1 vccd1 vccd1 _19851_/X sky130_fd_sc_hd__and3_1
XFILLER_141_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22080__A1 _21936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19481__C1 _19327_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12186_ _12184_/X _12185_/X _16674_/A vssd1 vssd1 vccd1 vccd1 _12186_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_122_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16834__A1 _15861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18802_ _18802_/A _18802_/B _18802_/C vssd1 vssd1 vccd1 vccd1 _18803_/A sky130_fd_sc_hd__nand3_1
X_19782_ _19625_/A _19447_/B _19625_/D _19768_/Y vssd1 vssd1 vccd1 vccd1 _19782_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_95_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16994_ _16994_/A _17376_/A _16994_/C _16994_/D vssd1 vssd1 vccd1 vccd1 _16997_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22907__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18733_ _18733_/A _18733_/B _18733_/C vssd1 vssd1 vccd1 vccd1 _18733_/Y sky130_fd_sc_hd__nand3_1
XFILLER_23_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15945_ _15725_/Y _15898_/X _16003_/A _15944_/Y vssd1 vssd1 vccd1 vccd1 _16268_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__20918__B1 _12571_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15662__D _15762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12320__A1 _11799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_612 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18664_ _18669_/A _18669_/B vssd1 vssd1 vccd1 vccd1 _18665_/C sky130_fd_sc_hd__nand2_1
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _19700_/D vssd1 vssd1 vccd1 vccd1 _19363_/D sky130_fd_sc_hd__buf_2
XFILLER_37_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _17609_/A _17609_/B _17612_/X _17614_/X vssd1 vssd1 vccd1 vccd1 _17616_/C
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_184_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14827_ _14236_/B _14826_/X _14235_/A vssd1 vssd1 vccd1 vccd1 _14831_/A sky130_fd_sc_hd__o21ai_1
XFILLER_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18595_ _18549_/Y _18547_/C _18554_/B vssd1 vssd1 vccd1 vccd1 _18717_/C sky130_fd_sc_hd__o21ai_1
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19536__B1 _19539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17546_ _17888_/A _17891_/A _17546_/C _19862_/A vssd1 vssd1 vccd1 vccd1 _17838_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14758_ _14886_/A vssd1 vssd1 vccd1 vccd1 _15254_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13709_ _13709_/A _22192_/D _13709_/C _21778_/D vssd1 vssd1 vccd1 vccd1 _13709_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_189_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17477_ _17477_/A _17477_/B vssd1 vssd1 vccd1 vccd1 _17477_/Y sky130_fd_sc_hd__nand2_1
X_14689_ _22968_/D vssd1 vssd1 vccd1 vccd1 _14689_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__23529__CLK _23558_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19216_ _19021_/X _19018_/X _19204_/X vssd1 vssd1 vccd1 vccd1 _19216_/Y sky130_fd_sc_hd__a21oi_2
X_16428_ _16416_/X _16420_/Y _16426_/Y _16427_/X vssd1 vssd1 vccd1 vccd1 _16428_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_165_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19303__A3 _19172_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19147_ _19147_/A _19147_/B vssd1 vssd1 vccd1 vccd1 _19256_/A sky130_fd_sc_hd__nand2_1
XFILLER_158_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16359_ _16396_/B _16397_/B vssd1 vssd1 vccd1 vccd1 _16359_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17314__A2 _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16117__A3 _18172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_956 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19078_ _19073_/Y _18882_/Y _19069_/Y _19071_/X vssd1 vssd1 vccd1 vccd1 _19078_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_173_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_926 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18029_ _17899_/A _17886_/X _17896_/Y vssd1 vssd1 vccd1 vccd1 _18032_/B sky130_fd_sc_hd__a21boi_1
XFILLER_117_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17078__A1 _12509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21040_ _21040_/A _21040_/B vssd1 vssd1 vccd1 vccd1 _21045_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13351__A3 _13349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20082__B1 _20164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14300__A2 _15075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20909__B1 _21054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22991_ _22991_/A vssd1 vssd1 vccd1 vccd1 _23327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14469__C _14469_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21942_ _21890_/X _21894_/X _21936_/Y _21941_/Y vssd1 vssd1 vccd1 vccd1 _21946_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__21871__B _22220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21873_ _21873_/A _22096_/C vssd1 vssd1 vccd1 vccd1 _21874_/B sky130_fd_sc_hd__xor2_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _13056_/X _12936_/A _20823_/Y vssd1 vssd1 vccd1 vccd1 _20828_/B sky130_fd_sc_hd__o21ai_1
XFILLER_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23543_ _23575_/CLK _23543_/D vssd1 vssd1 vccd1 vccd1 _23543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20755_ _13099_/Y _13100_/X _13208_/B _12987_/Y vssd1 vssd1 vccd1 vccd1 _20755_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23474_ _23499_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _23474_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20686_ _20509_/Y _20682_/Y _20678_/Y _20679_/Y vssd1 vssd1 vccd1 vccd1 _20688_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_137_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22425_ _22516_/A _22428_/D _22425_/C vssd1 vssd1 vccd1 vccd1 _22427_/B sky130_fd_sc_hd__nand3_1
XFILLER_148_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17305__A2 _11807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18502__A1 _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22356_ _22356_/A vssd1 vssd1 vccd1 vccd1 _22356_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13327__B1 _22392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21307_ _21307_/A _21307_/B _21386_/B _21307_/D vssd1 vssd1 vccd1 vccd1 _21308_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_108_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22287_ _22289_/C _22289_/D vssd1 vssd1 vccd1 vccd1 _22288_/B sky130_fd_sc_hd__nand2_1
XFILLER_105_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _18481_/C vssd1 vssd1 vccd1 vccd1 _12040_/X sky130_fd_sc_hd__buf_4
XFILLER_46_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21238_ _21154_/Y _21158_/Y _21237_/Y vssd1 vssd1 vccd1 vccd1 _21240_/A sky130_fd_sc_hd__a21oi_1
XFILLER_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13342__A3 _21987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13845__A _22420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21169_ _21169_/A vssd1 vssd1 vccd1 vccd1 _21438_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13991_ _13991_/A _13991_/B vssd1 vssd1 vccd1 vccd1 _13991_/Y sky130_fd_sc_hd__nand2_1
XFILLER_105_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _15864_/A _15729_/X _14553_/X vssd1 vssd1 vccd1 vccd1 _15731_/B sky130_fd_sc_hd__o21ai_4
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12942_ _12627_/X _12654_/A _12604_/Y _21121_/A _13181_/A vssd1 vssd1 vccd1 vccd1
+ _13107_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_86_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _23415_/Q vssd1 vssd1 vccd1 vccd1 _15662_/B sky130_fd_sc_hd__buf_2
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _23293_/Q _23291_/Q _12873_/C _23292_/Q vssd1 vssd1 vccd1 vccd1 _20897_/C
+ sky130_fd_sc_hd__nor4_4
XFILLER_73_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17400_ _17810_/C _17810_/D _17810_/A vssd1 vssd1 vccd1 vccd1 _17401_/B sky130_fd_sc_hd__nand3_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ input43/X _14549_/X _14647_/A _15921_/C vssd1 vssd1 vccd1 vccd1 _14612_/X
+ sky130_fd_sc_hd__a22o_1
X_18380_ _18338_/A _18338_/B _18341_/B vssd1 vssd1 vccd1 vccd1 _18382_/C sky130_fd_sc_hd__o21ai_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11824_ _23389_/Q vssd1 vssd1 vccd1 vccd1 _12403_/A sky130_fd_sc_hd__buf_2
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _23516_/Q _15592_/B vssd1 vssd1 vccd1 vccd1 _23504_/D sky130_fd_sc_hd__xor2_1
XFILLER_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22893__A _22895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17331_/A _17331_/B vssd1 vssd1 vccd1 vccd1 _17337_/C sky130_fd_sc_hd__nor2_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14543_ _23112_/D vssd1 vssd1 vccd1 vccd1 _14693_/A sky130_fd_sc_hd__buf_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11980_/A _11980_/B _11999_/A _12432_/A vssd1 vssd1 vccd1 vccd1 _11760_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17262_ _18607_/A vssd1 vssd1 vccd1 vccd1 _17587_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14474_ _14474_/A _14474_/B _14473_/X vssd1 vssd1 vccd1 vccd1 _14474_/Y sky130_fd_sc_hd__nor3b_1
X_11686_ _12282_/A _11686_/B vssd1 vssd1 vccd1 vccd1 _11686_/Y sky130_fd_sc_hd__nor2_2
X_19001_ _16032_/X _16033_/X _19308_/C _19163_/A vssd1 vssd1 vccd1 vccd1 _19191_/A
+ sky130_fd_sc_hd__o211ai_4
X_16213_ _16213_/A vssd1 vssd1 vccd1 vccd1 _17753_/B sky130_fd_sc_hd__buf_4
XFILLER_146_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13425_ _22521_/A _13810_/B _21883_/C _13600_/C vssd1 vssd1 vccd1 vccd1 _13425_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_128_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17193_ _17187_/A _17187_/B _17192_/X vssd1 vssd1 vccd1 vccd1 _17193_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12924__A _21035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16144_ _16817_/A _16144_/B vssd1 vssd1 vccd1 vccd1 _17055_/A sky130_fd_sc_hd__nand2_1
XFILLER_127_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13356_ _23326_/Q vssd1 vssd1 vccd1 vccd1 _13802_/B sky130_fd_sc_hd__buf_2
XFILLER_6_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12307_ _16526_/D vssd1 vssd1 vccd1 vccd1 _16500_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__19049__A2 _19048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16075_ _15852_/X _16075_/B _16075_/C _16539_/C vssd1 vssd1 vccd1 vccd1 _16335_/A
+ sky130_fd_sc_hd__and4b_2
X_13287_ _13287_/A _13287_/B vssd1 vssd1 vccd1 vccd1 _13303_/A sky130_fd_sc_hd__nor2_1
XFILLER_154_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19903_ _19903_/A _19903_/B _19903_/C vssd1 vssd1 vccd1 vccd1 _19903_/X sky130_fd_sc_hd__and3_1
XFILLER_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15026_ _15077_/A _15030_/B _15030_/C vssd1 vssd1 vccd1 vccd1 _15077_/B sky130_fd_sc_hd__nand3_1
XANTENNA__15954__B _16821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ _12238_/A vssd1 vssd1 vccd1 vccd1 _12238_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18330__B _18373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_992 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19834_ _19939_/A _19876_/B _19833_/X vssd1 vssd1 vccd1 vccd1 _19874_/A sky130_fd_sc_hd__a21o_1
X_12169_ _16856_/B vssd1 vssd1 vccd1 vccd1 _16122_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_150_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11895__A3 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16283__A2 _16278_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19765_ _19771_/B _19771_/C _19763_/X _19764_/Y vssd1 vssd1 vccd1 vccd1 _19928_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_16977_ _16663_/X _16704_/A _17202_/A _16969_/B vssd1 vssd1 vccd1 vccd1 _16979_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_110_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput5 wb_clk_i vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_6
X_18716_ _18714_/Y _18715_/X _18706_/A _18892_/A vssd1 vssd1 vccd1 vccd1 _18717_/B
+ sky130_fd_sc_hd__o211ai_1
X_15928_ _15928_/A _16113_/A _15928_/C _17753_/A vssd1 vssd1 vccd1 vccd1 _16281_/A
+ sky130_fd_sc_hd__nand4_4
X_19696_ _19698_/A vssd1 vssd1 vccd1 vccd1 _19903_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16035__A2 _16033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18647_ _18647_/A _18647_/B _18647_/C vssd1 vssd1 vccd1 vccd1 _18669_/D sky130_fd_sc_hd__nand3_4
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15859_ _15859_/A _15859_/B _15859_/C vssd1 vssd1 vccd1 vccd1 _15879_/B sky130_fd_sc_hd__nand3_2
XANTENNA__19161__B _19651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18578_ _12546_/B _18571_/Y _19090_/B _19090_/C vssd1 vssd1 vccd1 vccd1 _18578_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_178_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17529_ _23526_/Q _17529_/B vssd1 vssd1 vccd1 vccd1 _17534_/A sky130_fd_sc_hd__xnor2_1
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11804__B1 _19123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23069__A0 _14621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20540_ _20542_/A _20542_/B _20542_/C _20547_/C vssd1 vssd1 vccd1 vccd1 _20540_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_137_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20471_ _21493_/A _21493_/B vssd1 vssd1 vccd1 vccd1 _20471_/Y sky130_fd_sc_hd__nand2_2
X_22210_ _22215_/A _22215_/B _22177_/Y _22195_/Y _22200_/Y vssd1 vssd1 vccd1 vccd1
+ _22210_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_192_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23190_ _23190_/A vssd1 vssd1 vccd1 vccd1 _23415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13309__B1 _23323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15849__A2 _15975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22141_ _22141_/A _22141_/B _22141_/C _22141_/D vssd1 vssd1 vccd1 vccd1 _22186_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_134_948 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22072_ _21940_/B _21912_/A _21934_/Y _21933_/X vssd1 vssd1 vccd1 vccd1 _22073_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_126_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22043__A _22043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21023_ _23563_/Q vssd1 vssd1 vccd1 vccd1 _21025_/A sky130_fd_sc_hd__inv_2
XFILLER_114_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17137__A _19323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18015__A3 _17889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22974_ _22974_/A vssd1 vssd1 vccd1 vccd1 _23319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21925_ _22510_/A _21925_/B _22510_/C vssd1 vssd1 vccd1 vccd1 _21925_/X sky130_fd_sc_hd__and3_1
XFILLER_56_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21856_ _21856_/A _21856_/B _21856_/C _21856_/D vssd1 vssd1 vccd1 vccd1 _21857_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _20819_/A _20819_/B _20809_/A _20809_/B vssd1 vssd1 vccd1 vccd1 _20812_/A
+ sky130_fd_sc_hd__nand4_1
X_21787_ _13794_/Y _21785_/Y _13813_/A _21786_/Y vssd1 vssd1 vccd1 vccd1 _21789_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_24_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17600__A _17600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23526_ _23538_/CLK _23526_/D vssd1 vssd1 vccd1 vccd1 _23526_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20738_ _20738_/A vssd1 vssd1 vccd1 vccd1 _20867_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_bq_clk_i clkbuf_4_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _23584_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_196_686 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22218__A _22218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23040__C input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23457_ _23571_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 _23457_/Q sky130_fd_sc_hd__dfxtp_1
X_20669_ _20669_/A _21124_/B _20669_/C _20962_/B vssd1 vssd1 vccd1 vccd1 _20669_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_195_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13210_ _13210_/A _20465_/D _13210_/C vssd1 vssd1 vccd1 vccd1 _20611_/A sky130_fd_sc_hd__and3_1
XFILLER_51_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18487__B1 _18474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22408_ _22504_/B vssd1 vssd1 vccd1 vccd1 _22410_/A sky130_fd_sc_hd__inv_2
XFILLER_167_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ _14199_/A _14094_/A _23360_/Q vssd1 vssd1 vccd1 vccd1 _14886_/A sky130_fd_sc_hd__a21o_2
XFILLER_164_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23388_ _23391_/CLK _23388_/D vssd1 vssd1 vccd1 vccd1 _23388_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_125_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13141_ _13141_/A _13141_/B _13141_/C vssd1 vssd1 vccd1 vccd1 _13143_/B sky130_fd_sc_hd__nand3_1
XFILLER_174_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22339_ _22234_/A _22234_/B _22234_/C _22228_/Y _22238_/X vssd1 vssd1 vccd1 vccd1
+ _22341_/A sky130_fd_sc_hd__a32oi_2
XANTENNA__18431__A _23538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13072_ _13078_/A _13078_/B _13079_/B vssd1 vssd1 vccd1 vccd1 _13072_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16900_ _16900_/A _16900_/B vssd1 vssd1 vccd1 vccd1 _16900_/Y sky130_fd_sc_hd__nand2_1
X_12023_ _12021_/Y _12022_/X _11866_/Y vssd1 vssd1 vccd1 vccd1 _12023_/Y sky130_fd_sc_hd__a21oi_2
X_17880_ _17880_/A _17880_/B _17880_/C _17999_/A vssd1 vssd1 vccd1 vccd1 _17881_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_104_171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11877__A3 _11760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16831_ _16832_/A _17068_/A _16830_/X vssd1 vssd1 vccd1 vccd1 _16831_/X sky130_fd_sc_hd__a21o_1
XFILLER_66_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19550_ _19547_/X _19537_/X _19542_/X vssd1 vssd1 vccd1 vccd1 _19550_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__15790__A _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16762_ _16582_/C _16351_/Y _16283_/Y _16761_/Y vssd1 vssd1 vccd1 vccd1 _16762_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18006__A3 _17712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13974_ _14797_/C vssd1 vssd1 vccd1 vccd1 _13985_/D sky130_fd_sc_hd__buf_2
XFILLER_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18501_ _11760_/A _11760_/B _15882_/X _16604_/X _18500_/X vssd1 vssd1 vccd1 vccd1
+ _18501_/X sky130_fd_sc_hd__o32a_1
XFILLER_111_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15713_ _15713_/A _15713_/B _15713_/C vssd1 vssd1 vccd1 vccd1 _16856_/C sky130_fd_sc_hd__nand3_4
X_19481_ _18476_/X _18484_/X _19846_/A _19327_/B vssd1 vssd1 vccd1 vccd1 _19482_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_62_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12925_ _21050_/C vssd1 vssd1 vccd1 vccd1 _13156_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16693_ _16693_/A _16900_/B vssd1 vssd1 vccd1 vccd1 _16693_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18432_ _18420_/X _18425_/Y _18430_/Y _18431_/X vssd1 vssd1 vccd1 vccd1 _18433_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_62_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15644_ _15644_/A vssd1 vssd1 vccd1 vccd1 _15644_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _12725_/A _12854_/Y _12855_/Y _12728_/B vssd1 vssd1 vccd1 vccd1 _12858_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _23533_/Q vssd1 vssd1 vccd1 vccd1 _18363_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11807_ _11625_/A _11711_/B _11711_/C _11708_/Y vssd1 vssd1 vccd1 vccd1 _11807_/X
+ sky130_fd_sc_hd__a31o_4
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _15577_/A _23508_/Q _23509_/Q _15586_/C vssd1 vssd1 vccd1 vccd1 _15576_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _12824_/A vssd1 vssd1 vccd1 vccd1 _13119_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17314_ _12279_/X _17230_/A _12323_/X _16741_/A vssd1 vssd1 vccd1 vccd1 _17314_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14546_/A vssd1 vssd1 vccd1 vccd1 _14526_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18294_ _18244_/A _18245_/C _18293_/B vssd1 vssd1 vccd1 vccd1 _18305_/B sky130_fd_sc_hd__o21a_1
XFILLER_109_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11738_ _11918_/A vssd1 vssd1 vccd1 vccd1 _11738_/X sky130_fd_sc_hd__buf_4
XFILLER_159_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17245_ _17397_/A _17239_/X _17397_/B vssd1 vssd1 vccd1 vccd1 _17291_/A sky130_fd_sc_hd__a21oi_1
X_14457_ _14457_/A vssd1 vssd1 vccd1 vccd1 _14469_/C sky130_fd_sc_hd__clkbuf_2
X_11669_ _11669_/A vssd1 vssd1 vccd1 vccd1 _19203_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1038 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13408_ _13796_/A _13796_/B vssd1 vssd1 vccd1 vccd1 _13613_/A sky130_fd_sc_hd__nand2_1
X_17176_ _17179_/A _17179_/B _17179_/C vssd1 vssd1 vccd1 vccd1 _17350_/B sky130_fd_sc_hd__nand3_1
XFILLER_116_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14388_ _13972_/X _14458_/A _13985_/D _14246_/A _14876_/B vssd1 vssd1 vccd1 vccd1
+ _14388_/X sky130_fd_sc_hd__a32o_1
XFILLER_155_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16127_ _17712_/A _17092_/A _16314_/B _16314_/C vssd1 vssd1 vccd1 vccd1 _16592_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_143_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13339_ _13339_/A vssd1 vssd1 vccd1 vccd1 _13339_/X sky130_fd_sc_hd__buf_2
XFILLER_143_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16058_ _16058_/A vssd1 vssd1 vccd1 vccd1 _16479_/A sky130_fd_sc_hd__buf_2
XANTENNA__15700__A1 _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19156__B _19156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15009_ _14976_/Y _14979_/X _14987_/Y vssd1 vssd1 vccd1 vccd1 _15013_/A sky130_fd_sc_hd__o21ai_1
XFILLER_142_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21785__B1 _13797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19817_ _19803_/X _17763_/X _19815_/A vssd1 vssd1 vccd1 vccd1 _19992_/A sky130_fd_sc_hd__o21ai_1
XFILLER_110_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11717__B _11717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16796__A _16796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19172__A _19172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19748_ _19880_/B _19893_/B vssd1 vssd1 vccd1 vccd1 _19748_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13932__B _15353_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19679_ _19654_/X _19658_/Y _19672_/Y _19678_/Y vssd1 vssd1 vccd1 vccd1 _19688_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18953__A1 _11834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11733__A _23586_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19900__A _19900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21710_ _21723_/B _21723_/D vssd1 vssd1 vccd1 vccd1 _21711_/B sky130_fd_sc_hd__nand2_1
X_22690_ _23279_/Q _22690_/B _22690_/C vssd1 vssd1 vccd1 vccd1 _22818_/C sky130_fd_sc_hd__nand3b_1
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21641_ _21598_/A _21641_/B _21641_/C vssd1 vssd1 vccd1 vccd1 _21642_/B sky130_fd_sc_hd__nand3b_1
XFILLER_24_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17420__A _19949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21572_ _21570_/A _21569_/Y _21614_/C vssd1 vssd1 vccd1 vccd1 _21572_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1078 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20523_ _20523_/A _20523_/B _20523_/C vssd1 vssd1 vccd1 vccd1 _20524_/A sky130_fd_sc_hd__nand3_1
X_23311_ _23343_/CLK _23311_/D vssd1 vssd1 vccd1 vccd1 _23311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20454_ _20419_/X _20440_/Y _20453_/Y _20438_/A vssd1 vssd1 vccd1 vccd1 _20454_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_193_678 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23242_ _23439_/Q input24/X _23250_/S vssd1 vssd1 vccd1 vccd1 _23243_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_892 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15875__A _18755_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23173_ _23173_/A vssd1 vssd1 vccd1 vccd1 _23408_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13950__B1 _14188_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20815__A2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20385_ _20337_/A _20298_/A _20337_/C vssd1 vssd1 vccd1 vccd1 _20385_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13098__C _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17141__B1 _17898_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22124_ _21996_/Y _22122_/Y _22123_/Y _13410_/X vssd1 vssd1 vccd1 vccd1 _22135_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22055_ _22015_/X _22016_/X _22036_/X _22044_/Y _22197_/A vssd1 vssd1 vccd1 vccd1
+ _22208_/A sky130_fd_sc_hd__o221ai_4
XANTENNA__21776__B1 _21744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21006_ _20859_/Y _21004_/X _21005_/Y vssd1 vssd1 vccd1 vccd1 _21006_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_82_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19082__A _19082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12269__B1 _12093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19197__A1 _12053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22220__B _22263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21117__A _21159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16856__D _16856_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22957_ _22957_/A vssd1 vssd1 vccd1 vccd1 _23312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12710_ _12709_/X _12648_/X _12661_/A vssd1 vssd1 vccd1 vccd1 _12718_/A sky130_fd_sc_hd__o21ai_1
X_21908_ _21896_/A _22040_/A _22043_/A vssd1 vssd1 vccd1 vccd1 _21913_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13690_ _13743_/A _22713_/C _13864_/A vssd1 vssd1 vccd1 vccd1 _13691_/B sky130_fd_sc_hd__a21oi_1
XFILLER_70_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22888_ _22887_/B _22887_/C _23446_/Q vssd1 vssd1 vccd1 vccd1 _22889_/B sky130_fd_sc_hd__a21boi_1
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ _23288_/Q _23287_/Q vssd1 vssd1 vccd1 vccd1 _13011_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21839_ _21839_/A _21839_/B vssd1 vssd1 vccd1 vccd1 _21840_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_787 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15360_ _14184_/A _14184_/B _15357_/X _15358_/Y _15536_/A vssd1 vssd1 vccd1 vccd1
+ _15360_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ _23301_/Q vssd1 vssd1 vccd1 vccd1 _13014_/A sky130_fd_sc_hd__clkinv_2
XFILLER_184_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14311_ _14310_/A _14310_/C _14310_/D _14310_/B vssd1 vssd1 vccd1 vccd1 _14311_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23509_ _23518_/CLK input45/X vssd1 vssd1 vccd1 vccd1 _23509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15291_ _15291_/A _15291_/B vssd1 vssd1 vccd1 vccd1 _23276_/D sky130_fd_sc_hd__nor2_1
XANTENNA__15915__D1 _17098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17030_ _16781_/B _16665_/X _17029_/X _23428_/Q vssd1 vssd1 vccd1 vccd1 _17032_/A
+ sky130_fd_sc_hd__o211ai_2
X_14242_ _14459_/A _15082_/D _15415_/A _14377_/A vssd1 vssd1 vccd1 vccd1 _14256_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19657__C1 _19525_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14173_ _14173_/A _14173_/B _14384_/A vssd1 vssd1 vccd1 vccd1 _14174_/B sky130_fd_sc_hd__nand3_2
XANTENNA__17132__B1 _17303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22008__A1 _22218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13124_ _13133_/D _13124_/B _13124_/C vssd1 vssd1 vccd1 vccd1 _13125_/B sky130_fd_sc_hd__and3_1
XFILLER_194_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18981_ _18981_/A vssd1 vssd1 vccd1 vccd1 _19158_/A sky130_fd_sc_hd__clkbuf_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ _17932_/A _17932_/B vssd1 vssd1 vccd1 vccd1 _18139_/C sky130_fd_sc_hd__nand2_1
XFILLER_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13055_ _12828_/Y _20529_/A _13051_/X _13054_/Y vssd1 vssd1 vccd1 vccd1 _13055_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16238__A2 _15926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ _16033_/A vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__buf_4
X_17863_ _17863_/A _17863_/B vssd1 vssd1 vccd1 vccd1 _17880_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater108 _23298_/CLK vssd1 vssd1 vccd1 vccd1 _23297_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18632__B1 _18439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14249__A1 _14433_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater119 _23396_/CLK vssd1 vssd1 vccd1 vccd1 _23395_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19602_ _19600_/Y _19601_/X _19598_/Y _19609_/B vssd1 vssd1 vccd1 vccd1 _19605_/B
+ sky130_fd_sc_hd__o211ai_1
X_16814_ _16814_/A vssd1 vssd1 vccd1 vccd1 _16814_/X sky130_fd_sc_hd__clkbuf_2
X_17794_ _17792_/A _17792_/B _17792_/C vssd1 vssd1 vccd1 vccd1 _17919_/A sky130_fd_sc_hd__a21o_1
XFILLER_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19533_ _19534_/D _19532_/X _18673_/X _18096_/A vssd1 vssd1 vccd1 vccd1 _19533_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_16745_ _16745_/A vssd1 vssd1 vccd1 vccd1 _17898_/D sky130_fd_sc_hd__buf_2
X_13957_ _23501_/Q vssd1 vssd1 vccd1 vccd1 _14790_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18935__A1 _11875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1098 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19464_ _19116_/C _19425_/X _19428_/A _19424_/A _19116_/A vssd1 vssd1 vccd1 vccd1
+ _19464_/Y sky130_fd_sc_hd__o2111ai_1
X_12908_ _12908_/A _12908_/B _12908_/C vssd1 vssd1 vccd1 vccd1 _13101_/C sky130_fd_sc_hd__nand3_2
X_16676_ _15910_/X _16911_/A _16214_/Y vssd1 vssd1 vccd1 vccd1 _16676_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__20742__A1 _21455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13888_ _14863_/C _14024_/B vssd1 vssd1 vccd1 vccd1 _13889_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18415_ _18350_/A _18394_/A _18393_/B vssd1 vssd1 vccd1 vccd1 _18415_/Y sky130_fd_sc_hd__a21boi_1
X_15627_ _15618_/X _15621_/X _15652_/A vssd1 vssd1 vccd1 vccd1 _15797_/A sky130_fd_sc_hd__o21ai_4
X_19395_ _19389_/A _19389_/B _19389_/C _19355_/Y vssd1 vssd1 vccd1 vccd1 _19396_/A
+ sky130_fd_sc_hd__a31oi_1
X_12839_ _12836_/A _12836_/B _12770_/C _12845_/C vssd1 vssd1 vccd1 vccd1 _12988_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18346_ _18346_/A vssd1 vssd1 vccd1 vccd1 _18388_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17240__A _19949_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15558_ _15558_/A _15558_/B _15558_/C vssd1 vssd1 vccd1 vccd1 _15559_/B sky130_fd_sc_hd__nor3_4
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19360__A1 _12324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14509_ _16167_/C vssd1 vssd1 vccd1 vccd1 _16549_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_187_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18277_ _18274_/X _20317_/A _18277_/C _18277_/D vssd1 vssd1 vccd1 vccd1 _18277_/X
+ sky130_fd_sc_hd__and4b_1
X_15489_ _15446_/D _15369_/A _15369_/B _15533_/A _15420_/C vssd1 vssd1 vccd1 vccd1
+ _15489_/X sky130_fd_sc_hd__a32o_1
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14185__B1 _15175_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17228_ _11971_/X _11972_/X _15612_/A _15612_/B vssd1 vssd1 vccd1 vccd1 _17228_/X
+ sky130_fd_sc_hd__a22o_2
Xinput30 wb_dat_i[30] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_4
Xinput41 x[0] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_4
Xinput52 x[9] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_4
XANTENNA__19112__A1 _18941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12735__A1 _12634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17159_ _17179_/B vssd1 vssd1 vccd1 vccd1 _17350_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_851 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20170_ _20175_/A _20283_/B _20175_/C vssd1 vssd1 vccd1 vccd1 _20170_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20106__A _20106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11728__A _16661_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16229__A2 _17625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17977__A2 _18096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15988__A1 _15858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22811_ _22808_/B _22808_/C _22810_/Y _22808_/A vssd1 vssd1 vccd1 vccd1 _22812_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_72_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17134__B _17134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14660__A1 _18434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14660__B2 _16780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22742_ _22820_/A vssd1 vssd1 vccd1 vccd1 _22743_/B sky130_fd_sc_hd__inv_2
XFILLER_164_1104 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16401__A2 _15884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22673_ _22549_/A _22549_/B _22598_/A vssd1 vssd1 vccd1 vccd1 _22676_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__11613__D _12308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20495__B _23297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21624_ _21624_/A _21624_/B vssd1 vssd1 vccd1 vccd1 _21660_/C sky130_fd_sc_hd__nor2_1
XFILLER_194_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20497__B1 _23297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21555_ _21555_/A _21555_/B vssd1 vssd1 vccd1 vccd1 _21556_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22238__A1 _22237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20506_ _12644_/X _12711_/Y _12763_/A _12714_/A vssd1 vssd1 vccd1 vccd1 _20506_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_154_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21486_ _21418_/Y _21422_/B _21413_/X _21409_/X vssd1 vssd1 vccd1 vccd1 _21487_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20437_ _20452_/B _20452_/C _20452_/A vssd1 vssd1 vccd1 vccd1 _20449_/B sky130_fd_sc_hd__a21o_1
XFILLER_10_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23225_ _23225_/A vssd1 vssd1 vccd1 vccd1 _23431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16468__A2 _16539_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20368_ _20368_/A _20368_/B _20368_/C _20368_/D vssd1 vssd1 vccd1 vccd1 _20371_/A
+ sky130_fd_sc_hd__or4_1
X_23156_ _23401_/Q input17/X _23156_/S vssd1 vssd1 vccd1 vccd1 _23157_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11638__A _16591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22107_ _22107_/A _22107_/B _22107_/C _22107_/D vssd1 vssd1 vccd1 vccd1 _22249_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19805__A _19805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23087_ _23370_/Q input19/X _23095_/S vssd1 vssd1 vccd1 vccd1 _23088_/A sky130_fd_sc_hd__mux2_1
X_20299_ _20293_/X _20294_/X _20343_/A vssd1 vssd1 vccd1 vccd1 _20300_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22038_ _22038_/A vssd1 vssd1 vccd1 vccd1 _22153_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14860_ _23361_/Q _23360_/Q _15111_/A _15111_/B vssd1 vssd1 vccd1 vccd1 _14860_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_57_76 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13811_ _13616_/A _13616_/B _13810_/Y _13620_/X vssd1 vssd1 vccd1 vccd1 _13812_/C
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__16640__A2 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A wb_dat_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ _14798_/B _14791_/B _14791_/C vssd1 vssd1 vccd1 vccd1 _14791_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__22174__B1 _22276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16530_ _16530_/A _16530_/B _16530_/C vssd1 vssd1 vccd1 vccd1 _16531_/A sky130_fd_sc_hd__nand3_4
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13742_ _13563_/X _13741_/X _22192_/C _13582_/B vssd1 vssd1 vccd1 vccd1 _13744_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_64 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16461_ _16452_/Y _16453_/X _16404_/A _16405_/A vssd1 vssd1 vccd1 vccd1 _16467_/B
+ sky130_fd_sc_hd__o211ai_1
X_13673_ _13673_/A vssd1 vssd1 vccd1 vccd1 _13680_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13206__A2 _20464_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18200_ _18122_/Y _18192_/Y _18154_/X _18302_/C _18195_/Y vssd1 vssd1 vccd1 vccd1
+ _18200_/X sky130_fd_sc_hd__o221a_1
X_15412_ _15412_/A _15412_/B vssd1 vssd1 vccd1 vccd1 _15413_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19180_ _19969_/A _19180_/B _19180_/C _19180_/D vssd1 vssd1 vccd1 vccd1 _19332_/B
+ sky130_fd_sc_hd__and4_2
XANTENNA__22477__A1 _21997_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12624_ _12687_/B vssd1 vssd1 vccd1 vccd1 _12624_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16392_ _16383_/X _16386_/X _16324_/Y _16391_/Y vssd1 vssd1 vccd1 vccd1 _16392_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_197_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18131_ _18122_/Y _18127_/Y _18155_/A vssd1 vssd1 vccd1 vccd1 _18136_/A sky130_fd_sc_hd__o21ai_1
XFILLER_106_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17889__D1 _17723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15343_ _15478_/A _15442_/B _15442_/D vssd1 vssd1 vccd1 vccd1 _15344_/B sky130_fd_sc_hd__o21ai_1
XFILLER_169_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12555_ _12553_/X _12554_/Y _12540_/B _18565_/A vssd1 vssd1 vccd1 vccd1 _12555_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater158_A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18062_ _23528_/Q _17828_/A _17828_/B _17951_/C _17946_/X vssd1 vssd1 vccd1 vccd1
+ _18062_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_11_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15274_ _15293_/B _15275_/B _15272_/Y _15294_/A vssd1 vssd1 vccd1 vccd1 _15276_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_156_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12486_ _12199_/A _12198_/B _12218_/Y _12217_/X vssd1 vssd1 vccd1 vccd1 _12487_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_156_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17013_ _23520_/Q _17006_/Y _17008_/Y _17012_/Y vssd1 vssd1 vccd1 vccd1 _17014_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_22_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14225_ _14227_/A _14227_/B _14215_/Y _14218_/Y _14816_/A vssd1 vssd1 vccd1 vccd1
+ _14229_/C sky130_fd_sc_hd__o221ai_2
XFILLER_172_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19645__A2 _19505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12932__A _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output87_A _23581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14156_ _14230_/A _14156_/B _14156_/C vssd1 vssd1 vccd1 vccd1 _14302_/B sky130_fd_sc_hd__nand3_2
XFILLER_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _13107_/A _13107_/B _13107_/C vssd1 vssd1 vccd1 vccd1 _13109_/A sky130_fd_sc_hd__nand3_1
XFILLER_112_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ _18964_/A _18964_/B _19410_/B vssd1 vssd1 vccd1 vccd1 _18969_/D sky130_fd_sc_hd__nand3_2
XFILLER_112_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _23355_/Q vssd1 vssd1 vccd1 vccd1 _14863_/A sky130_fd_sc_hd__buf_4
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _17915_/A vssd1 vssd1 vccd1 vccd1 _17917_/B sky130_fd_sc_hd__inv_2
XFILLER_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21204__A2 _12862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13031_/Y _13037_/Y _13030_/Y vssd1 vssd1 vccd1 vccd1 _13038_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_67_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18895_ _18904_/A _18904_/B vssd1 vssd1 vccd1 vccd1 _18895_/X sky130_fd_sc_hd__and2_1
XANTENNA__12496__A3 _12181_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17235__A _17235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17846_ _17975_/A vssd1 vssd1 vccd1 vccd1 _17846_/X sky130_fd_sc_hd__buf_2
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20963__A1 _21545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17777_ _17776_/Y _17656_/C _17656_/A vssd1 vssd1 vccd1 vccd1 _17779_/B sky130_fd_sc_hd__o21ai_1
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14989_ _14889_/A _14889_/B _15001_/A vssd1 vssd1 vccd1 vccd1 _15099_/A sky130_fd_sc_hd__a21o_1
XFILLER_47_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19516_ _19525_/A _19525_/B _19524_/B vssd1 vssd1 vccd1 vccd1 _19519_/C sky130_fd_sc_hd__nand3_1
XFILLER_34_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_743 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16728_ _16262_/X _16260_/Y _16268_/D vssd1 vssd1 vccd1 vccd1 _16732_/B sky130_fd_sc_hd__o21ai_1
XFILLER_81_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19447_ _19447_/A _19447_/B vssd1 vssd1 vccd1 vccd1 _19778_/D sky130_fd_sc_hd__nand2_1
X_16659_ _15932_/A _16665_/A _23427_/Q vssd1 vssd1 vccd1 vccd1 _17722_/A sky130_fd_sc_hd__o21bai_4
XFILLER_90_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19378_ _19534_/B vssd1 vssd1 vccd1 vccd1 _19800_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__19333__A1 _11926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19333__B2 _19482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18329_ _20265_/A vssd1 vssd1 vccd1 vccd1 _20368_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21340_ _21340_/A _21340_/B vssd1 vssd1 vccd1 vccd1 _21340_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17895__A1 _20217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21271_ _21387_/C _21271_/B vssd1 vssd1 vccd1 vccd1 _21274_/A sky130_fd_sc_hd__nand2_1
XFILLER_191_968 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16314__A _19161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22035__B _22392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20222_ _20222_/A vssd1 vssd1 vccd1 vccd1 _20287_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17647__A1 _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23010_ _23336_/Q input16/X _23012_/S vssd1 vssd1 vccd1 vccd1 _23011_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16855__C1 _16856_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20153_ _20158_/C _20158_/D vssd1 vssd1 vccd1 vccd1 _20153_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23147__A _23169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20084_ _12237_/X _20263_/A _20164_/B _20043_/A _20083_/Y vssd1 vssd1 vccd1 vccd1
+ _20086_/A sky130_fd_sc_hd__o311a_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1008 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16083__B1 _16062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16622__A2 _23595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12289__A _12289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15830__B1 _18481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19021__B1 _12464_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ _20846_/A _20847_/A _20847_/B vssd1 vssd1 vccd1 vccd1 _20986_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_129_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22725_ _22725_/A _22725_/B vssd1 vssd1 vccd1 vccd1 _22726_/B sky130_fd_sc_hd__nand2_1
XFILLER_198_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16386__A1 _16377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23585__CLK _23588_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22656_ _22656_/A _22656_/B _22700_/A _22656_/D vssd1 vssd1 vccd1 vccd1 _22710_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19324__A1 _19491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21607_ _21666_/A _21607_/B vssd1 vssd1 vccd1 vccd1 _21612_/C sky130_fd_sc_hd__and2_1
XANTENNA__16138__A1 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22587_ _22362_/B _22486_/Y _22489_/C _22663_/B _22586_/Y vssd1 vssd1 vccd1 vccd1
+ _22587_/Y sky130_fd_sc_hd__o2111ai_2
XFILLER_194_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17886__A1 _18016_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ _12339_/A _12339_/B _12339_/C vssd1 vssd1 vccd1 vccd1 _12340_/X sky130_fd_sc_hd__a21o_1
X_21538_ _21422_/B _21485_/A _21422_/A _21485_/B _21537_/Y vssd1 vssd1 vccd1 vccd1
+ _21540_/C sky130_fd_sc_hd__a41oi_4
XFILLER_139_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12271_ _12271_/A _12508_/D _19675_/C _12271_/D vssd1 vssd1 vccd1 vccd1 _12335_/D
+ sky130_fd_sc_hd__nand4_2
X_21469_ _21397_/A _21399_/B _21397_/B _21424_/A vssd1 vssd1 vccd1 vccd1 _21472_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_49_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _23357_/Q vssd1 vssd1 vccd1 vccd1 _14588_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23208_ _23254_/S vssd1 vssd1 vccd1 vccd1 _23217_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_88_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15649__B1 _16044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11922__A2 _11634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12902__D _12902_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23139_ _18997_/B input9/X _23145_/S vssd1 vssd1 vccd1 vccd1 _23140_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15961_ _11916_/X _16795_/C _17963_/C _12514_/B vssd1 vssd1 vccd1 vccd1 _16612_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_122_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_770 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14872__A1 _14097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17700_ _17700_/A _17700_/B vssd1 vssd1 vccd1 vccd1 _17832_/B sky130_fd_sc_hd__nand2_1
X_14912_ _13994_/A _13994_/B _15084_/A vssd1 vssd1 vccd1 vccd1 _14912_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13583__A _21891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18680_ _12184_/X _12185_/X _18678_/Y _19664_/B _18677_/Y vssd1 vssd1 vccd1 vccd1
+ _18681_/C sky130_fd_sc_hd__o2111ai_1
X_15892_ _15889_/X _15890_/Y _15867_/Y _15891_/Y vssd1 vssd1 vccd1 vccd1 _15892_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__12883__B1 _13151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_70 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22896__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17631_ _17631_/A vssd1 vssd1 vccd1 vccd1 _17960_/B sky130_fd_sc_hd__buf_2
X_14843_ _14844_/A _14844_/B _14844_/C vssd1 vssd1 vccd1 vccd1 _15065_/A sky130_fd_sc_hd__a21o_1
XFILLER_63_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_732 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17562_ _17562_/A _17562_/B vssd1 vssd1 vccd1 vccd1 _17562_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14774_ _14774_/A _14774_/B _14774_/C vssd1 vssd1 vccd1 vccd1 _14774_/Y sky130_fd_sc_hd__nand3_1
XFILLER_189_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11986_ _12105_/C vssd1 vssd1 vccd1 vccd1 _19000_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_523 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19301_ _19176_/Y _19179_/Y _19230_/B _19189_/X vssd1 vssd1 vccd1 vccd1 _19471_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16513_ _16483_/Y _16518_/C _16512_/Y vssd1 vssd1 vccd1 vccd1 _16522_/A sky130_fd_sc_hd__a21o_1
X_13725_ _13723_/Y _13727_/A _13727_/B vssd1 vssd1 vccd1 vccd1 _13730_/B sky130_fd_sc_hd__a21oi_1
X_17493_ _17493_/A _17493_/B _17493_/C vssd1 vssd1 vccd1 vccd1 _17497_/A sky130_fd_sc_hd__nand3_1
XFILLER_32_724 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12927__A _21050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11831__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19232_ _19232_/A _19240_/A _19240_/B vssd1 vssd1 vccd1 vccd1 _19256_/B sky130_fd_sc_hd__nand3_2
X_16444_ _16445_/A _16445_/B _16225_/X _16479_/A vssd1 vssd1 vccd1 vccd1 _16446_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1018 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13656_ _13680_/A _13656_/B vssd1 vssd1 vccd1 vccd1 _13674_/A sky130_fd_sc_hd__nand2_2
XANTENNA__19315__A1 _16437_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12938__A1 _12709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19163_ _19163_/A vssd1 vssd1 vccd1 vccd1 _19652_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12607_ _12683_/B vssd1 vssd1 vccd1 vccd1 _20495_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_157_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16129__A1 _11935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16375_ _16370_/X _16384_/A _17454_/B _16457_/D _16457_/A vssd1 vssd1 vccd1 vccd1
+ _16379_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_13_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21122__A1 _20773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _13698_/B _13587_/B vssd1 vssd1 vccd1 vccd1 _13587_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18114_ _18114_/A _18114_/B _18156_/A _18114_/D vssd1 vssd1 vccd1 vccd1 _18156_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_158_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ _15326_/A _15326_/B vssd1 vssd1 vccd1 vccd1 _15328_/A sky130_fd_sc_hd__nand2_1
X_19094_ _19094_/A _19094_/B vssd1 vssd1 vccd1 vccd1 _19106_/B sky130_fd_sc_hd__nand2_1
XFILLER_145_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12538_ _12531_/X _12533_/Y _12535_/Y _12537_/Y vssd1 vssd1 vccd1 vccd1 _12540_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_157_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15888__B1 _16423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18045_ _18045_/A _18045_/B vssd1 vssd1 vccd1 vccd1 _18129_/A sky130_fd_sc_hd__xor2_4
X_15257_ _15319_/C _15257_/B _15305_/A vssd1 vssd1 vccd1 vccd1 _15259_/B sky130_fd_sc_hd__and3_1
XFILLER_145_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12469_ _12469_/A _12469_/B _12469_/C vssd1 vssd1 vccd1 vccd1 _12478_/A sky130_fd_sc_hd__nand3_2
XANTENNA__19148__C _19148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17629__A1 _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14208_ _23360_/Q vssd1 vssd1 vccd1 vccd1 _15112_/C sky130_fd_sc_hd__clkinv_2
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14560__B1 _14693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15188_ _15188_/A _15188_/B _15188_/C _15188_/D vssd1 vssd1 vccd1 vccd1 _15190_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_bq_clk_i clkbuf_3_7_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _23578_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_98_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14139_ _14139_/A _14139_/B _14217_/C _14218_/A vssd1 vssd1 vccd1 vccd1 _14141_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19996_ _19996_/A _19996_/B _19996_/C vssd1 vssd1 vccd1 vccd1 _20003_/C sky130_fd_sc_hd__nand3_1
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16301__B2 _16055_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18947_ _18947_/A _18947_/B _18947_/C vssd1 vssd1 vccd1 vccd1 _18947_/X sky130_fd_sc_hd__and3_1
XANTENNA__19164__B _19652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18054__A1 _17943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22302__C _22392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18878_ _18889_/A _18889_/B _18867_/Y _19062_/A vssd1 vssd1 vccd1 vccd1 _18878_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20936__A1 _12709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_985 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17829_ _17820_/Y _17825_/Y _18148_/A vssd1 vssd1 vccd1 vccd1 _17831_/A sky130_fd_sc_hd__o21a_1
XANTENNA__22138__B1 _22139_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14101__B _14777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19180__A _19969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19003__B1 _19191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20840_ _20840_/A vssd1 vssd1 vccd1 vccd1 _20847_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21215__A _21215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20771_ _20688_/C _20680_/Y _20688_/B vssd1 vssd1 vccd1 vccd1 _20773_/B sky130_fd_sc_hd__o21ai_2
X_22510_ _22510_/A _22510_/B _22510_/C vssd1 vssd1 vccd1 vccd1 _22510_/X sky130_fd_sc_hd__and3_1
XFILLER_167_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23490_ _23510_/CLK _23502_/Q vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22441_ _22538_/A _22538_/B _22730_/B vssd1 vssd1 vccd1 vccd1 _22443_/A sky130_fd_sc_hd__a21o_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17317__B1 _17029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22372_ _22297_/B _22368_/Y _22365_/X _22362_/Y vssd1 vssd1 vccd1 vccd1 _22372_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21323_ _21317_/Y _21318_/X _21319_/Y vssd1 vssd1 vccd1 vccd1 _21327_/C sky130_fd_sc_hd__a21o_1
XFILLER_108_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16540__A1 _16558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12572__A _23301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16044__A _16044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21254_ _21246_/X _21247_/X _21345_/C vssd1 vssd1 vccd1 vccd1 _21254_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_190_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12291__B _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20205_ _20205_/A vssd1 vssd1 vccd1 vccd1 _20205_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15883__A _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19355__A _19391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19490__B1 _19847_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21185_ _21187_/A _21173_/X _21186_/A _21210_/B vssd1 vssd1 vccd1 vccd1 _21185_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20136_ _20151_/D _20151_/B _19803_/X _18328_/A vssd1 vssd1 vccd1 vccd1 _20136_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_89_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20067_ _20067_/A _20067_/B vssd1 vssd1 vccd1 vccd1 _20071_/A sky130_fd_sc_hd__nor2_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22129__B1 _22264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14606__A1 _23581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14606__B2 _14883_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17603__A _17761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11840_ _12432_/A vssd1 vssd1 vccd1 vccd1 _11840_/X sky130_fd_sc_hd__buf_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11771_ _23387_/Q vssd1 vssd1 vccd1 vccd1 _12245_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ _20969_/A vssd1 vssd1 vccd1 vccd1 _21356_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12747__A _23447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ _13400_/Y _13482_/A _22388_/B _13440_/Y _13650_/A vssd1 vssd1 vccd1 vccd1
+ _13555_/B sky130_fd_sc_hd__o2111ai_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22708_ _22754_/C _22754_/D vssd1 vssd1 vccd1 vccd1 _22800_/C sky130_fd_sc_hd__nor2_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14490_ _15082_/D vssd1 vssd1 vccd1 vccd1 _15446_/C sky130_fd_sc_hd__buf_2
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ _21793_/C _13810_/B _21793_/B vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__nand3_2
XANTENNA__21104__A1 _12640_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22639_ _22644_/A _22461_/X _22703_/A _22646_/A _22638_/Y vssd1 vssd1 vccd1 vccd1
+ _22642_/B sky130_fd_sc_hd__o221ai_1
XANTENNA__17308__B1 _17307_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18434__A _18434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17006__A_N _23519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17859__A1 _16684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16160_ _16160_/A vssd1 vssd1 vccd1 vccd1 _16499_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ _23326_/Q vssd1 vssd1 vccd1 vccd1 _13783_/B sky130_fd_sc_hd__inv_2
XFILLER_142_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15111_ _15111_/A _15111_/B vssd1 vssd1 vccd1 vccd1 _15112_/A sky130_fd_sc_hd__nor2_1
XFILLER_154_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12323_ _12323_/A vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__buf_4
XFILLER_181_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16091_ _16469_/A _16071_/Y _16062_/Y _16063_/X vssd1 vssd1 vccd1 vccd1 _16091_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_182_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15042_ _15044_/C _15195_/B _15038_/Y _15041_/Y vssd1 vssd1 vccd1 vccd1 _15045_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_181_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12254_ _12254_/A vssd1 vssd1 vccd1 vccd1 _12393_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_181_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19850_ _19855_/A _19855_/B _19855_/C vssd1 vssd1 vccd1 vccd1 _19850_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_122_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19481__B1 _19846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12185_ _12185_/A vssd1 vssd1 vccd1 vccd1 _12185_/X sky130_fd_sc_hd__buf_2
XANTENNA__22080__A2 _21994_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15098__A1 _14181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18801_ _18796_/X _18790_/X _18792_/Y _19511_/A _15928_/C vssd1 vssd1 vccd1 vccd1
+ _18802_/C sky130_fd_sc_hd__o2111ai_1
XANTENNA__16834__A2 _16058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19781_ _19781_/A _19781_/B _23547_/Q vssd1 vssd1 vccd1 vccd1 _19923_/A sky130_fd_sc_hd__nand3_1
XFILLER_110_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16993_ _17365_/C _17026_/C _17026_/D _17369_/A _17025_/A vssd1 vssd1 vccd1 vccd1
+ _16994_/C sky130_fd_sc_hd__a311o_1
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18732_ _19090_/B _19091_/A _18910_/A _18909_/C vssd1 vssd1 vccd1 vccd1 _18732_/Y
+ sky130_fd_sc_hd__nand4_2
X_15944_ _15948_/A _16246_/B _15859_/A _15943_/Y vssd1 vssd1 vccd1 vccd1 _15944_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__14202__A _14911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12320__A2 _11801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15875_ _18755_/D vssd1 vssd1 vccd1 vccd1 _19700_/D sky130_fd_sc_hd__buf_2
X_18663_ _11814_/A _12053_/A _12187_/Y _18656_/Y _18959_/A vssd1 vssd1 vccd1 vccd1
+ _18669_/B sky130_fd_sc_hd__o221ai_4
XANTENNA__15017__B _15225_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17614_ _17958_/A _17285_/X _17605_/Y _17606_/X _17607_/X vssd1 vssd1 vccd1 vccd1
+ _17614_/X sky130_fd_sc_hd__o311a_1
XFILLER_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14826_ _14826_/A _14826_/B _14826_/C vssd1 vssd1 vccd1 vccd1 _14826_/X sky130_fd_sc_hd__and3_1
X_18594_ _18545_/Y _18548_/Y _18557_/B vssd1 vssd1 vccd1 vccd1 _18728_/B sky130_fd_sc_hd__o21ai_1
XFILLER_184_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19536__A1 _17591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21035__A _21358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17545_ _19675_/C vssd1 vssd1 vccd1 vccd1 _19862_/A sky130_fd_sc_hd__buf_2
X_14757_ _14178_/B _14458_/A _14178_/A _14128_/A _14876_/B vssd1 vssd1 vccd1 vccd1
+ _14757_/Y sky130_fd_sc_hd__a32oi_4
X_11969_ _11969_/A _11969_/B _12227_/A vssd1 vssd1 vccd1 vccd1 _12227_/B sky130_fd_sc_hd__nand3_1
X_13708_ _22145_/C vssd1 vssd1 vccd1 vccd1 _22192_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_60_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17476_ _17487_/A _17487_/B _17480_/A _17481_/D vssd1 vssd1 vccd1 vccd1 _17482_/A
+ sky130_fd_sc_hd__a22o_1
X_14688_ _14688_/A vssd1 vssd1 vccd1 vccd1 _14688_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__21894__A2 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19215_ _19176_/Y _19179_/Y _19189_/X _19230_/B vssd1 vssd1 vccd1 vccd1 _19215_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15968__A _15968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16427_ _16422_/B _16336_/X _16424_/Y _16425_/Y vssd1 vssd1 vccd1 vccd1 _16427_/X
+ sky130_fd_sc_hd__o211a_1
X_13639_ _13434_/B _13434_/A _13414_/B vssd1 vssd1 vccd1 vccd1 _13639_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_81_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19146_ _19146_/A _19410_/C vssd1 vssd1 vccd1 vccd1 _19147_/B sky130_fd_sc_hd__nand2_1
X_16358_ _12379_/X _16356_/X _15802_/A _16757_/B vssd1 vssd1 vccd1 vccd1 _16572_/B
+ sky130_fd_sc_hd__o31a_2
XANTENNA__15687__B _23429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16117__A4 _18219_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15309_ _15419_/B vssd1 vssd1 vccd1 vccd1 _15511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19077_ _18893_/A _18893_/B _18893_/C _18895_/X vssd1 vssd1 vccd1 vccd1 _19077_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_146_968 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16289_ _17226_/D vssd1 vssd1 vccd1 vccd1 _17243_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_118_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18028_ _18028_/A _18028_/B _18028_/C vssd1 vssd1 vccd1 vccd1 _18033_/B sky130_fd_sc_hd__nand3_1
XFILLER_160_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22016__D _22276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17078__A2 _16377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15089__A1 _14097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20082__A1 _18016_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19979_ _20062_/B vssd1 vssd1 vccd1 vccd1 _20212_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14836__A1 _14298_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15208__A _15208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14112__A _14858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22990_ _13603_/X input38/X _22990_/S vssd1 vssd1 vccd1 vccd1 _22991_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21941_ _21941_/A _21994_/A _21994_/B vssd1 vssd1 vccd1 vccd1 _21941_/Y sky130_fd_sc_hd__nand3_2
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21871__C _21987_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17423__A _17625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21872_ _21801_/A _21801_/C _21801_/B vssd1 vssd1 vccd1 vccd1 _22096_/C sky130_fd_sc_hd__a21boi_1
XFILLER_36_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20823_ _20676_/B _20821_/X _20955_/A vssd1 vssd1 vccd1 vccd1 _20823_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23542_ _23582_/CLK _23542_/D vssd1 vssd1 vccd1 vccd1 _23542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20754_ _20754_/A vssd1 vssd1 vccd1 vccd1 _20754_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11902__C _11902_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23087__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23473_ _23499_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 _23473_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20685_ _20672_/X _20520_/Y _20678_/Y _20679_/Y vssd1 vssd1 vccd1 vccd1 _20688_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22424_ _22428_/A _22428_/B vssd1 vssd1 vccd1 vccd1 _22425_/C sky130_fd_sc_hd__nand2_1
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18502__A2 _19040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13398__A _23472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22355_ _22355_/A _22355_/B vssd1 vssd1 vccd1 vccd1 _23564_/D sky130_fd_sc_hd__xor2_4
XFILLER_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_776 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21306_ _21306_/A vssd1 vssd1 vccd1 vccd1 _21386_/B sky130_fd_sc_hd__clkbuf_2
X_22286_ _22279_/A _22386_/A _22656_/B _22284_/Y _22716_/A vssd1 vssd1 vccd1 vccd1
+ _22289_/D sky130_fd_sc_hd__o2111ai_4
XFILLER_85_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21237_ _21402_/A _21354_/A vssd1 vssd1 vccd1 vccd1 _21237_/Y sky130_fd_sc_hd__nand2_1
XFILLER_137_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21168_ _21083_/Y _21087_/Y _21089_/Y vssd1 vssd1 vccd1 vccd1 _21215_/A sky130_fd_sc_hd__o21ai_2
XFILLER_132_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11646__A _23587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20119_ _20032_/A _20032_/B _20029_/Y _20117_/X _20118_/X vssd1 vssd1 vccd1 vccd1
+ _20119_/Y sky130_fd_sc_hd__o311ai_2
XANTENNA__15118__A _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ _13985_/X _13989_/Y _13971_/X vssd1 vssd1 vccd1 vccd1 _13991_/B sky130_fd_sc_hd__o21bai_1
X_21099_ _21096_/X _21097_/X _21092_/Y _21098_/Y vssd1 vssd1 vccd1 vccd1 _21109_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__19766__A1 _19380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ _12941_/A vssd1 vssd1 vccd1 vccd1 _13181_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15660_ _15660_/A vssd1 vssd1 vccd1 vccd1 _17233_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12872_ _12872_/A vssd1 vssd1 vccd1 vccd1 _20907_/A sky130_fd_sc_hd__buf_2
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14055__A2 _14911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14611_ _23425_/Q vssd1 vssd1 vccd1 vccd1 _15921_/C sky130_fd_sc_hd__buf_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11823_ _11823_/A _11823_/B _11983_/A _12282_/A vssd1 vssd1 vccd1 vccd1 _11841_/A
+ sky130_fd_sc_hd__nand4_4
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15591_ _23514_/Q _23515_/Q _15586_/A hold23/A vssd1 vssd1 vccd1 vccd1 _15592_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22893__B _22895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17330_ _17330_/A _17330_/B _17330_/C vssd1 vssd1 vccd1 vccd1 _17331_/B sky130_fd_sc_hd__and3_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _16510_/C _14516_/X _14528_/X _14541_/X vssd1 vssd1 vccd1 vccd1 _14542_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11754_/A vssd1 vssd1 vccd1 vccd1 _12432_/A sky130_fd_sc_hd__buf_2
XFILLER_198_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12471__D1 _12260_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12196__B _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _18607_/C vssd1 vssd1 vccd1 vccd1 _17586_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14108_/Y _14933_/A _14436_/A _14436_/C _14472_/Y vssd1 vssd1 vccd1 vccd1
+ _14473_/X sky130_fd_sc_hd__o2111a_1
XANTENNA__23078__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11685_ _23388_/Q vssd1 vssd1 vccd1 vccd1 _12282_/A sky130_fd_sc_hd__inv_2
XANTENNA__16752__B2 _16275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19000_ _19163_/A _19000_/B _19308_/C vssd1 vssd1 vccd1 vccd1 _19000_/Y sky130_fd_sc_hd__nand3_1
X_16212_ _16201_/X _16205_/Y _16206_/Y _16211_/Y vssd1 vssd1 vccd1 vccd1 _16233_/B
+ sky130_fd_sc_hd__o211ai_4
X_13424_ _22039_/C vssd1 vssd1 vccd1 vccd1 _13810_/B sky130_fd_sc_hd__clkbuf_4
X_17192_ _16924_/Y _17166_/B _16937_/Y _16942_/X vssd1 vssd1 vccd1 vccd1 _17192_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_167_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16143_ _12497_/A _16142_/B _11723_/A vssd1 vssd1 vccd1 vccd1 _16817_/A sky130_fd_sc_hd__o21bai_2
XFILLER_154_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13355_ _13355_/A vssd1 vssd1 vccd1 vccd1 _22186_/C sky130_fd_sc_hd__buf_2
XFILLER_182_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ _12306_/A vssd1 vssd1 vccd1 vccd1 _16526_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_182_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16074_ _12174_/X _12173_/X _16462_/D _12175_/X vssd1 vssd1 vccd1 vccd1 _16539_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_6_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13286_ _13471_/A _13269_/X _13516_/A _13285_/X vssd1 vssd1 vccd1 vccd1 _13287_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_142_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19902_ _19894_/Y _19899_/Y _19901_/X vssd1 vssd1 vccd1 vccd1 _19902_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15025_ _14912_/X _14911_/Y _14910_/X vssd1 vssd1 vccd1 vccd1 _15030_/C sky130_fd_sc_hd__a21boi_2
XANTENNA__17508__A _18211_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12237_ _12237_/A vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__buf_4
XFILLER_30_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23250__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16412__A _19494_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20064__A1 _12113_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18330__C _20368_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_716 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19833_ _19876_/C vssd1 vssd1 vccd1 vccd1 _19833_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12168_ _12168_/A vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19764_ _19764_/A vssd1 vssd1 vccd1 vccd1 _19764_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16976_ _16970_/Y _16972_/X _16969_/C vssd1 vssd1 vccd1 vccd1 _16979_/A sky130_fd_sc_hd__o21ai_1
XFILLER_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12099_ _19155_/B _18469_/B _18998_/C _12099_/D vssd1 vssd1 vccd1 vccd1 _12100_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_65_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18715_ _18715_/A _18715_/B _18904_/A vssd1 vssd1 vccd1 vccd1 _18715_/X sky130_fd_sc_hd__and3_1
Xinput6 wb_cyc_i vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
XFILLER_77_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15927_ _15927_/A vssd1 vssd1 vccd1 vccd1 _17753_/A sky130_fd_sc_hd__buf_4
X_19695_ _12243_/X _17846_/X _11670_/X _17565_/A vssd1 vssd1 vccd1 vccd1 _19698_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17243__A _19949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18646_ _19196_/B _18453_/X _18462_/B _18634_/A vssd1 vssd1 vccd1 vccd1 _18647_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15858_ _15858_/A _15858_/B vssd1 vssd1 vccd1 vccd1 _15859_/C sky130_fd_sc_hd__nand2_1
XANTENNA__19161__C _19163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_487 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14809_ _14814_/A _14814_/B _14814_/C vssd1 vssd1 vccd1 vccd1 _14809_/Y sky130_fd_sc_hd__a21oi_1
X_18577_ _18912_/B vssd1 vssd1 vccd1 vccd1 _19090_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15789_ _15651_/Y _15670_/X _15786_/Y vssd1 vssd1 vccd1 vccd1 _15796_/A sky130_fd_sc_hd__o21ai_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17528_ _17528_/A _17528_/B vssd1 vssd1 vccd1 vccd1 _17529_/B sky130_fd_sc_hd__and2_1
XANTENNA__11804__A1 _11799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23069__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15698__A _15698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17459_ _20049_/A _17605_/A _17605_/B vssd1 vssd1 vccd1 vccd1 _17460_/B sky130_fd_sc_hd__and3_1
XANTENNA__16743__A1 _16480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14754__B1 _14181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20470_ _20628_/B vssd1 vssd1 vccd1 vccd1 _21493_/B sky130_fd_sc_hd__buf_2
XFILLER_146_721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19129_ _18953_/X _18952_/Y _18938_/X vssd1 vssd1 vccd1 vccd1 _19129_/X sky130_fd_sc_hd__a21bo_1
XFILLER_69_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_968 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22140_ _22153_/A vssd1 vssd1 vccd1 vccd1 _22474_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22071_ _22211_/A _22211_/B _22036_/X _22044_/Y _22054_/A vssd1 vssd1 vccd1 vccd1
+ _22073_/B sky130_fd_sc_hd__o221ai_1
XFILLER_99_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21022_ _21353_/A _21019_/C _21020_/Y _21021_/X vssd1 vssd1 vccd1 vccd1 _21029_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19646__A1_N _16032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17137__B _17625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22973_ _13226_/X input18/X _22979_/S vssd1 vssd1 vccd1 vccd1 _22974_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14777__A _14777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21924_ _21924_/A vssd1 vssd1 vccd1 vccd1 _22510_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_76_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ _21842_/A _21858_/D _13870_/Y vssd1 vssd1 vccd1 vccd1 _21859_/A sky130_fd_sc_hd__a21o_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20806_ _12765_/A _12862_/A _12877_/Y _20814_/A _20973_/A vssd1 vssd1 vccd1 vccd1
+ _20809_/B sky130_fd_sc_hd__o221ai_1
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14993__B1 _15338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21786_ _21786_/A _21786_/B vssd1 vssd1 vccd1 vccd1 _21786_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23525_ _23578_/CLK _23525_/D vssd1 vssd1 vccd1 vccd1 _23525_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20737_ _20737_/A _20737_/B _20737_/C vssd1 vssd1 vccd1 vccd1 _20738_/A sky130_fd_sc_hd__nand3_1
XFILLER_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22218__B _22218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13548__A1 _13547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15401__A _15442_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14745__B1 _14738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23456_ _23571_/CLK hold21/X vssd1 vssd1 vccd1 vccd1 _23456_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_167_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20668_ _20699_/A _20699_/B vssd1 vssd1 vccd1 vccd1 _20668_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22407_ _22406_/Y _22313_/X _22323_/A vssd1 vssd1 vccd1 vccd1 _22417_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__18487__A1 _11670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15120__B _15120_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18487__B2 _19491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23387_ _23389_/CLK _23387_/D vssd1 vssd1 vccd1 vccd1 _23387_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_192_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20599_ _20585_/A _20598_/X _21008_/A _20593_/C vssd1 vssd1 vccd1 vccd1 _20614_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12463__C _18756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20294__B2 _20243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13140_ _12962_/C _13140_/B _13140_/C vssd1 vssd1 vccd1 vccd1 _13141_/A sky130_fd_sc_hd__nand3b_1
X_22338_ _22357_/A _22357_/B _22356_/A vssd1 vssd1 vccd1 vccd1 _22341_/B sky130_fd_sc_hd__a21o_1
XFILLER_164_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13071_ _13077_/A _13077_/B vssd1 vssd1 vccd1 vccd1 _13079_/B sky130_fd_sc_hd__nand2_2
XFILLER_152_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22269_ _22566_/A _22566_/B _22269_/C vssd1 vssd1 vccd1 vccd1 _22269_/Y sky130_fd_sc_hd__nand3_2
XFILLER_151_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_982 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12022_ _12022_/A vssd1 vssd1 vccd1 vccd1 _12022_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18644__D1 _17134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input49_A x[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19543__A _19543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16830_ _12222_/X _12223_/X _15972_/X vssd1 vssd1 vccd1 vccd1 _16830_/X sky130_fd_sc_hd__a21o_1
XFILLER_66_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21758__A1_N _13797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16761_ _16755_/Y _16435_/C _16774_/B _17010_/B vssd1 vssd1 vccd1 vccd1 _16761_/Y
+ sky130_fd_sc_hd__o211ai_2
X_13973_ _14191_/A _14191_/B _13966_/X vssd1 vssd1 vccd1 vccd1 _14797_/C sky130_fd_sc_hd__a21o_1
XFILLER_47_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18500_ _18500_/A vssd1 vssd1 vccd1 vccd1 _18500_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15712_ _15712_/A _16187_/B _15712_/C _15712_/D vssd1 vssd1 vccd1 vccd1 _15713_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12924_ _21035_/C vssd1 vssd1 vccd1 vccd1 _21050_/C sky130_fd_sc_hd__clkbuf_2
X_19480_ _19480_/A vssd1 vssd1 vccd1 vccd1 _19480_/X sky130_fd_sc_hd__clkbuf_2
X_16692_ _16054_/A _16055_/A _15610_/X _16684_/X _15660_/A vssd1 vssd1 vccd1 vccd1
+ _16900_/B sky130_fd_sc_hd__o221a_1
XFILLER_34_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12919__B _21268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18431_ _23538_/Q _18431_/B vssd1 vssd1 vccd1 vccd1 _18431_/X sky130_fd_sc_hd__xor2_1
XFILLER_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12855_ _12677_/X _12704_/X _21035_/C _12705_/X vssd1 vssd1 vccd1 vccd1 _12855_/Y
+ sky130_fd_sc_hd__o211ai_4
X_15643_ _15630_/Y _15631_/Y _15791_/A vssd1 vssd1 vccd1 vccd1 _15647_/A sky130_fd_sc_hd__o21a_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16973__A1 _16663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11806_ _11916_/A vssd1 vssd1 vccd1 vccd1 _11853_/A sky130_fd_sc_hd__clkbuf_4
X_18362_ _18362_/A _18362_/B vssd1 vssd1 vccd1 vccd1 _18362_/Y sky130_fd_sc_hd__nand2_1
X_15574_ _15574_/A vssd1 vssd1 vccd1 vccd1 _15586_/C sky130_fd_sc_hd__clkbuf_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12668_/X _20493_/D _12618_/A vssd1 vssd1 vccd1 vccd1 _12824_/A sky130_fd_sc_hd__a21o_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _17313_/A _17313_/B _17313_/C vssd1 vssd1 vccd1 vccd1 _17326_/C sky130_fd_sc_hd__nand3_2
XFILLER_109_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14525_ _22896_/D vssd1 vssd1 vccd1 vccd1 _14546_/A sky130_fd_sc_hd__clkbuf_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11764_/A vssd1 vssd1 vccd1 vccd1 _16360_/A sky130_fd_sc_hd__clkbuf_4
X_18293_ _18293_/A _18293_/B vssd1 vssd1 vccd1 vccd1 _18305_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17244_ _19957_/D _18093_/A _17096_/X _17243_/X vssd1 vssd1 vccd1 vccd1 _17397_/B
+ sky130_fd_sc_hd__a31o_1
X_14456_ _14819_/A _14456_/B _14456_/C _15175_/C vssd1 vssd1 vccd1 vccd1 _14461_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_70_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11668_ _19363_/A _19363_/B vssd1 vssd1 vccd1 vccd1 _11669_/A sky130_fd_sc_hd__nand2_1
X_13407_ _13349_/X _13365_/Y _13367_/Y _22145_/C vssd1 vssd1 vccd1 vccd1 _13407_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_190_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17175_ _17179_/B _17179_/C _17179_/A vssd1 vssd1 vccd1 vccd1 _17334_/B sky130_fd_sc_hd__a21o_1
XFILLER_127_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14387_ _14114_/X _13969_/Y _14385_/Y _14396_/B vssd1 vssd1 vccd1 vccd1 _14390_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11599_ _11610_/C vssd1 vssd1 vccd1 vccd1 _18947_/B sky130_fd_sc_hd__buf_2
XFILLER_143_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16126_ _16126_/A vssd1 vssd1 vccd1 vccd1 _17712_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13338_ _13377_/B vssd1 vssd1 vccd1 vccd1 _13338_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13766__A _13766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16057_ _16054_/X _16055_/X _16056_/X _16028_/A _16028_/B vssd1 vssd1 vccd1 vccd1
+ _16060_/B sky130_fd_sc_hd__o2111ai_2
X_13269_ _13269_/A vssd1 vssd1 vccd1 vccd1 _13269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15700__A2 _16315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15008_ _14967_/X _14968_/X _15006_/Y _15007_/X vssd1 vssd1 vccd1 vccd1 _15035_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_155_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22982__A0 _13304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19816_ _19975_/B _19809_/X _19810_/Y _19815_/Y vssd1 vssd1 vccd1 vccd1 _19823_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_111_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16796__B _23597_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19747_ _19747_/A vssd1 vssd1 vccd1 vccd1 _19747_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19172__B _19172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16959_ _16944_/X _16949_/Y _17184_/A vssd1 vssd1 vccd1 vccd1 _16961_/A sky130_fd_sc_hd__a21o_1
XFILLER_110_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19678_ _19673_/Y _19676_/X _19682_/C vssd1 vssd1 vccd1 vccd1 _19678_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16413__B1 _17723_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18953__A2 _11834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18629_ _12130_/A _18490_/A _18446_/A _18443_/A vssd1 vssd1 vccd1 vccd1 _18804_/B
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__19900__B _20369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18219__D _18219_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21640_ _21668_/A _21641_/B _21635_/C _21502_/D _21641_/C vssd1 vssd1 vccd1 vccd1
+ _21642_/A sky130_fd_sc_hd__a41o_1
XFILLER_36_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21571_ _21577_/A _21611_/A _21568_/A _21568_/B vssd1 vssd1 vccd1 vccd1 _21614_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__17420__B _17420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23310_ _23345_/CLK _23310_/D vssd1 vssd1 vccd1 vccd1 _23310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20522_ _20501_/X _20520_/Y _20521_/Y _20518_/X _20492_/B vssd1 vssd1 vccd1 vccd1
+ _20523_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23241_ _23241_/A vssd1 vssd1 vccd1 vccd1 _23250_/S sky130_fd_sc_hd__clkbuf_2
X_20453_ _20453_/A _20453_/B vssd1 vssd1 vccd1 vccd1 _20453_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22265__A2 _22263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18532__A _19543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23172_ _23408_/Q input25/X _23178_/S vssd1 vssd1 vccd1 vccd1 _23173_/A sky130_fd_sc_hd__mux2_1
X_20384_ _20384_/A _20384_/B _20384_/C vssd1 vssd1 vccd1 vccd1 _20415_/B sky130_fd_sc_hd__nand3_1
XANTENNA__17141__A1 _16908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22123_ _22510_/A _22363_/A _22361_/C _22510_/C vssd1 vssd1 vccd1 vccd1 _22123_/Y
+ sky130_fd_sc_hd__nand4_2
XANTENNA__15152__B1 _13960_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22054_ _22054_/A vssd1 vssd1 vccd1 vccd1 _22197_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__22422__C1 _13431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22973__A0 _13226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21005_ _21157_/B _21157_/C vssd1 vssd1 vccd1 vccd1 _21005_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19363__A _19363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18641__A1 _12311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19082__B _19082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19197__A2 _11926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22220__C _22220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22956_ _23312_/Q input25/X _22962_/S vssd1 vssd1 vccd1 vccd1 _22957_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21907_ _22045_/A _22040_/A _21913_/B _22043_/A vssd1 vssd1 vccd1 vccd1 _21911_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_43_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_919 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22887_ _23446_/Q _22887_/B _22887_/C vssd1 vssd1 vccd1 vccd1 _22895_/A sky130_fd_sc_hd__and3b_4
XFILLER_102_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12640_ _12640_/A vssd1 vssd1 vccd1 vccd1 _12640_/X sky130_fd_sc_hd__buf_2
XFILLER_188_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21838_ _21836_/Y _21837_/Y _21834_/Y _21826_/X vssd1 vssd1 vccd1 vccd1 _21838_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20675__C _23453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12571_ _12571_/A vssd1 vssd1 vccd1 vccd1 _12571_/X sky130_fd_sc_hd__clkbuf_4
X_21769_ _13465_/X _22126_/A _13814_/Y _21783_/A _21984_/A vssd1 vssd1 vccd1 vccd1
+ _21769_/X sky130_fd_sc_hd__o311a_1
XFILLER_157_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_985 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14310_ _14310_/A _14310_/B _14310_/C _14310_/D vssd1 vssd1 vccd1 vccd1 _14310_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_184_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23508_ _23510_/CLK input44/X vssd1 vssd1 vccd1 vccd1 _23508_/Q sky130_fd_sc_hd__dfxtp_1
X_15290_ _15402_/A _14749_/X _15402_/B vssd1 vssd1 vccd1 vccd1 _15291_/B sky130_fd_sc_hd__a21oi_1
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15915__C1 _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ _15356_/A vssd1 vssd1 vccd1 vccd1 _15415_/A sky130_fd_sc_hd__buf_2
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23439_ _23441_/CLK _23439_/D vssd1 vssd1 vccd1 vccd1 _23439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20267__A1 _20055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14172_ _14172_/A _14172_/B _14429_/A vssd1 vssd1 vccd1 vccd1 _14756_/A sky130_fd_sc_hd__nand3_4
XFILLER_124_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17132__A1 _16480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17132__B2 _12311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13123_ _13133_/D _13124_/B _13124_/C vssd1 vssd1 vccd1 vccd1 _13125_/A sky130_fd_sc_hd__a21oi_1
XFILLER_125_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18980_ _18980_/A vssd1 vssd1 vccd1 vccd1 _20080_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15694__A1 _15674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17931_ _17928_/Y _17929_/X _17930_/Y vssd1 vssd1 vccd1 vccd1 _17932_/B sky130_fd_sc_hd__a21o_1
XFILLER_140_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13054_ _20961_/A _12766_/A _13053_/X vssd1 vssd1 vccd1 vccd1 _13054_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_121_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12005_ _11649_/X _16619_/A _11711_/C vssd1 vssd1 vccd1 vccd1 _16033_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__18632__A1 _11864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17862_ _20142_/D _17959_/A _17959_/B vssd1 vssd1 vccd1 vccd1 _17863_/B sky130_fd_sc_hd__and3_1
XANTENNA_repeater103_A _23481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater109 _23295_/CLK vssd1 vssd1 vccd1 vccd1 _23296_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18632__B2 _18440_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19601_ _19601_/A _19601_/B _19755_/A vssd1 vssd1 vccd1 vccd1 _19601_/X sky130_fd_sc_hd__and3_1
X_16813_ _16627_/X _17039_/A _16811_/X _16814_/A vssd1 vssd1 vccd1 vccd1 _17073_/B
+ sky130_fd_sc_hd__o211a_1
X_17793_ _17798_/A _17798_/C vssd1 vssd1 vccd1 vccd1 _17919_/B sky130_fd_sc_hd__nand2_1
XFILLER_120_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13457__B1 _22269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19532_ _19534_/A vssd1 vssd1 vccd1 vccd1 _19532_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11834__A _11834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16744_ _16744_/A _16744_/B _16784_/A vssd1 vssd1 vccd1 vccd1 _16744_/Y sky130_fd_sc_hd__nand3_2
X_13956_ _14796_/B vssd1 vssd1 vccd1 vccd1 _14911_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19463_ _19447_/A _19447_/B _19295_/A vssd1 vssd1 vccd1 vccd1 _19916_/A sky130_fd_sc_hd__a21oi_2
X_12907_ _12903_/Y _12904_/X _12905_/Y _12906_/Y vssd1 vssd1 vccd1 vccd1 _12908_/C
+ sky130_fd_sc_hd__o22ai_2
XFILLER_59_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16946__A1 _16934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13887_ _14863_/D _13939_/A _14863_/C vssd1 vssd1 vccd1 vccd1 _13890_/A sky130_fd_sc_hd__nand3b_2
X_16675_ _16675_/A vssd1 vssd1 vccd1 vccd1 _16911_/A sky130_fd_sc_hd__buf_2
XFILLER_185_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20742__A2 _20726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18414_ _18411_/X _18414_/B _18414_/C vssd1 vssd1 vccd1 vccd1 _18417_/B sky130_fd_sc_hd__nand3b_1
XFILLER_59_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12838_ _12904_/A vssd1 vssd1 vccd1 vccd1 _12991_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15626_ _15644_/A _15645_/A _15664_/C vssd1 vssd1 vccd1 vccd1 _15652_/A sky130_fd_sc_hd__a21o_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ _19401_/A _19398_/B _19390_/X _19393_/Y vssd1 vssd1 vccd1 vccd1 _19399_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_50_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23141__A0 _18799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18345_ _18345_/A _18388_/A _18346_/A vssd1 vssd1 vccd1 vccd1 _18348_/A sky130_fd_sc_hd__and3_1
XFILLER_159_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15557_ _15558_/A _15558_/C _15558_/B vssd1 vssd1 vccd1 vccd1 _15559_/A sky130_fd_sc_hd__o21a_2
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _23452_/Q vssd1 vssd1 vccd1 vccd1 _21054_/B sky130_fd_sc_hd__buf_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_624 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14508_ _16462_/D vssd1 vssd1 vccd1 vccd1 _16167_/C sky130_fd_sc_hd__clkbuf_2
X_18276_ _20265_/A _18328_/A _18276_/C _18330_/A vssd1 vssd1 vccd1 vccd1 _18277_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_148_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15488_ _15488_/A _15488_/B _15488_/C _15536_/B vssd1 vssd1 vccd1 vccd1 _15488_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__15906__C1 _16866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17227_ _16604_/X _17409_/A _17093_/Y vssd1 vssd1 vccd1 vccd1 _17236_/C sky130_fd_sc_hd__o21ai_2
Xinput20 wb_dat_i[21] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
X_14439_ _14443_/B _14442_/B _14439_/C vssd1 vssd1 vccd1 vccd1 _14441_/B sky130_fd_sc_hd__nand3_1
Xinput31 wb_dat_i[31] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 x[10] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_8
XFILLER_174_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19112__A2 _17581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12735__A2 _12722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17158_ _17220_/A _17220_/B _17220_/C vssd1 vssd1 vccd1 vccd1 _17179_/B sky130_fd_sc_hd__nand3_1
XFILLER_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_724 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11943__B1 _11942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16109_ _16549_/D vssd1 vssd1 vccd1 vccd1 _17326_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_171_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17089_ _17089_/A _17089_/B _17089_/C _17089_/D vssd1 vssd1 vccd1 vccd1 _17126_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__15220__D_N _15219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18623__A1 _18778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16229__A3 _17625_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18623__B2 _18615_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15988__A2 _15969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22810_ _22810_/A _22810_/B vssd1 vssd1 vccd1 vccd1 _22810_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13999__A1 _14331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21915__D1 _22364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17729__A3 _18017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22741_ _22738_/A _22738_/B _22740_/Y vssd1 vssd1 vccd1 vccd1 _22820_/A sky130_fd_sc_hd__a21oi_1
XFILLER_26_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17431__A _17431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22672_ _22676_/B _22720_/B vssd1 vssd1 vccd1 vccd1 _22675_/A sky130_fd_sc_hd__nand2_1
XFILLER_179_930 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23132__A0 _12121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20495__C _20495_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21623_ _21621_/Y _21622_/Y _21615_/X _21619_/Y vssd1 vssd1 vccd1 vccd1 _21624_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20497__A1 _20495_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21554_ _21595_/C _21554_/B _21554_/C _21554_/D vssd1 vssd1 vccd1 vccd1 _21555_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_193_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16285__B1_N _16856_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20505_ _20502_/X _20504_/X _20496_/X vssd1 vssd1 vccd1 vccd1 _21169_/A sky130_fd_sc_hd__o21a_1
XFILLER_193_454 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22238__A2 _22096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21485_ _21485_/A _21485_/B vssd1 vssd1 vccd1 vccd1 _21487_/A sky130_fd_sc_hd__nand2_1
XFILLER_181_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13384__C1 _13379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23224_ _23431_/Q input15/X _23228_/S vssd1 vssd1 vccd1 vccd1 _23225_/A sky130_fd_sc_hd__mux2_1
X_20436_ _20446_/B _20446_/C vssd1 vssd1 vccd1 vccd1 _20452_/A sky130_fd_sc_hd__nand2_1
XFILLER_134_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_830 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23155_ _23155_/A vssd1 vssd1 vccd1 vccd1 _23400_/D sky130_fd_sc_hd__clkbuf_1
X_20367_ _18376_/C _20265_/B _20318_/X _20366_/X vssd1 vssd1 vccd1 vccd1 _20379_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_122_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22106_ _22117_/D _22106_/B _22439_/D _22118_/B vssd1 vssd1 vccd1 vccd1 _22348_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__11638__B _16591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23086_ _23097_/A vssd1 vssd1 vccd1 vccd1 _23095_/S sky130_fd_sc_hd__clkbuf_2
X_20298_ _20298_/A vssd1 vssd1 vccd1 vccd1 _20343_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18614__A1 _12374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22037_ _22037_/A vssd1 vssd1 vccd1 vccd1 _22037_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_974 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11654__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ _22014_/A _13810_/B _21927_/A _22159_/C vssd1 vssd1 vccd1 vccd1 _13810_/Y
+ sky130_fd_sc_hd__nand4_2
X_14790_ _14796_/A _14790_/B _14790_/C vssd1 vssd1 vccd1 vccd1 _14798_/B sky130_fd_sc_hd__nand3_1
XANTENNA__14030__A _23498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__B1 _12104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13741_ _22474_/A _13741_/B _13741_/C vssd1 vssd1 vccd1 vccd1 _13741_/X sky130_fd_sc_hd__and3_1
X_22939_ _22939_/A vssd1 vssd1 vccd1 vccd1 _23304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16460_ _16404_/A _16405_/A _16457_/X _16459_/X vssd1 vssd1 vccd1 vccd1 _16467_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_13672_ _13680_/A _13680_/B _13672_/C vssd1 vssd1 vccd1 vccd1 _13672_/X sky130_fd_sc_hd__and3_1
XFILLER_189_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23123__A0 _11784_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_76 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15411_ _15366_/Y _15379_/A _15508_/A _15363_/A vssd1 vssd1 vccd1 vccd1 _15412_/B
+ sky130_fd_sc_hd__o211a_1
X_12623_ _20799_/A _13019_/C _13019_/B vssd1 vssd1 vccd1 vccd1 _12687_/B sky130_fd_sc_hd__o21bai_1
X_16391_ _16395_/A _16395_/B _16395_/C vssd1 vssd1 vccd1 vccd1 _16391_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12414__A1 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22477__A2 _22059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18130_ _18045_/B _18132_/C _18129_/Y _17957_/Y vssd1 vssd1 vccd1 vccd1 _18155_/A
+ sky130_fd_sc_hd__o22ai_4
X_15342_ _15528_/A vssd1 vssd1 vccd1 vccd1 _15478_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17889__C1 _17406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ _12537_/B _12537_/A _12531_/X _12533_/Y vssd1 vssd1 vccd1 vccd1 _12554_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_157_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18550__B1 _18526_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18061_ _18054_/Y _18057_/Y _23530_/Q _18060_/Y vssd1 vssd1 vccd1 vccd1 _18149_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_157_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15273_ _15190_/A _15193_/B _15271_/Y vssd1 vssd1 vccd1 vccd1 _15294_/A sky130_fd_sc_hd__a21o_1
XFILLER_145_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ _12480_/A _12480_/B _12483_/Y _12484_/Y _12490_/A vssd1 vssd1 vccd1 vccd1
+ _12487_/B sky130_fd_sc_hd__o221ai_1
XFILLER_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18172__A _18172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17012_ _17012_/A _17012_/B _17012_/C vssd1 vssd1 vccd1 vccd1 _17012_/Y sky130_fd_sc_hd__nand3_1
X_14224_ _14224_/A _14224_/B _14224_/C vssd1 vssd1 vccd1 vccd1 _14816_/A sky130_fd_sc_hd__nand3_2
XFILLER_184_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18838__D1 _19180_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14155_ _14152_/X _14005_/B _14154_/Y vssd1 vssd1 vccd1 vccd1 _14156_/C sky130_fd_sc_hd__o21a_1
XFILLER_180_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15667__A1 _15920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13106_ _13106_/A _13106_/B vssd1 vssd1 vccd1 vccd1 _13147_/B sky130_fd_sc_hd__nand2_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18963_ _18954_/Y _18955_/Y _18950_/Y _19410_/A vssd1 vssd1 vccd1 vccd1 _19410_/B
+ sky130_fd_sc_hd__o211ai_2
X_14086_ _14086_/A _14086_/B _14094_/A vssd1 vssd1 vccd1 vccd1 _14203_/A sky130_fd_sc_hd__nand3_2
XFILLER_152_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _17915_/A _17912_/X _17913_/Y vssd1 vssd1 vccd1 vccd1 _17919_/C sky130_fd_sc_hd__o21ai_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _12862_/A _12851_/Y _13029_/B _13029_/A vssd1 vssd1 vccd1 vccd1 _13037_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_79_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18894_ _18619_/A _18619_/B _18619_/C _18715_/A vssd1 vssd1 vccd1 vccd1 _18904_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_26_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14859__B _14980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17845_ _19534_/B _19799_/C _17845_/C _17845_/D vssd1 vssd1 vccd1 vccd1 _17855_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16092__A1 _16089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20963__A2 _12722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17776_ _17616_/B _17616_/C _17616_/A vssd1 vssd1 vccd1 vccd1 _17776_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_82_828 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22165__A1 _22474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14988_ _14976_/A _15422_/A _14985_/X _14987_/Y vssd1 vssd1 vccd1 vccd1 _15124_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_75_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19515_ _19525_/C _19525_/D vssd1 vssd1 vccd1 vccd1 _19524_/B sky130_fd_sc_hd__nand2_2
X_16727_ _16721_/Y _16724_/X _16735_/C vssd1 vssd1 vccd1 vccd1 _16732_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__16919__A1 _15932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13939_ _13939_/A vssd1 vssd1 vccd1 vccd1 _14091_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17577__D1 _17845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19446_ _19625_/B vssd1 vssd1 vccd1 vccd1 _19447_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_50_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16658_ _23426_/Q _16658_/B _16658_/C vssd1 vssd1 vccd1 vccd1 _16665_/A sky130_fd_sc_hd__nor3_4
XFILLER_23_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15609_ _15715_/A _16658_/B vssd1 vssd1 vccd1 vccd1 _16683_/A sky130_fd_sc_hd__nor2_1
X_19377_ _19219_/X _19220_/Y _19205_/X _19202_/Y vssd1 vssd1 vccd1 vccd1 _19385_/B
+ sky130_fd_sc_hd__o22ai_2
X_16589_ _16598_/A _16598_/B _16588_/X vssd1 vssd1 vccd1 vccd1 _16590_/B sky130_fd_sc_hd__o21ai_2
XFILLER_15_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19333__A2 _19803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18328_ _18328_/A vssd1 vssd1 vccd1 vccd1 _18373_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18259_ _18364_/B _23533_/Q _18364_/A vssd1 vssd1 vccd1 vccd1 _18319_/B sky130_fd_sc_hd__nand3_1
XFILLER_148_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18082__A _20215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16552__C1 _16510_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21858__D _21858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21270_ _21270_/A _21270_/B _21270_/C vssd1 vssd1 vccd1 vccd1 _21274_/C sky130_fd_sc_hd__nand3_1
XFILLER_144_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16314__B _16314_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20221_ _20222_/A _20277_/B _20219_/X _20220_/Y vssd1 vssd1 vccd1 vccd1 _20221_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__22035__C _22035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17647__A2 _18276_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20651__A1 _12675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20152_ _19539_/A _20151_/C _19539_/B _20151_/B _20134_/A vssd1 vssd1 vccd1 vccd1
+ _20158_/D sky130_fd_sc_hd__a32o_1
XFILLER_171_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20083_ _20083_/A _20083_/B vssd1 vssd1 vccd1 vccd1 _20083_/Y sky130_fd_sc_hd__nand2_2
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19006__D1 _19180_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22156__A1 _13732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12289__B _12289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19021__B2 _11961_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20985_ _21111_/B _20987_/B _21111_/A vssd1 vssd1 vccd1 vccd1 _20985_/X sky130_fd_sc_hd__and3_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17161__A _17161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22724_ _22586_/Y _22657_/Y _22664_/X _22484_/X _22237_/X vssd1 vssd1 vccd1 vccd1
+ _22725_/B sky130_fd_sc_hd__a311o_1
XFILLER_81_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11921__B _23256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22655_ _22577_/Y _22573_/Y _22713_/D _22712_/A vssd1 vssd1 vccd1 vccd1 _22656_/D
+ sky130_fd_sc_hd__o211ai_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21606_ _21645_/B _21605_/B _21605_/C vssd1 vssd1 vccd1 vccd1 _21607_/B sky130_fd_sc_hd__o21ai_1
XFILLER_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16138__A2 _16056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22586_ _22469_/X _22567_/Y _22468_/X _22579_/Y _22650_/B vssd1 vssd1 vccd1 vccd1
+ _22586_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_21_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21537_ _21535_/X _21485_/B _21536_/Y vssd1 vssd1 vccd1 vccd1 _21537_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_194_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17886__A2 _20164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12270_ _12508_/D _19675_/C _12271_/A _12271_/D vssd1 vssd1 vccd1 vccd1 _12335_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21468_ _21468_/A _21468_/B vssd1 vssd1 vccd1 vccd1 _21472_/B sky130_fd_sc_hd__xor2_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17099__B1 _11935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23207_ _23207_/A vssd1 vssd1 vccd1 vccd1 _23423_/D sky130_fd_sc_hd__clkbuf_1
X_20419_ _23556_/Q _20419_/B vssd1 vssd1 vccd1 vccd1 _20419_/X sky130_fd_sc_hd__or2_1
XFILLER_88_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21399_ _21424_/A _21399_/B _21399_/C vssd1 vssd1 vccd1 vccd1 _21400_/B sky130_fd_sc_hd__nand3b_1
XFILLER_134_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23138_ _23138_/A vssd1 vssd1 vccd1 vccd1 _23392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15960_ _16141_/D vssd1 vssd1 vccd1 vccd1 _17963_/C sky130_fd_sc_hd__buf_2
X_23069_ _14621_/X input10/X _23073_/S vssd1 vssd1 vccd1 vccd1 _23070_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input31_A wb_dat_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ _14911_/A _14911_/B _14911_/C _15075_/A vssd1 vssd1 vccd1 vccd1 _14911_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_49_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15891_ _15985_/C _15866_/B _15879_/Y vssd1 vssd1 vccd1 vccd1 _15891_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17630_ _17410_/Y _17625_/Y _17629_/Y vssd1 vssd1 vccd1 vccd1 _17634_/A sky130_fd_sc_hd__o21ai_1
XFILLER_124_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14842_ _14842_/A _14842_/B vssd1 vssd1 vccd1 vccd1 _14844_/C sky130_fd_sc_hd__nand2_1
XFILLER_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17561_ _17475_/A _17475_/B _17475_/C _17481_/C _17487_/Y vssd1 vssd1 vccd1 vccd1
+ _17653_/A sky130_fd_sc_hd__a32oi_1
XFILLER_17_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14773_ _14990_/A _14990_/B _15116_/B vssd1 vssd1 vccd1 vccd1 _14773_/Y sky130_fd_sc_hd__nand3_2
X_11985_ _12426_/C vssd1 vssd1 vccd1 vccd1 _19019_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_17_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19300_ _19239_/X _19240_/Y _19226_/A _19242_/Y vssd1 vssd1 vccd1 vccd1 _19399_/A
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16512_ _16512_/A _16532_/C _16532_/B vssd1 vssd1 vccd1 vccd1 _16512_/Y sky130_fd_sc_hd__nand3_1
XFILLER_1_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13724_ _13723_/C _13723_/B _13717_/Y vssd1 vssd1 vccd1 vccd1 _13727_/B sky130_fd_sc_hd__a21boi_1
XFILLER_189_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17492_ _17386_/X _17387_/Y _17490_/Y _17491_/X vssd1 vssd1 vccd1 vccd1 _17502_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_189_546 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19231_ _19052_/B _19037_/A _19048_/Y _19046_/Y vssd1 vssd1 vccd1 vccd1 _19240_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__14388__A1 _13972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16443_ _17134_/B _16499_/A _16443_/C _19503_/C vssd1 vssd1 vccd1 vccd1 _16445_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14388__B2 _14876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13655_ _13655_/A vssd1 vssd1 vccd1 vccd1 _13671_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_176_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19315__A2 _19858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19162_ _19162_/A _19162_/B vssd1 vssd1 vccd1 vccd1 _19167_/B sky130_fd_sc_hd__nand2_1
X_12606_ _12606_/A _12606_/B _12606_/C vssd1 vssd1 vccd1 vccd1 _12606_/Y sky130_fd_sc_hd__nand3_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16129__A2 _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16374_ _16374_/A vssd1 vssd1 vccd1 vccd1 _16457_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13586_ _13686_/A _22700_/D _13756_/A _13756_/B vssd1 vssd1 vccd1 vccd1 _13587_/B
+ sky130_fd_sc_hd__a211oi_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21122__A2 _20773_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _18114_/A _18114_/B _18156_/A _18114_/D vssd1 vssd1 vccd1 vccd1 _18118_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_157_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12537_ _12537_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _12537_/Y sky130_fd_sc_hd__nand2_1
X_15325_ _15324_/A _15324_/B _15380_/A _15323_/X vssd1 vssd1 vccd1 vccd1 _15328_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_19093_ _19094_/A _19109_/A _19094_/B vssd1 vssd1 vccd1 vccd1 _19106_/A sky130_fd_sc_hd__a21o_1
XANTENNA__18480__A_N _18474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15888__A1 _15878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ _18132_/A _18132_/B vssd1 vssd1 vccd1 vccd1 _18045_/B sky130_fd_sc_hd__or2_2
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ _11766_/A _11926_/A _12177_/B _18675_/C _12461_/Y vssd1 vssd1 vccd1 vccd1
+ _12469_/C sky130_fd_sc_hd__o221ai_2
X_15256_ _15265_/A _15353_/A _15353_/B _15303_/A _15303_/D vssd1 vssd1 vccd1 vccd1
+ _15259_/A sky130_fd_sc_hd__a32o_1
XFILLER_32_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14207_ _14031_/X _14061_/X _14312_/C vssd1 vssd1 vccd1 vccd1 _14207_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__14560__A1 input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17629__A2 _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14560__B2 _11677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15187_ _15249_/A _15250_/A _15187_/C vssd1 vssd1 vccd1 vccd1 _15188_/D sky130_fd_sc_hd__nand3_1
XFILLER_153_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12399_ _12399_/A _12399_/B _12399_/C vssd1 vssd1 vccd1 vccd1 _12399_/X sky130_fd_sc_hd__and3_1
XFILLER_125_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_991 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14218_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19995_ _19992_/X _19835_/Y _19987_/Y _19991_/Y vssd1 vssd1 vccd1 vccd1 _19996_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_152_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17891__D _19957_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12459__B1_N _12110_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18946_ _11815_/A _17975_/A _12353_/A _17431_/A vssd1 vssd1 vccd1 vccd1 _19261_/A
+ sky130_fd_sc_hd__o22ai_4
X_14069_ _14069_/A vssd1 vssd1 vccd1 vccd1 _14069_/X sky130_fd_sc_hd__buf_2
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20397__B1 _20384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18877_ _18868_/X _18870_/Y _18875_/X _18884_/A vssd1 vssd1 vccd1 vccd1 _19062_/A
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__20936__A2 _21592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17828_ _17828_/A _17828_/B _23528_/Q vssd1 vssd1 vccd1 vccd1 _18148_/A sky130_fd_sc_hd__nand3_1
XFILLER_95_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17759_ _17759_/A _17759_/B _17759_/C vssd1 vssd1 vccd1 vccd1 _17773_/A sky130_fd_sc_hd__nand3_2
XANTENNA__19003__B2 _19210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20770_ _20669_/X _20670_/X _20683_/X _20769_/Y _20688_/A vssd1 vssd1 vccd1 vccd1
+ _20770_/X sky130_fd_sc_hd__o311a_1
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21361__A2 _20471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19429_ _19116_/C _19425_/X _19116_/A vssd1 vssd1 vccd1 vccd1 _19616_/B sky130_fd_sc_hd__o21ai_2
XFILLER_23_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22440_ _22342_/A _22438_/Y _22246_/B _22439_/Y vssd1 vssd1 vccd1 vccd1 _22730_/B
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__22846__C1 _22858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17317__A1 _16054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17317__B2 _16665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18524__B _18524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20773__C _20773_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22371_ _13527_/X _22479_/A _22279_/A _22386_/A vssd1 vssd1 vccd1 vccd1 _22371_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_191_700 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21322_ _21225_/X _21221_/B _21321_/Y vssd1 vssd1 vccd1 vccd1 _21322_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16540__A2 _16530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21253_ _21342_/B _21253_/B vssd1 vssd1 vccd1 vccd1 _21345_/C sky130_fd_sc_hd__nand2_1
XFILLER_150_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20204_ _23552_/Q vssd1 vssd1 vccd1 vccd1 _20255_/A sky130_fd_sc_hd__inv_2
XFILLER_144_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23158__A _23169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21184_ _21184_/A _21184_/B _21184_/C _21184_/D vssd1 vssd1 vccd1 vccd1 _21210_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_145_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13684__A _23480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20135_ _20151_/A _20151_/B _20212_/D _20151_/D vssd1 vssd1 vccd1 vccd1 _20135_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_132_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16698__C _16706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20066_ _20066_/A _20066_/B _20066_/C vssd1 vssd1 vccd1 vccd1 _20067_/B sky130_fd_sc_hd__and3_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17253__B1 _16370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23552__CLK _23558_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15803__A1 _17465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17005__B1 _23520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11823_/A _11823_/B _11999_/A vssd1 vssd1 vccd1 vccd1 _11861_/A sky130_fd_sc_hd__nand3_4
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ _20973_/A _20973_/B _21101_/B _21101_/C vssd1 vssd1 vccd1 vccd1 _20975_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_54_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22707_ _22707_/A _22707_/B vssd1 vssd1 vccd1 vccd1 _22754_/D sky130_fd_sc_hd__nand2_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17041__D _20317_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20899_ _21174_/A _20905_/C _21174_/C vssd1 vssd1 vccd1 vccd1 _20899_/Y sky130_fd_sc_hd__nand3_1
XFILLER_16_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ _13440_/A _13440_/B vssd1 vssd1 vccd1 vccd1 _13440_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22638_ _13547_/X _22164_/A _22637_/Y vssd1 vssd1 vccd1 vccd1 _22638_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_186_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17308__A1 _17140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13042__A1 _13122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18505__B1 _18504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21104__A2 _12637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22301__A1 _22644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18434__B _18434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13371_ _13354_/Y _22186_/C _13802_/B _13486_/A vssd1 vssd1 vccd1 vccd1 _13376_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_194_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17859__A2 _16683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22569_ _22569_/A _22569_/B _22569_/C vssd1 vssd1 vccd1 vccd1 _22577_/B sky130_fd_sc_hd__nand3_2
XFILLER_154_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12322_ _12360_/A _12360_/B _12381_/C _12381_/B vssd1 vssd1 vccd1 vccd1 _12336_/A
+ sky130_fd_sc_hd__a22o_1
X_15110_ _15253_/A vssd1 vssd1 vccd1 vccd1 _15110_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16090_ _16094_/A _16052_/X _16326_/A vssd1 vssd1 vccd1 vccd1 _16090_/X sky130_fd_sc_hd__o21a_1
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15041_ _15041_/A _15041_/B vssd1 vssd1 vccd1 vccd1 _15041_/Y sky130_fd_sc_hd__nor2_1
X_12253_ _12253_/A vssd1 vssd1 vccd1 vccd1 _12393_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__14542__A1 _16510_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12184_ _12184_/A vssd1 vssd1 vccd1 vccd1 _12184_/X sky130_fd_sc_hd__buf_2
XFILLER_107_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16295__A1 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18800_ _18800_/A _18800_/B vssd1 vssd1 vccd1 vccd1 _19511_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17066__A _19700_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19780_ _19783_/A _19793_/A _19916_/D vssd1 vssd1 vccd1 vccd1 _19781_/B sky130_fd_sc_hd__a21o_1
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16992_ _17011_/C vssd1 vssd1 vccd1 vccd1 _17376_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ _19091_/A _18910_/A _18909_/C _19090_/B vssd1 vssd1 vccd1 vccd1 _18731_/X
+ sky130_fd_sc_hd__a22o_1
X_15943_ _15943_/A _15943_/B vssd1 vssd1 vccd1 vccd1 _15943_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20918__A2 _14615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13744__D _21832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18662_ _18662_/A _18662_/B vssd1 vssd1 vccd1 vccd1 _18669_/A sky130_fd_sc_hd__nand2_2
XFILLER_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _18600_/B vssd1 vssd1 vccd1 vccd1 _18755_/D sky130_fd_sc_hd__buf_2
XFILLER_95_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15017__C _15253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21591__A2 _21432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17613_ _17613_/A vssd1 vssd1 vccd1 vccd1 _17958_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _14825_/A _14825_/B _14825_/C vssd1 vssd1 vccd1 vccd1 _14830_/A sky130_fd_sc_hd__nand3_1
XFILLER_92_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _18593_/A _18593_/B vssd1 vssd1 vccd1 vccd1 _23520_/D sky130_fd_sc_hd__nand2_1
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19536__A2 _17593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17544_ _17663_/A _17663_/B _17483_/A _17543_/X vssd1 vssd1 vccd1 vccd1 _17661_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_45_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _14756_/A _14756_/B vssd1 vssd1 vccd1 vccd1 _14756_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21035__B _21358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17547__A1 _17546_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ _11968_/A vssd1 vssd1 vccd1 vccd1 _12227_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_189_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17547__B2 _19862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13707_ _21778_/C _21987_/C _21987_/A _13736_/A _22192_/C vssd1 vssd1 vccd1 vccd1
+ _13707_/X sky130_fd_sc_hd__a32o_1
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17475_ _17475_/A _17475_/B _17475_/C vssd1 vssd1 vccd1 vccd1 _17481_/D sky130_fd_sc_hd__nand3_2
X_11899_ _11670_/X _11898_/X _11891_/A vssd1 vssd1 vccd1 vccd1 _11902_/B sky130_fd_sc_hd__o21ai_4
X_14687_ _23404_/Q _14672_/X _14677_/X _23436_/Q _14686_/X vssd1 vssd1 vccd1 vccd1
+ _14687_/X sky130_fd_sc_hd__a221o_1
XANTENNA__21894__A3 _21892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19214_ _19202_/Y _19206_/X _19213_/Y vssd1 vssd1 vccd1 vccd1 _19230_/B sky130_fd_sc_hd__o21ai_2
XFILLER_34_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16426_ _16421_/Y _16422_/Y _16424_/Y _16425_/Y vssd1 vssd1 vccd1 vccd1 _16426_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_13638_ _13645_/A _13645_/B _13633_/X _13637_/X vssd1 vssd1 vccd1 vccd1 _13646_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_160_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19145_ _19409_/A _19409_/B _19409_/C _19144_/X vssd1 vssd1 vccd1 vccd1 _19146_/A
+ sky130_fd_sc_hd__a31oi_2
X_16357_ _16356_/X _15800_/Y _18172_/D _14735_/A _16046_/Y vssd1 vssd1 vccd1 vccd1
+ _16757_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_146_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13569_ _13569_/A _13569_/B _13569_/C vssd1 vssd1 vccd1 vccd1 _13569_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__12673__A _23451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15308_ _15308_/A _15363_/D _15409_/A _15308_/D vssd1 vssd1 vccd1 vccd1 _15311_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_172_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19076_ _18617_/X _18928_/X _19087_/B vssd1 vssd1 vccd1 vccd1 _19076_/Y sky130_fd_sc_hd__o21ai_1
X_16288_ _17845_/C vssd1 vssd1 vccd1 vccd1 _17974_/D sky130_fd_sc_hd__clkbuf_4
X_18027_ _17902_/B _17881_/Y _17873_/Y _17868_/Y vssd1 vssd1 vccd1 vccd1 _18028_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_15239_ _15171_/Y _15238_/Y _15234_/Y vssd1 vssd1 vccd1 vccd1 _15239_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__15730__B1 _14553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18275__A2 _18211_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1043 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19978_ _19980_/C _19972_/A _19973_/X vssd1 vssd1 vccd1 vccd1 _20073_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__18680__C1 _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14836__A2 _15054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18929_ _18708_/B _18751_/X _18892_/A vssd1 vssd1 vccd1 vccd1 _18929_/X sky130_fd_sc_hd__o21a_1
XFILLER_140_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15208__B _15408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17704__A _18059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19191__A _19191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21940_ _21940_/A _21940_/B vssd1 vssd1 vccd1 vccd1 _21994_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13009__A _23296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21871_ _21987_/A _22220_/C _21987_/C vssd1 vssd1 vccd1 vccd1 _21873_/A sky130_fd_sc_hd__and3_1
XFILLER_83_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20822_ _12784_/A _12722_/A _20674_/Y vssd1 vssd1 vccd1 vccd1 _20955_/A sky130_fd_sc_hd__o21ai_1
XFILLER_78_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1052 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23541_ _23566_/CLK _23541_/D vssd1 vssd1 vccd1 vccd1 _23541_/Q sky130_fd_sc_hd__dfxtp_1
X_20753_ _20615_/Y _20616_/Y _20605_/B _21011_/A vssd1 vssd1 vccd1 vccd1 _20754_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1096 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23472_ _23499_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 _23472_/Q sky130_fd_sc_hd__dfxtp_4
X_20684_ _20669_/X _20670_/X _20680_/Y _20683_/X vssd1 vssd1 vccd1 vccd1 _20715_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22423_ _22237_/A _13431_/X _22419_/Y _22421_/X vssd1 vssd1 vccd1 vccd1 _22428_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_176_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16055__A _16055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22354_ _22354_/A _22452_/B vssd1 vssd1 vccd1 vccd1 _22355_/B sky130_fd_sc_hd__or2_2
XFILLER_136_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21305_ _21307_/A _21307_/B _21306_/A _21307_/D vssd1 vssd1 vccd1 vccd1 _21308_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22285_ _22479_/A vssd1 vssd1 vccd1 vccd1 _22716_/A sky130_fd_sc_hd__buf_2
XFILLER_191_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21236_ _21236_/A _21236_/B _21236_/C vssd1 vssd1 vccd1 vccd1 _21354_/A sky130_fd_sc_hd__nand3_1
XFILLER_137_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11927__A _16593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21167_ _21162_/Y _21165_/X _21166_/Y vssd1 vssd1 vccd1 vccd1 _21221_/A sky130_fd_sc_hd__o21ai_1
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20118_ _20306_/A vssd1 vssd1 vccd1 vccd1 _20118_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16682__D1 _17420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21098_ _21097_/X _21087_/Y _21083_/Y vssd1 vssd1 vccd1 vccd1 _21098_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_172_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20049_ _20049_/A _20215_/B _20215_/C vssd1 vssd1 vccd1 vccd1 _20049_/Y sky130_fd_sc_hd__nand3_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12940_ _20955_/C vssd1 vssd1 vccd1 vccd1 _21121_/A sky130_fd_sc_hd__buf_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15788__B1 _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _12871_/A vssd1 vssd1 vccd1 vccd1 _20906_/A sky130_fd_sc_hd__buf_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14055__A3 _14760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14610_ _23393_/Q vssd1 vssd1 vccd1 vccd1 _18997_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11822_/A vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14996__D1 _14469_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15590_ _23515_/Q _15590_/B vssd1 vssd1 vccd1 vccd1 _23503_/D sky130_fd_sc_hd__xnor2_1
XFILLER_45_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14460__B1 _14181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _21832_/A _14532_/X _14534_/X _14540_/X vssd1 vssd1 vccd1 vccd1 _14541_/X
+ sky130_fd_sc_hd__a211o_1
X_11753_ _11977_/B vssd1 vssd1 vccd1 vccd1 _11999_/A sky130_fd_sc_hd__inv_2
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16201__A1 _11822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16201__B2 _11848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17260_ _17260_/A _17260_/B vssd1 vssd1 vccd1 vccd1 _17260_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_886 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14472_ _14933_/A _14472_/B _14472_/C _14472_/D vssd1 vssd1 vccd1 vccd1 _14472_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _11684_/A vssd1 vssd1 vccd1 vccd1 _12282_/B sky130_fd_sc_hd__buf_2
XFILLER_187_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14212__B1 _14097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23448__CLK _23462_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16211_ _11766_/B _15655_/X _16217_/A vssd1 vssd1 vccd1 vccd1 _16211_/Y sky130_fd_sc_hd__o21ai_1
X_13423_ _13423_/A vssd1 vssd1 vccd1 vccd1 _22521_/A sky130_fd_sc_hd__clkbuf_2
X_17191_ _17184_/A _16944_/X _16949_/Y _16961_/C vssd1 vssd1 vccd1 vccd1 _17191_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16142_ _17964_/C _16142_/B vssd1 vssd1 vccd1 vccd1 _17742_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13354_ _13308_/Y _13354_/B _13354_/C _13783_/C vssd1 vssd1 vccd1 vccd1 _13354_/Y
+ sky130_fd_sc_hd__nand4b_1
XFILLER_139_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17162__C1 _17152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12305_ _12547_/A _12303_/Y _12547_/B vssd1 vssd1 vccd1 vccd1 _12305_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_127_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15459__C_N _15353_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13285_ _13465_/A _13257_/A _13284_/Y vssd1 vssd1 vccd1 vccd1 _13285_/X sky130_fd_sc_hd__o21a_1
X_16073_ _16073_/A _16073_/B vssd1 vssd1 vccd1 vccd1 _16073_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__23598__CLK _23598_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19901_ _19903_/C _19903_/B _19903_/A _19900_/X vssd1 vssd1 vccd1 vccd1 _19901_/X
+ sky130_fd_sc_hd__a31o_1
X_12236_ _16408_/A vssd1 vssd1 vccd1 vccd1 _12237_/A sky130_fd_sc_hd__buf_2
X_15024_ _15081_/B _15022_/C _15022_/A vssd1 vssd1 vccd1 vccd1 _15030_/B sky130_fd_sc_hd__a21o_1
XANTENNA__18257__A2 _18417_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20215__A _20215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19832_ _19723_/C _19831_/X _19723_/B vssd1 vssd1 vccd1 vccd1 _19876_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__18330__D _18376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ _12167_/A vssd1 vssd1 vccd1 vccd1 _12167_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19763_ _19380_/X _19621_/X _19620_/X vssd1 vssd1 vccd1 vccd1 _19763_/X sky130_fd_sc_hd__o21a_1
XANTENNA__19206__A1 _19013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16975_ _16975_/A _16975_/B vssd1 vssd1 vccd1 vccd1 _16975_/Y sky130_fd_sc_hd__nand2_1
X_12098_ _18649_/A vssd1 vssd1 vccd1 vccd1 _19155_/B sky130_fd_sc_hd__buf_2
X_18714_ _18715_/B _18904_/A _18715_/A vssd1 vssd1 vccd1 vccd1 _18714_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15926_ _12052_/A _17409_/A _15917_/Y _15923_/X _15925_/Y vssd1 vssd1 vccd1 vccd1
+ _15926_/X sky130_fd_sc_hd__o311a_2
X_19694_ _19694_/A _19799_/C _19967_/A _19900_/D vssd1 vssd1 vccd1 vccd1 _19698_/C
+ sky130_fd_sc_hd__nand4_2
Xinput7 wb_dat_i[0] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_6
XFILLER_37_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22761__A1 _21997_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18645_ _18645_/A vssd1 vssd1 vccd1 vccd1 _19196_/B sky130_fd_sc_hd__buf_2
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17243__B _17243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15857_ _12174_/X _12173_/X _15855_/Y _15856_/Y _12175_/X vssd1 vssd1 vccd1 vccd1
+ _15858_/B sky130_fd_sc_hd__o221a_2
XFILLER_65_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20772__B1 _20775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12668__A _20495_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16440__A1 _19512_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14808_ _14928_/A _14928_/B vssd1 vssd1 vccd1 vccd1 _14814_/C sky130_fd_sc_hd__xnor2_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18576_ _18576_/A _18576_/B vssd1 vssd1 vccd1 vccd1 _18576_/Y sky130_fd_sc_hd__nand2_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _15724_/Y _15725_/Y _15890_/A _15787_/Y vssd1 vssd1 vccd1 vccd1 _16022_/A
+ sky130_fd_sc_hd__o211ai_4
X_17527_ _17537_/A _17537_/B _17527_/C _18059_/B vssd1 vssd1 vccd1 vccd1 _17528_/B
+ sky130_fd_sc_hd__nand4_1
X_14739_ _14734_/X _16749_/C _14738_/X vssd1 vssd1 vccd1 vccd1 _23262_/D sky130_fd_sc_hd__a21o_1
XANTENNA__11804__A2 _11801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17458_ _17454_/Y _17597_/A _17457_/Y vssd1 vssd1 vccd1 vccd1 _17460_/A sky130_fd_sc_hd__o21ai_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15698__B _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16743__A2 _18276_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16409_ _18503_/A vssd1 vssd1 vccd1 vccd1 _17406_/A sky130_fd_sc_hd__buf_4
XFILLER_192_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17389_ _12323_/X _17304_/A _17305_/Y vssd1 vssd1 vccd1 vccd1 _17392_/A sky130_fd_sc_hd__o21ai_1
XFILLER_119_936 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19128_ _19121_/X _19123_/Y _19126_/X vssd1 vssd1 vccd1 vccd1 _19128_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_146_733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13962__C1 _13977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19059_ _19059_/A _19059_/B vssd1 vssd1 vccd1 vccd1 _19060_/B sky130_fd_sc_hd__nand2_2
XANTENNA__13011__B _20798_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19186__A _19186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22070_ _22061_/Y _22054_/A _22015_/X _22016_/X vssd1 vssd1 vccd1 vccd1 _22073_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_195_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12850__B _12850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21021_ _20865_/Y _20870_/X _20754_/X _21015_/X _21006_/Y vssd1 vssd1 vccd1 vccd1
+ _21021_/X sky130_fd_sc_hd__o311a_1
XFILLER_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22972_ _22972_/A vssd1 vssd1 vccd1 vccd1 _23318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14777__B _14777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21923_ _21923_/A vssd1 vssd1 vccd1 vccd1 _22510_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21854_ _21854_/A _21854_/B vssd1 vssd1 vccd1 vccd1 _22455_/A sky130_fd_sc_hd__nor2_2
XFILLER_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13245__A1 _13523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12297__B _12297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20795__A _23299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20805_ _20805_/A _21065_/A _20805_/C vssd1 vssd1 vccd1 vccd1 _20809_/A sky130_fd_sc_hd__nand3_1
XANTENNA__14993__A1 _14879_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21785_ _13616_/Y _13621_/Y _13797_/B _13797_/A vssd1 vssd1 vccd1 vccd1 _21785_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_196_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_858 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23524_ _23538_/CLK _23524_/D vssd1 vssd1 vccd1 vccd1 _23524_/Q sky130_fd_sc_hd__dfxtp_4
X_20736_ _20736_/A _20736_/B vssd1 vssd1 vccd1 vccd1 _20737_/C sky130_fd_sc_hd__nand2_1
XFILLER_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23455_ _23571_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 _23455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20667_ _20667_/A _20667_/B vssd1 vssd1 vccd1 vccd1 _20699_/B sky130_fd_sc_hd__nand2_2
XFILLER_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13202__A _13202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22406_ _22406_/A _22406_/B vssd1 vssd1 vccd1 vccd1 _22406_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18487__A2 _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23386_ _23389_/CLK _23386_/D vssd1 vssd1 vccd1 vccd1 _23386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20598_ _12991_/A _12991_/B _12991_/C _20583_/Y vssd1 vssd1 vccd1 vccd1 _20598_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_100_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23110__S _23110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12463__D _19017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22337_ _22756_/C _22226_/B _22226_/C _22221_/B vssd1 vssd1 vccd1 vccd1 _22356_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_124_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13070_ _13065_/Y _13070_/B _20565_/D vssd1 vssd1 vccd1 vccd1 _13077_/B sky130_fd_sc_hd__nand3b_1
XFILLER_151_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22268_ _22268_/A vssd1 vssd1 vccd1 vccd1 _22566_/B sky130_fd_sc_hd__buf_2
XFILLER_152_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12021_ _12018_/X _12020_/X _18755_/A _18755_/B vssd1 vssd1 vccd1 vccd1 _12021_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_151_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21219_ _21218_/C _21319_/A _21218_/B vssd1 vssd1 vccd1 vccd1 _21219_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_133_994 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22199_ _22199_/A _22290_/B vssd1 vssd1 vccd1 vccd1 _22200_/C sky130_fd_sc_hd__nand2_1
XFILLER_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_622 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19543__B _19543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13872__A _21732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16760_ _16763_/B _16570_/Y _16759_/Y _16765_/A vssd1 vssd1 vccd1 vccd1 _17010_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_24_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13972_ _13972_/A vssd1 vssd1 vccd1 vccd1 _13972_/X sky130_fd_sc_hd__buf_2
XFILLER_46_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15711_ _23420_/Q vssd1 vssd1 vccd1 vccd1 _15712_/D sky130_fd_sc_hd__inv_2
X_12923_ _13138_/C _13138_/D _12923_/C vssd1 vssd1 vccd1 vccd1 _12962_/B sky130_fd_sc_hd__nand3_1
X_16691_ _11766_/B _16686_/A _16911_/A _16911_/B _16900_/A vssd1 vssd1 vccd1 vccd1
+ _16691_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18430_ _18430_/A vssd1 vssd1 vccd1 vccd1 _18430_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15642_ _15642_/A _15931_/A vssd1 vssd1 vccd1 vccd1 _15791_/A sky130_fd_sc_hd__nor2_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _12677_/X _12704_/A _20782_/C _12851_/C vssd1 vssd1 vccd1 vccd1 _12854_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23270__CLK _23492_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _18403_/A _18403_/B _23535_/Q vssd1 vssd1 vccd1 vccd1 _18405_/A sky130_fd_sc_hd__a21oi_1
X_11805_ _11805_/A _11805_/B _11805_/C vssd1 vssd1 vccd1 vccd1 _12297_/B sky130_fd_sc_hd__nand3_2
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15573_ _23509_/Q _15573_/B vssd1 vssd1 vccd1 vccd1 _23497_/D sky130_fd_sc_hd__xnor2_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _12815_/B vssd1 vssd1 vccd1 vccd1 _12785_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17312_ _17150_/B _17140_/Y _16908_/X _17307_/A vssd1 vssd1 vccd1 vccd1 _17313_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14524_ _14535_/A _14538_/A _14538_/B _14538_/C vssd1 vssd1 vccd1 vccd1 _22896_/D
+ sky130_fd_sc_hd__nor4b_2
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18292_ _18292_/A _18292_/B vssd1 vssd1 vccd1 vccd1 _18293_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _11736_/A vssd1 vssd1 vccd1 vccd1 _11764_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17243_ _19949_/A _17243_/B _19674_/B _17243_/D vssd1 vssd1 vccd1 vccd1 _17243_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_30_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14455_ _14430_/D _15238_/C _14430_/A _15094_/C vssd1 vssd1 vccd1 vccd1 _14456_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15933__B1 _15921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11667_ _12024_/B vssd1 vssd1 vccd1 vccd1 _19363_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_128_733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13406_ _21778_/C _22264_/B _13376_/A _13443_/B _13446_/B vssd1 vssd1 vccd1 vccd1
+ _13414_/B sky130_fd_sc_hd__a32o_1
XFILLER_70_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17174_ _16934_/X _16936_/Y _17166_/A vssd1 vssd1 vccd1 vccd1 _17179_/A sky130_fd_sc_hd__o21ai_2
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14386_ _14386_/A _14386_/B _14751_/B _14458_/A vssd1 vssd1 vccd1 vccd1 _14396_/B
+ sky130_fd_sc_hd__nand4_2
X_11598_ _11618_/C vssd1 vssd1 vccd1 vccd1 _11610_/C sky130_fd_sc_hd__clkbuf_2
X_16125_ _16121_/Y _16610_/A _16124_/X vssd1 vssd1 vccd1 vccd1 _16125_/Y sky130_fd_sc_hd__a21oi_1
X_13337_ _13308_/Y _22028_/B _13354_/B vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__a21o_1
XFILLER_182_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16423__A _16423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16056_ _17062_/B vssd1 vssd1 vccd1 vccd1 _16056_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13766__B _13766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13268_ _13766_/A _13766_/B _13268_/C vssd1 vssd1 vccd1 vccd1 _13269_/A sky130_fd_sc_hd__nand3_1
XFILLER_124_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17438__B1 _16027_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15007_ _15124_/A _15124_/B _15013_/C _15013_/D vssd1 vssd1 vccd1 vccd1 _15007_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12219_ _12217_/X _12218_/Y _12198_/B _12199_/A vssd1 vssd1 vccd1 vccd1 _12531_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__15039__A _15208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13199_ _13199_/A _13199_/B vssd1 vssd1 vccd1 vccd1 _13201_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22982__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19815_ _19815_/A _19815_/B vssd1 vssd1 vccd1 vccd1 _19815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11717__D _19648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14267__A3 _14863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19746_ _19598_/B _19598_/C _19598_/A vssd1 vssd1 vccd1 vccd1 _19746_/Y sky130_fd_sc_hd__a21oi_1
X_16958_ _16952_/Y _16955_/X _16961_/C vssd1 vssd1 vccd1 vccd1 _16964_/A sky130_fd_sc_hd__o21bai_2
XFILLER_111_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19172__C _19172_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15909_ _15719_/B _15908_/Y _15721_/X vssd1 vssd1 vccd1 vccd1 _16236_/B sky130_fd_sc_hd__o21ai_1
X_19677_ _19670_/C _19480_/X _19486_/B _19482_/Y vssd1 vssd1 vccd1 vccd1 _19682_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21207__C _21207_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16889_ _16655_/B _16655_/C _16655_/D _16650_/Y vssd1 vssd1 vccd1 vccd1 _16895_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__16413__A1 _16167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16413__B2 _16549_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18628_ _18482_/Y _18487_/X _18465_/A vssd1 vssd1 vccd1 vccd1 _18628_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18559_ _18559_/A _18559_/B vssd1 vssd1 vccd1 vccd1 _18559_/X sky130_fd_sc_hd__and2_1
XFILLER_178_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21570_ _21570_/A vssd1 vssd1 vccd1 vccd1 _21577_/A sky130_fd_sc_hd__inv_2
XFILLER_127_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16177__B1 _16176_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17420__C _19674_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21170__B1 _20786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1055 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20521_ _20501_/X _20509_/Y _20805_/C _12980_/A vssd1 vssd1 vccd1 vccd1 _20521_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_193_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19115__B1 _19116_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23240_ _23240_/A vssd1 vssd1 vccd1 vccd1 _23438_/D sky130_fd_sc_hd__clkbuf_1
X_20452_ _20452_/A _20452_/B _20452_/C vssd1 vssd1 vccd1 vccd1 _20453_/A sky130_fd_sc_hd__and3_1
XANTENNA__19666__A1 _19675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20781__C _20781_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23171_ _23171_/A vssd1 vssd1 vccd1 vccd1 _23407_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13957__A _23501_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20383_ _20411_/A _20383_/B vssd1 vssd1 vccd1 vccd1 _20384_/C sky130_fd_sc_hd__nand2_2
XFILLER_161_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22122_ _22508_/A _22508_/B _22361_/C vssd1 vssd1 vccd1 vccd1 _22122_/Y sky130_fd_sc_hd__nand3_2
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15152__A1 _14184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22053_ _22045_/Y _22046_/Y _22050_/Y _22052_/Y vssd1 vssd1 vccd1 vccd1 _22054_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_82_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21004_ _20857_/Y _20851_/Y _20863_/Y vssd1 vssd1 vccd1 vccd1 _21004_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22973__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19363__B _19363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18641__A2 _19670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19082__C _20368_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__A2 _16523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22955_ _22955_/A vssd1 vssd1 vccd1 vccd1 _23311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21933__C1 _22043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21906_ _21906_/A _22037_/A vssd1 vssd1 vccd1 vccd1 _22043_/A sky130_fd_sc_hd__nand2_2
XFILLER_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22886_ _22882_/X _22873_/Y _22881_/Y vssd1 vssd1 vccd1 vccd1 _22891_/C sky130_fd_sc_hd__o21ai_2
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21837_ _21844_/A _21844_/C vssd1 vssd1 vccd1 vccd1 _21837_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16508__A _16530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23150__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11940__A _16591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12570_ _20628_/C vssd1 vssd1 vccd1 vccd1 _12571_/A sky130_fd_sc_hd__inv_2
X_21768_ _22508_/A _22508_/B _22172_/C _13816_/A _22381_/C vssd1 vssd1 vccd1 vccd1
+ _21984_/A sky130_fd_sc_hd__a32o_2
XFILLER_24_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23507_ _23510_/CLK input41/X vssd1 vssd1 vccd1 vccd1 _23507_/Q sky130_fd_sc_hd__dfxtp_1
X_20719_ _20512_/A _20512_/B _20518_/X _20695_/B _20695_/C vssd1 vssd1 vccd1 vccd1
+ _20719_/X sky130_fd_sc_hd__o2111a_1
XFILLER_180_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21699_ _21716_/B _21716_/C _23574_/Q vssd1 vssd1 vccd1 vccd1 _21717_/A sky130_fd_sc_hd__a21boi_2
XFILLER_141_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14240_ _14911_/C vssd1 vssd1 vccd1 vccd1 _15356_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__19657__A1 _19304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23438_ _23441_/CLK _23438_/D vssd1 vssd1 vccd1 vccd1 _23438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20267__A2 _20055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14171_ _14133_/B _14121_/Y _14116_/X _14118_/X vssd1 vssd1 vccd1 vccd1 _14180_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_164_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23369_ _23401_/CLK _23369_/D vssd1 vssd1 vccd1 vccd1 _23369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_831 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11952__A1 _11948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13122_ _13166_/A _13122_/B vssd1 vssd1 vccd1 vccd1 _13124_/C sky130_fd_sc_hd__nor2_1
XFILLER_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17930_ _17922_/X _17924_/X _17925_/Y vssd1 vssd1 vccd1 vccd1 _17930_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_127_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _13058_/B vssd1 vssd1 vccd1 vccd1 _13053_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_152_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_994 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22964__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ _16032_/A vssd1 vssd1 vccd1 vccd1 _12004_/X sky130_fd_sc_hd__buf_4
XFILLER_61_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17861_ _17760_/B _17858_/Y _17859_/Y _17860_/Y vssd1 vssd1 vccd1 vccd1 _17863_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18632__A2 _11865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14698__A _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19600_ _19600_/A vssd1 vssd1 vccd1 vccd1 _19600_/Y sky130_fd_sc_hd__inv_2
X_16812_ _16812_/A _16812_/B vssd1 vssd1 vccd1 vccd1 _16814_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17792_ _17792_/A _17792_/B _17792_/C vssd1 vssd1 vccd1 vccd1 _17798_/C sky130_fd_sc_hd__nand3_1
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1012 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19531_ _18859_/C _17443_/A _17444_/A _17972_/A _12343_/A vssd1 vssd1 vccd1 vccd1
+ _19534_/A sky130_fd_sc_hd__a32o_1
XANTENNA__11834__B _11834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16743_ _16480_/X _18276_/C _16194_/C _16192_/X _16183_/X vssd1 vssd1 vccd1 vccd1
+ _16784_/A sky130_fd_sc_hd__o32a_1
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13955_ _23502_/Q vssd1 vssd1 vccd1 vccd1 _14796_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19462_ _19456_/B _19456_/A _19636_/A vssd1 vssd1 vccd1 vccd1 _19635_/A sky130_fd_sc_hd__a21o_1
X_12906_ _12896_/B _12896_/C _12896_/A vssd1 vssd1 vccd1 vccd1 _12906_/Y sky130_fd_sc_hd__a21oi_4
X_16674_ _16674_/A _19011_/A _17108_/B _17098_/B vssd1 vssd1 vccd1 vccd1 _16674_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _14024_/B vssd1 vssd1 vccd1 vccd1 _13939_/A sky130_fd_sc_hd__buf_2
XFILLER_61_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18413_ _18413_/A _18413_/B vssd1 vssd1 vccd1 vccd1 _18414_/B sky130_fd_sc_hd__xor2_1
XFILLER_146_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15625_ _15761_/A _16187_/C _15631_/B _15637_/D vssd1 vssd1 vccd1 vccd1 _15644_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19393_ _19601_/A _19601_/B _19468_/A _19600_/A vssd1 vssd1 vccd1 vccd1 _19393_/Y
+ sky130_fd_sc_hd__a22oi_2
X_12837_ _12837_/A _12837_/B vssd1 vssd1 vccd1 vccd1 _12904_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23141__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22139__B _22139_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12968__B1 _21295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18344_ _18344_/A _18344_/B vssd1 vssd1 vccd1 vccd1 _18346_/A sky130_fd_sc_hd__or2_1
XFILLER_187_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15556_ _15556_/A _15564_/B vssd1 vssd1 vccd1 vccd1 _15558_/B sky130_fd_sc_hd__xor2_2
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _20670_/C vssd1 vssd1 vccd1 vccd1 _13179_/A sky130_fd_sc_hd__buf_2
XFILLER_159_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _15964_/B vssd1 vssd1 vccd1 vccd1 _16462_/D sky130_fd_sc_hd__clkbuf_2
X_18275_ _20265_/C _18211_/C _18272_/X _18274_/X vssd1 vssd1 vccd1 vccd1 _18275_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19360__A3 _19357_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ _11969_/B _11907_/B _11908_/A vssd1 vssd1 vccd1 vccd1 _11719_/X sky130_fd_sc_hd__or3_1
XFILLER_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15906__B1 _15618_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15487_ _15511_/C _15485_/D _15483_/X _15486_/Y vssd1 vssd1 vccd1 vccd1 _15493_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12699_ _20663_/C vssd1 vssd1 vccd1 vccd1 _21054_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_675 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17226_ _19840_/A _17860_/A _19664_/B _17226_/D vssd1 vssd1 vccd1 vccd1 _17236_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_35_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput10 wb_dat_i[12] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_4
X_14438_ _14438_/A _14438_/B vssd1 vssd1 vccd1 vccd1 _14443_/B sky130_fd_sc_hd__nor2_1
Xinput21 wb_dat_i[22] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
Xinput32 wb_dat_i[3] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_8
Xinput43 x[11] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__19112__A3 _18778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17157_ _17154_/X _17155_/X _17152_/B _17161_/B vssd1 vssd1 vccd1 vccd1 _17220_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_122_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14369_ _14420_/A _14422_/B _14422_/C vssd1 vssd1 vccd1 vccd1 _14369_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__12681__A _23447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16153__A _16153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_736 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11943__A1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16108_ _16108_/A _16108_/B _16108_/C vssd1 vssd1 vccd1 vccd1 _16581_/A sky130_fd_sc_hd__nand3_2
X_17088_ _17068_/X _17069_/X _17070_/X _20049_/A _17454_/B vssd1 vssd1 vccd1 vccd1
+ _17089_/D sky130_fd_sc_hd__o2111ai_4
XFILLER_116_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16039_ _16039_/A vssd1 vssd1 vccd1 vccd1 _16309_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18623__A2 _18778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19729_ _19560_/Y _19728_/X _19719_/Y _19893_/A vssd1 vssd1 vccd1 vccd1 _19730_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21915__C1 _22043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17712__A _17712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22740_ _22738_/A _22738_/B _23280_/Q vssd1 vssd1 vccd1 vccd1 _22740_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_93_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22671_ _22671_/A _22720_/A _22671_/C _22671_/D vssd1 vssd1 vccd1 vccd1 _22720_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_164_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23132__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__A _11760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21622_ _21616_/A _21617_/A _21614_/Y _21630_/A vssd1 vssd1 vccd1 vccd1 _21622_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21553_ _21554_/D _21358_/A _21358_/B _21554_/B _21554_/C vssd1 vssd1 vccd1 vccd1
+ _21555_/A sky130_fd_sc_hd__a32o_1
XANTENNA__20497__A2 _23296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_675 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20504_ _20504_/A vssd1 vssd1 vccd1 vccd1 _20504_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__15373__A1 _15310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21484_ _21484_/A _23568_/Q _21484_/C vssd1 vssd1 vccd1 vccd1 _21485_/B sky130_fd_sc_hd__nand3_2
XFILLER_119_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15373__B2 _15371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22238__A3 _22090_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23223_ _23223_/A vssd1 vssd1 vccd1 vccd1 _23430_/D sky130_fd_sc_hd__clkbuf_1
X_20435_ _20446_/B _20446_/C _20446_/A vssd1 vssd1 vccd1 vccd1 _20449_/A sky130_fd_sc_hd__a21o_1
XFILLER_14_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11934__A1 _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23154_ _23400_/Q input16/X _23156_/S vssd1 vssd1 vccd1 vccd1 _23155_/A sky130_fd_sc_hd__mux2_1
X_20366_ _20366_/A _20366_/B _20366_/C _20368_/C vssd1 vssd1 vccd1 vccd1 _20366_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_162_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22105_ _22102_/A _22240_/B _22102_/C vssd1 vssd1 vccd1 vccd1 _22439_/D sky130_fd_sc_hd__a21o_1
XFILLER_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23085_ _23085_/A vssd1 vssd1 vccd1 vccd1 _23369_/D sky130_fd_sc_hd__clkbuf_1
X_20297_ _20243_/A _20243_/B _20295_/X _20296_/Y vssd1 vssd1 vccd1 vccd1 _20298_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22036_ _22025_/Y _22032_/Y _22035_/X vssd1 vssd1 vccd1 vccd1 _22036_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18614__A2 _18604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_986 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11935__A _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13740_ _13738_/X _13739_/Y _13686_/A _22465_/D vssd1 vssd1 vccd1 vccd1 _13744_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22938_ _23304_/Q input16/X _22940_/S vssd1 vssd1 vccd1 vccd1 _22939_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13671_ _13671_/A _13671_/B _13671_/C vssd1 vssd1 vccd1 vccd1 _13676_/B sky130_fd_sc_hd__nand3_1
XFILLER_32_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22869_ _22859_/Y _22849_/X _22828_/A _22828_/B _22868_/Y vssd1 vssd1 vccd1 vccd1
+ _22869_/Y sky130_fd_sc_hd__a41oi_4
XANTENNA__23123__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_88 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15410_ _15225_/B _15254_/C _15254_/A _15366_/Y _15379_/A vssd1 vssd1 vccd1 vccd1
+ _15412_/A sky130_fd_sc_hd__a311oi_1
X_12622_ _12687_/A vssd1 vssd1 vccd1 vccd1 _12622_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16390_ _16389_/X _16322_/B _16402_/B _16323_/A vssd1 vssd1 vccd1 vccd1 _16395_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_169_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17889__B1 _17406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15341_ _15442_/D _15528_/A _15442_/B vssd1 vssd1 vccd1 vccd1 _15344_/A sky130_fd_sc_hd__or3_1
X_12553_ _18557_/B _12523_/B _12528_/A _12528_/B vssd1 vssd1 vccd1 vccd1 _12553_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14981__A _15353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_956 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18060_ _18060_/A _18060_/B vssd1 vssd1 vccd1 vccd1 _18060_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15272_ _15192_/B _15192_/A _15271_/Y _15190_/A vssd1 vssd1 vccd1 vccd1 _15272_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16561__B1 _16560_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12484_ _12484_/A _12484_/B vssd1 vssd1 vccd1 vccd1 _12484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12178__A1 _15882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18172__B _20151_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17011_ _17011_/A _17011_/B _17011_/C vssd1 vssd1 vccd1 vccd1 _17012_/C sky130_fd_sc_hd__nand3_1
XFILLER_144_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21437__A1 _20957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14223_ _14222_/Y _14218_/A _14217_/C vssd1 vssd1 vccd1 vccd1 _14224_/C sky130_fd_sc_hd__a21boi_1
XFILLER_125_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18838__C1 _19543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17105__A2 _15655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14154_ _14153_/Y _14152_/X _14003_/A _14253_/B vssd1 vssd1 vccd1 vccd1 _14154_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_152_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13105_ _12978_/Y _12984_/B _12984_/A vssd1 vssd1 vccd1 vccd1 _13147_/A sky130_fd_sc_hd__o21ai_1
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18962_ _19410_/A _18944_/Y _18950_/Y vssd1 vssd1 vccd1 vccd1 _18964_/B sky130_fd_sc_hd__a21o_1
XFILLER_152_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _14980_/A _14068_/X _14069_/X _14083_/Y _14084_/X vssd1 vssd1 vccd1 vccd1
+ _14139_/A sky130_fd_sc_hd__a32o_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14875__B1 _15120_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17913_ _17796_/Y _17786_/Y _17779_/Y vssd1 vssd1 vccd1 vccd1 _17913_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_140_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11689__B1 _11665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13036_ _12952_/X _13025_/X _13041_/B _13022_/Y _20955_/C vssd1 vssd1 vccd1 vccd1
+ _13036_/X sky130_fd_sc_hd__o2111a_1
X_18893_ _18893_/A _18893_/B _18893_/C vssd1 vssd1 vccd1 vccd1 _18897_/D sky130_fd_sc_hd__nand3_2
XFILLER_121_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1043 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16616__A1 _12509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17844_ _17972_/A vssd1 vssd1 vccd1 vccd1 _19799_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_113_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17775_ _17781_/A _17838_/C _17782_/B _17782_/C vssd1 vssd1 vccd1 vccd1 _17779_/A
+ sky130_fd_sc_hd__a22o_1
X_14987_ _15262_/A _15010_/A vssd1 vssd1 vccd1 vccd1 _14987_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22165__A2 _22754_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19514_ _19514_/A _19514_/B _19514_/C vssd1 vssd1 vccd1 vccd1 _19525_/D sky130_fd_sc_hd__nand3_4
X_16726_ _16243_/A _16246_/C _16725_/Y vssd1 vssd1 vccd1 vccd1 _16735_/C sky130_fd_sc_hd__a21oi_2
X_13938_ _13908_/C _13937_/X _13911_/C _13901_/B vssd1 vssd1 vccd1 vccd1 _13994_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16919__A2 _16665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19445_ _19442_/Y _19443_/Y _19444_/X vssd1 vssd1 vccd1 vccd1 _19625_/B sky130_fd_sc_hd__o21ai_2
XFILLER_35_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16657_ _23427_/Q _16657_/B vssd1 vssd1 vccd1 vccd1 _17029_/A sky130_fd_sc_hd__nand2_2
X_13869_ _21856_/C _21856_/D _13763_/A _13763_/B vssd1 vssd1 vccd1 vccd1 _13870_/B
+ sky130_fd_sc_hd__a22oi_4
XANTENNA__16148__A _17431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__A _23589_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15608_ _15729_/A vssd1 vssd1 vccd1 vccd1 _15931_/A sky130_fd_sc_hd__buf_2
X_19376_ _19376_/A _19387_/A vssd1 vssd1 vccd1 vccd1 _19385_/A sky130_fd_sc_hd__nand2_1
X_16588_ _12222_/X _12223_/X _15883_/A vssd1 vssd1 vccd1 vccd1 _16588_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20893__A _23300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18327_ _20366_/A _18376_/B _18274_/X _18277_/C vssd1 vssd1 vccd1 vccd1 _18338_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_148_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _15539_/A _15539_/B vssd1 vssd1 vccd1 vccd1 _15540_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18363__A _23533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _18364_/A _18364_/B _23533_/Q vssd1 vssd1 vccd1 vccd1 _18319_/A sky130_fd_sc_hd__a21o_1
XFILLER_175_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14158__A2 _15019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_926 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17209_ _17943_/A _17374_/C _17208_/Y _16987_/A vssd1 vssd1 vccd1 vccd1 _17212_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_128_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18189_ _18298_/A _18298_/B _18134_/C _18209_/A vssd1 vssd1 vccd1 vccd1 _18191_/A
+ sky130_fd_sc_hd__o211ai_1
X_20220_ _20146_/C _20148_/A _20216_/X _20218_/Y vssd1 vssd1 vccd1 vccd1 _20220_/Y
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__16314__C _16314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16304__B1 _15742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16855__A1 _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20151_ _20151_/A _20151_/B _20151_/C _20151_/D vssd1 vssd1 vccd1 vccd1 _20158_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_144_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20082_ _18016_/C _19862_/B _19862_/C _20164_/C _20269_/C vssd1 vssd1 vccd1 vccd1
+ _20083_/B sky130_fd_sc_hd__a32o_1
XFILLER_44_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19006__C1 _19703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19557__B1 _19203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22156__A2 _22164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ _20984_/A _20984_/B _20984_/C vssd1 vssd1 vccd1 vccd1 _21111_/A sky130_fd_sc_hd__nand3_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17568__C1 _17567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22723_ _22723_/A _22723_/B vssd1 vssd1 vccd1 vccd1 _22726_/A sky130_fd_sc_hd__or2_1
XFILLER_14_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16058__A _16058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22654_ _22643_/A _22712_/A _22712_/B vssd1 vssd1 vccd1 vccd1 _22656_/A sky130_fd_sc_hd__a21bo_1
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21605_ _21645_/B _21605_/B _21605_/C vssd1 vssd1 vccd1 vccd1 _21666_/A sky130_fd_sc_hd__or3_2
X_22585_ _22559_/X _22478_/X _22580_/Y _22581_/X vssd1 vssd1 vccd1 vccd1 _22585_/Y
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__18273__A _20210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21536_ _21484_/C _21484_/A _23568_/Q vssd1 vssd1 vccd1 vccd1 _21536_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_166_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13357__B1 _13802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22226__C _22226_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21467_ _21465_/X _21467_/B vssd1 vssd1 vccd1 vccd1 _21468_/B sky130_fd_sc_hd__and2b_1
XFILLER_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20418_ _20419_/B _23556_/Q vssd1 vssd1 vccd1 vccd1 _20418_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17099__B2 _15655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23206_ _14599_/X input38/X _23206_/S vssd1 vssd1 vccd1 vccd1 _23207_/A sky130_fd_sc_hd__mux2_1
X_21398_ _21424_/A _21424_/B _21399_/C vssd1 vssd1 vccd1 vccd1 _21400_/A sky130_fd_sc_hd__o21bai_1
XFILLER_104_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20349_ _20356_/A _20356_/B _23554_/Q vssd1 vssd1 vccd1 vccd1 _20359_/D sky130_fd_sc_hd__nand3_1
XFILLER_175_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23137_ _18997_/A input8/X _23145_/S vssd1 vssd1 vccd1 vccd1 _23138_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23068_ _23068_/A vssd1 vssd1 vccd1 vccd1 _23361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12332__A1 _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17256__D1 _17450_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22019_ _23331_/Q vssd1 vssd1 vccd1 vccd1 _22021_/A sky130_fd_sc_hd__inv_2
X_14910_ _14777_/A _14911_/B _14777_/C _14793_/C _14791_/B vssd1 vssd1 vccd1 vccd1
+ _14910_/X sky130_fd_sc_hd__a32o_1
XANTENNA__11665__A _11665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15890_ _15890_/A _15890_/B vssd1 vssd1 vccd1 vccd1 _15890_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_336 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17271__A1 _16447_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22896__C input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A wb_dat_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ _14306_/A _14306_/B _14306_/C _14310_/A vssd1 vssd1 vccd1 vccd1 _14842_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14085__A1 _14980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_870 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17560_ _17806_/B _17556_/X _17559_/Y vssd1 vssd1 vccd1 vccd1 _17667_/A sky130_fd_sc_hd__o21ai_1
XFILLER_112_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14772_ _14774_/B vssd1 vssd1 vccd1 vccd1 _14990_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11984_ _11757_/A _18812_/B _18470_/C _18468_/A vssd1 vssd1 vccd1 vccd1 _12426_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16511_ _16510_/C _18017_/D _16539_/A _16539_/B vssd1 vssd1 vccd1 vccd1 _16532_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13723_ _13717_/Y _13723_/B _13723_/C vssd1 vssd1 vccd1 vccd1 _13723_/Y sky130_fd_sc_hd__nand3b_1
X_17491_ _17663_/A _17663_/B _17497_/C _17497_/D vssd1 vssd1 vccd1 vccd1 _17491_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19230_ _19230_/A _19230_/B vssd1 vssd1 vccd1 vccd1 _19240_/A sky130_fd_sc_hd__nand2_1
XFILLER_95_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16442_ _15884_/A _12373_/A _11898_/X _16311_/X vssd1 vssd1 vccd1 vccd1 _16445_/A
+ sky130_fd_sc_hd__o22ai_4
X_13654_ _13647_/X _13648_/Y _13649_/Y _13653_/Y vssd1 vssd1 vccd1 vccd1 _13655_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19315__A3 _19491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19161_ _19161_/A _19651_/A _19163_/A vssd1 vssd1 vccd1 vccd1 _19162_/B sky130_fd_sc_hd__and3_1
X_12605_ _12873_/C _12678_/C vssd1 vssd1 vccd1 vccd1 _12606_/B sky130_fd_sc_hd__nor2_1
XANTENNA__19279__A _19279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _11871_/A _15698_/A _15698_/B _18461_/A _15972_/X vssd1 vssd1 vccd1 vccd1
+ _16374_/A sky130_fd_sc_hd__o32ai_2
XFILLER_9_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13585_/A vssd1 vssd1 vccd1 vccd1 _13686_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_197_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18112_ _18109_/Y _18110_/X _18022_/B _18028_/B vssd1 vssd1 vccd1 vccd1 _18114_/D
+ sky130_fd_sc_hd__o211ai_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15324_ _15324_/A _15324_/B _15380_/A _15323_/X vssd1 vssd1 vccd1 vccd1 _15380_/B
+ sky130_fd_sc_hd__or4bb_2
XFILLER_185_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19092_ _19090_/Y _18915_/Y _19091_/Y vssd1 vssd1 vccd1 vccd1 _19094_/B sky130_fd_sc_hd__a21oi_1
X_12536_ _12536_/A _12536_/B vssd1 vssd1 vccd1 vccd1 _12537_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18043_ _18043_/A _18043_/B _18043_/C vssd1 vssd1 vccd1 vccd1 _18132_/B sky130_fd_sc_hd__and3_2
XFILLER_184_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15255_ _15255_/A _15255_/B vssd1 vssd1 vccd1 vccd1 _15303_/D sky130_fd_sc_hd__nand2_1
XFILLER_172_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12467_ _16122_/A _16122_/B _18755_/A _18755_/B vssd1 vssd1 vccd1 vccd1 _18675_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_172_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output92_A _23266_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ _14017_/X _14050_/A _14089_/Y vssd1 vssd1 vccd1 vccd1 _14312_/C sky130_fd_sc_hd__a21oi_2
XFILLER_193_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15186_ _15250_/A _15187_/C _15249_/A vssd1 vssd1 vccd1 vccd1 _15188_/C sky130_fd_sc_hd__a21o_1
X_12398_ _12563_/B _12398_/B _12398_/C _12546_/A vssd1 vssd1 vccd1 vccd1 _19089_/A
+ sky130_fd_sc_hd__nand4b_4
XFILLER_153_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21291__C1 _21431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ _14137_/A _14137_/B _14137_/C vssd1 vssd1 vccd1 vccd1 _14138_/A sky130_fd_sc_hd__nand3_1
X_19994_ _19987_/Y _19991_/Y _19993_/X vssd1 vssd1 vccd1 vccd1 _19996_/B sky130_fd_sc_hd__a21o_1
XFILLER_141_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18945_ _19381_/B _19113_/C _18945_/C _19262_/A vssd1 vssd1 vccd1 vccd1 _18945_/Y
+ sky130_fd_sc_hd__nand4_1
X_14068_ _14068_/A vssd1 vssd1 vccd1 vccd1 _14068_/X sky130_fd_sc_hd__buf_2
XFILLER_67_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13019_ _20897_/C _13019_/B _13019_/C _20798_/C vssd1 vssd1 vccd1 vccd1 _13019_/Y
+ sky130_fd_sc_hd__nand4_4
X_18876_ _18875_/C _18875_/A _18875_/B vssd1 vssd1 vccd1 vccd1 _18884_/A sky130_fd_sc_hd__a21oi_4
XFILLER_95_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20888__A _21121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17827_ _18072_/D _18072_/C _18253_/B _18256_/A vssd1 vssd1 vccd1 vccd1 _17828_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__22138__A2 _22139_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13790__A _22064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17262__A _18607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17758_ _17773_/B _17773_/C _17773_/D vssd1 vssd1 vccd1 vccd1 _17758_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__19180__C _19180_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16709_ _16709_/A _16709_/B _16709_/C vssd1 vssd1 vccd1 vccd1 _16956_/A sky130_fd_sc_hd__nand3_2
XFILLER_63_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17689_ _17945_/A _17945_/B _17693_/A vssd1 vssd1 vccd1 vccd1 _17689_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19428_ _19428_/A _19616_/A vssd1 vssd1 vccd1 vccd1 _19428_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14379__A2 _15358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19359_ _18673_/A _17846_/X _19358_/Y vssd1 vssd1 vccd1 vccd1 _19614_/B sky130_fd_sc_hd__o21ai_2
XFILLER_148_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18093__A _18093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17317__A2 _16055_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22370_ _22366_/Y _22370_/B _22496_/B vssd1 vssd1 vccd1 vccd1 _22409_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__16525__B1 _16526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21321_ _21319_/B _21215_/C _21215_/A vssd1 vssd1 vccd1 vccd1 _21321_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_159_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21252_ _21012_/X _21251_/Y _21237_/Y _21154_/Y vssd1 vssd1 vccd1 vccd1 _21253_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_117_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20203_ _20203_/A _20203_/B vssd1 vssd1 vccd1 vccd1 _23531_/D sky130_fd_sc_hd__xor2_1
XFILLER_117_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_503 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21183_ _12571_/X _21592_/A _21178_/C vssd1 vssd1 vccd1 vccd1 _21184_/D sky130_fd_sc_hd__o21ai_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20134_ _20134_/A vssd1 vssd1 vccd1 vccd1 _20151_/D sky130_fd_sc_hd__buf_2
XANTENNA__16698__D _16706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20065_ _20066_/C _20066_/A _20066_/B vssd1 vssd1 vccd1 vccd1 _20067_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__19652__A _19652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17789__C1 _19862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20798__A _20798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17253__B2 _17565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22129__A2 _22126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15803__A2 _15800_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17005__A1 _23519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_851 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ _20967_/A _20967_/B vssd1 vssd1 vccd1 vccd1 _21101_/C sky130_fd_sc_hd__nand2_1
XFILLER_54_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17410__D1 _17233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22706_ _22701_/A _22701_/B _22830_/A _22754_/B vssd1 vssd1 vccd1 vccd1 _22754_/C
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _20902_/A _23300_/Q _21047_/B vssd1 vssd1 vccd1 vccd1 _21174_/C sky130_fd_sc_hd__nand3_2
XFILLER_198_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22637_ _22637_/A _22637_/B _22637_/C vssd1 vssd1 vccd1 vccd1 _22637_/Y sky130_fd_sc_hd__nand3_1
XFILLER_110_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17308__A2 _17305_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18505__A1 _12214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22301__A2 _13599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _21905_/B vssd1 vssd1 vccd1 vccd1 _13486_/A sky130_fd_sc_hd__clkinv_2
XFILLER_194_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22568_ _22057_/X _22168_/X _22361_/C _22392_/A vssd1 vssd1 vccd1 vccd1 _22577_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_16_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12321_ _12321_/A vssd1 vssd1 vccd1 vccd1 _12381_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_155_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21519_ _21468_/A _21467_/B _21465_/X vssd1 vssd1 vccd1 vccd1 _21521_/A sky130_fd_sc_hd__a21oi_1
XFILLER_166_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22499_ _22499_/A _22499_/B _22499_/C vssd1 vssd1 vccd1 vccd1 _22513_/A sky130_fd_sc_hd__nand3_1
XFILLER_5_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15040_ _14926_/A _14926_/C _15037_/Y vssd1 vssd1 vccd1 vccd1 _15041_/B sky130_fd_sc_hd__a21oi_1
X_12252_ _12254_/A _12253_/A _12251_/X vssd1 vssd1 vccd1 vccd1 _12300_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12002__B1 _16198_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15566__S _15566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12183_ _12183_/A _12187_/A _19539_/A _16674_/A vssd1 vssd1 vccd1 vccd1 _12183_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_135_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17066__B _19700_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16991_ _17217_/A _17218_/A vssd1 vssd1 vccd1 vccd1 _17011_/C sky130_fd_sc_hd__or2_1
XFILLER_96_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18730_ _19089_/A _12545_/Y _19089_/B _19090_/C vssd1 vssd1 vccd1 vccd1 _18909_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_122_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15942_ _15948_/A _16246_/B _15948_/C vssd1 vssd1 vccd1 vccd1 _16003_/A sky130_fd_sc_hd__nand3_1
XFILLER_49_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17244__A1 _19957_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18661_ _12113_/X _18660_/X _11686_/Y _19011_/A _11849_/C vssd1 vssd1 vccd1 vccd1
+ _18662_/B sky130_fd_sc_hd__o311a_1
XANTENNA__18441__B1 _18788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _19700_/C vssd1 vssd1 vccd1 vccd1 _19363_/C sky130_fd_sc_hd__buf_2
XFILLER_37_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15017__D _15017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ _17610_/X _17611_/X _17589_/Y _17597_/Y vssd1 vssd1 vccd1 vccd1 _17612_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__21591__A3 _21432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14824_ _14825_/A _14825_/B _14825_/C vssd1 vssd1 vccd1 vccd1 _14824_/X sky130_fd_sc_hd__a21o_1
XFILLER_92_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _23539_/Q _18733_/A _18589_/Y _18590_/X vssd1 vssd1 vccd1 vccd1 _18593_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ _17478_/X _17477_/Y _17290_/A _17486_/Y _17488_/X vssd1 vssd1 vccd1 vccd1
+ _17543_/X sky130_fd_sc_hd__o2111a_1
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11816__B1 _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14755_ _14174_/B _14887_/A _14753_/Y _14754_/X vssd1 vssd1 vccd1 vccd1 _14762_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _11967_/A _11967_/B _11967_/C vssd1 vssd1 vccd1 vccd1 _11968_/A sky130_fd_sc_hd__nand3_1
XANTENNA__21035__C _21035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17547__A2 _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16204__C1 _19165_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ _22159_/C vssd1 vssd1 vccd1 vccd1 _22192_/C sky130_fd_sc_hd__clkbuf_2
X_17474_ _17473_/A _17473_/B _17473_/C _17473_/D vssd1 vssd1 vccd1 vccd1 _17475_/C
+ sky130_fd_sc_hd__a22o_1
X_14686_ _23372_/Q _14667_/X _14685_/X vssd1 vssd1 vccd1 vccd1 _14686_/X sky130_fd_sc_hd__o21a_1
X_11898_ _18461_/A vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__buf_4
XFILLER_189_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19213_ _19202_/Y _19212_/Y _19205_/X vssd1 vssd1 vccd1 vccd1 _19213_/Y sky130_fd_sc_hd__o21ai_1
X_16425_ _16425_/A _16425_/B _16425_/C vssd1 vssd1 vccd1 vccd1 _16425_/Y sky130_fd_sc_hd__nand3_1
X_13637_ _13495_/X _13313_/X _13630_/B _13634_/X _13636_/X vssd1 vssd1 vccd1 vccd1
+ _13637_/X sky130_fd_sc_hd__o311a_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19144_ _18944_/C _19141_/Y _19410_/B vssd1 vssd1 vccd1 vccd1 _19144_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16356_ _16356_/A vssd1 vssd1 vccd1 vccd1 _16356_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13568_ _22474_/A _13471_/A _21892_/A _13487_/Y _13482_/Y vssd1 vssd1 vccd1 vccd1
+ _13569_/C sky130_fd_sc_hd__o221ai_2
XFILLER_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15307_ _15363_/D _15109_/X _15110_/X _15308_/A _15308_/D vssd1 vssd1 vccd1 vccd1
+ _15311_/A sky130_fd_sc_hd__a32o_1
XFILLER_172_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19075_ _19075_/A _19075_/B _19075_/C vssd1 vssd1 vccd1 vccd1 _19087_/B sky130_fd_sc_hd__nand3_2
X_12519_ _12374_/A _12509_/X _12518_/X _12089_/A vssd1 vssd1 vccd1 vccd1 _12520_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16287_ _17108_/B vssd1 vssd1 vccd1 vccd1 _17845_/C sky130_fd_sc_hd__buf_2
X_13499_ _13663_/C vssd1 vssd1 vccd1 vccd1 _13709_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18026_ _18026_/A _18026_/B vssd1 vssd1 vccd1 vccd1 _18033_/A sky130_fd_sc_hd__nand2_1
XFILLER_161_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15238_ _15369_/A _15369_/B _15238_/C vssd1 vssd1 vccd1 vccd1 _15238_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__15730__A1 _15864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17468__D1 _18172_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15169_ _15369_/A _15369_/B vssd1 vssd1 vccd1 vccd1 _15375_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19977_ _19977_/A _19977_/B vssd1 vssd1 vccd1 vccd1 _19977_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18928_ _17050_/X _16819_/X _16804_/A _16804_/B _19082_/B vssd1 vssd1 vccd1 vccd1
+ _18928_/X sky130_fd_sc_hd__a221o_4
XFILLER_80_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19903__C _19903_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20411__A _20411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18859_ _18859_/A _18859_/B _18859_/C _18859_/D vssd1 vssd1 vccd1 vccd1 _18859_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_95_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18088__A _18163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15505__A _15527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21870_ _13741_/B _13741_/C _22236_/A vssd1 vssd1 vccd1 vccd1 _21874_/A sky130_fd_sc_hd__a21o_1
XFILLER_36_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20821_ _12689_/X _12850_/B _12827_/A _12692_/Y vssd1 vssd1 vccd1 vccd1 _20821_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23540_ _23566_/CLK _23540_/D vssd1 vssd1 vccd1 vccd1 _23540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20752_ _21157_/A _20752_/B vssd1 vssd1 vccd1 vccd1 _21011_/A sky130_fd_sc_hd__and2_1
XFILLER_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18940__A_N _18944_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23471_ _23499_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 _23471_/Q sky130_fd_sc_hd__dfxtp_4
X_20683_ _20509_/Y _20682_/Y _20678_/Y _20679_/Y vssd1 vssd1 vccd1 vccd1 _20683_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22422_ _22419_/Y _22421_/X _22237_/A _13431_/X vssd1 vssd1 vccd1 vccd1 _22428_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22353_ _23275_/Q _22353_/B vssd1 vssd1 vccd1 vccd1 _22452_/B sky130_fd_sc_hd__nor2_1
XFILLER_163_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21304_ _21300_/X _21301_/X _21173_/X _21303_/X vssd1 vssd1 vccd1 vccd1 _21307_/D
+ sky130_fd_sc_hd__o211ai_4
XFILLER_124_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23169__A _23169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22284_ _13465_/X _22059_/X _22283_/X vssd1 vssd1 vccd1 vccd1 _22284_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21235_ _21229_/Y _21333_/B _21233_/X vssd1 vssd1 vccd1 vccd1 _21236_/B sky130_fd_sc_hd__o21ai_2
XFILLER_105_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16071__A _16075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21166_ _21164_/X _21162_/Y _21387_/C _12981_/C vssd1 vssd1 vccd1 vccd1 _21166_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_85_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20117_ _20207_/B vssd1 vssd1 vccd1 vccd1 _20117_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16682__C1 _17149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19215__A2 _19179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12104__A _18756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21097_ _21097_/A _21097_/B _21097_/C vssd1 vssd1 vccd1 vccd1 _21097_/X sky130_fd_sc_hd__and3_1
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20048_ _17593_/X _17591_/X _17595_/X _20215_/B _20215_/C vssd1 vssd1 vccd1 vccd1
+ _20048_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23108__S _23110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15415__A _15415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _12688_/B _12756_/B _12875_/B vssd1 vssd1 vccd1 vccd1 _12871_/A sky130_fd_sc_hd__a21o_1
XFILLER_171_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _12144_/A vssd1 vssd1 vccd1 vccd1 _11822_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21999_ _21884_/B _21996_/Y _22476_/C _21877_/A _21998_/Y vssd1 vssd1 vccd1 vccd1
+ _21999_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14298_/C _14545_/A _14539_/X _19261_/C vssd1 vssd1 vccd1 vccd1 _14540_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12471__B1 _18506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _23386_/Q vssd1 vssd1 vccd1 vccd1 _11977_/B sky130_fd_sc_hd__buf_2
XFILLER_57_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16201__A2 _16319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14471_ _14377_/A _15233_/C _14835_/C _14469_/C vssd1 vssd1 vccd1 vccd1 _14472_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _12260_/C vssd1 vssd1 vccd1 vccd1 _18945_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_42_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _15902_/B _16202_/Y _16209_/Y vssd1 vssd1 vccd1 vccd1 _16217_/A sky130_fd_sc_hd__o21ai_1
X_13422_ _13453_/A vssd1 vssd1 vccd1 vccd1 _13430_/A sky130_fd_sc_hd__buf_2
XFILLER_174_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17190_ _16955_/X _17185_/Y _17189_/Y vssd1 vssd1 vccd1 vccd1 _17190_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__19151__A1 _19149_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _16141_/A _16795_/A _16620_/C _16141_/D vssd1 vssd1 vccd1 vccd1 _16142_/B
+ sky130_fd_sc_hd__nand4_2
X_13353_ _23325_/Q vssd1 vssd1 vccd1 vccd1 _13783_/C sky130_fd_sc_hd__inv_2
XFILLER_139_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17162__B1 _17154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18461__A _18461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12304_ _19082_/A _12237_/X _12289_/B _12547_/A _12303_/Y vssd1 vssd1 vccd1 vccd1
+ _12304_/X sky130_fd_sc_hd__o311a_1
X_16072_ _16062_/Y _16063_/X _16469_/A _16071_/Y vssd1 vssd1 vccd1 vccd1 _16072_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_182_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13284_ _13634_/A _13634_/B _22280_/B vssd1 vssd1 vccd1 vccd1 _13284_/Y sky130_fd_sc_hd__nand3_1
X_19900_ _19900_/A _20369_/A _19967_/A _19900_/D vssd1 vssd1 vccd1 vccd1 _19900_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_182_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15023_ _15023_/A vssd1 vssd1 vccd1 vccd1 _15077_/A sky130_fd_sc_hd__clkbuf_1
X_12235_ _16066_/C vssd1 vssd1 vccd1 vccd1 _16408_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21797__B1 _22365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19831_ _19831_/A _19831_/B _19831_/C vssd1 vssd1 vccd1 vccd1 _19831_/X sky130_fd_sc_hd__and3_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12166_ _12166_/A _12166_/B vssd1 vssd1 vccd1 vccd1 _12181_/A sky130_fd_sc_hd__nand2_1
XFILLER_123_686 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19762_ _19762_/A _19762_/B vssd1 vssd1 vccd1 vccd1 _19771_/C sky130_fd_sc_hd__nand2_2
XFILLER_110_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12097_ _23385_/Q _23384_/Q _23382_/Q _23383_/Q vssd1 vssd1 vccd1 vccd1 _18649_/A
+ sky130_fd_sc_hd__nor4_4
X_16974_ _16740_/A _16784_/Y _16733_/A vssd1 vssd1 vccd1 vccd1 _16975_/B sky130_fd_sc_hd__a21bo_1
X_18713_ _18721_/B vssd1 vssd1 vccd1 vccd1 _18715_/A sky130_fd_sc_hd__inv_2
XFILLER_77_762 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15925_ _11871_/A _15774_/A _16194_/C vssd1 vssd1 vccd1 vccd1 _15925_/Y sky130_fd_sc_hd__o21ai_2
X_19693_ _19483_/Y _19692_/Y _19521_/B _19521_/C vssd1 vssd1 vccd1 vccd1 _19719_/A
+ sky130_fd_sc_hd__a22o_1
Xinput8 wb_dat_i[10] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_4
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12949__A _20905_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14867__C _14867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18644_ _19859_/A _18453_/X _20146_/B _18804_/A _17134_/B vssd1 vssd1 vccd1 vccd1
+ _18647_/B sky130_fd_sc_hd__o2111ai_4
X_15856_ _15630_/Y _15645_/A _15672_/C vssd1 vssd1 vccd1 vccd1 _15856_/Y sky130_fd_sc_hd__a21oi_4
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17243__C _19674_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14807_ _14167_/A _15019_/A _14819_/A _14806_/X vssd1 vssd1 vccd1 vccd1 _14928_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_80_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18575_ _18568_/B _18568_/C _18568_/A vssd1 vssd1 vccd1 vccd1 _18576_/B sky130_fd_sc_hd__a21oi_1
X_15787_ _15773_/Y _15775_/X _15786_/Y vssd1 vssd1 vccd1 vccd1 _15787_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _12633_/A _21061_/A _13029_/A vssd1 vssd1 vccd1 vccd1 _12999_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17526_ _17934_/B vssd1 vssd1 vccd1 vccd1 _17527_/C sky130_fd_sc_hd__clkbuf_2
X_14738_ _14738_/A vssd1 vssd1 vccd1 vccd1 _14738_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17457_ _17285_/A _17600_/A _17260_/B vssd1 vssd1 vccd1 vccd1 _17457_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_177_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14669_ _23336_/Q _14668_/X _14642_/X _23304_/Q _14657_/X vssd1 vssd1 vccd1 vccd1
+ _14669_/X sky130_fd_sc_hd__a221o_1
XANTENNA__16156__A _19363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16408_ _16408_/A vssd1 vssd1 vccd1 vccd1 _16408_/X sky130_fd_sc_hd__buf_2
XFILLER_193_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17388_ _17388_/A _19675_/C _19512_/D _17898_/D vssd1 vssd1 vccd1 vccd1 _17549_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_119_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19142__A1 _18944_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19127_ _19118_/Y _19119_/Y _19126_/X _19121_/X vssd1 vssd1 vccd1 vccd1 _19127_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16339_ _16340_/B _16296_/Y _16338_/Y vssd1 vssd1 vccd1 vccd1 _16339_/X sky130_fd_sc_hd__o21a_1
XFILLER_158_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17153__B1 _17161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23542__CLK _23582_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19058_ _19058_/A _19058_/B vssd1 vssd1 vccd1 vccd1 _19060_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11605__B1_N _11604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18009_ _18004_/X _18005_/X _18006_/X _18008_/X vssd1 vssd1 vccd1 vccd1 _18114_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_133_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21020_ _21012_/X _21006_/Y _21015_/X vssd1 vssd1 vccd1 vccd1 _21020_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15219__B _15219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22971_ _21832_/A input7/X _22979_/S vssd1 vssd1 vccd1 vccd1 _22972_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13493__A2 _13732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14777__C _14777_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21922_ _21922_/A _21922_/B vssd1 vssd1 vccd1 vccd1 _21922_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21853_ _21853_/A _23482_/Q vssd1 vssd1 vccd1 vccd1 _21854_/B sky130_fd_sc_hd__and2_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13245__A2 _22476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12297__C _12297_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17450__A _19534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20804_ _12877_/Y _20814_/A _20973_/A vssd1 vssd1 vccd1 vccd1 _20805_/A sky130_fd_sc_hd__o21ai_1
XFILLER_169_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21784_ _21755_/A _21760_/A _21783_/X vssd1 vssd1 vccd1 vccd1 _21875_/A sky130_fd_sc_hd__a21o_1
XFILLER_24_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_342 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23523_ _23575_/CLK _23523_/D vssd1 vssd1 vccd1 vccd1 _23523_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20735_ _20853_/A _20854_/A _20853_/B vssd1 vssd1 vccd1 vccd1 _20737_/B sky130_fd_sc_hd__nand3_1
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16066__A _16066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14745__A2 _16815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23454_ _23571_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 _23454_/Q sky130_fd_sc_hd__dfxtp_2
X_20666_ _20666_/A _20666_/B vssd1 vssd1 vccd1 vccd1 _20667_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22405_ _22405_/A _22405_/B _22405_/C vssd1 vssd1 vccd1 vccd1 _22406_/B sky130_fd_sc_hd__nand3_1
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20597_ _20597_/A _20597_/B _20597_/C vssd1 vssd1 vccd1 vccd1 _20605_/A sky130_fd_sc_hd__nand3_4
X_23385_ _23385_/CLK _23385_/D vssd1 vssd1 vccd1 vccd1 _23385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23217__A0 _23428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22336_ _22716_/D vssd1 vssd1 vccd1 vccd1 _22756_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_152_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17695__B2 _23525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14902__C1 _14980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22267_ _22267_/A vssd1 vssd1 vccd1 vccd1 _22566_/A sky130_fd_sc_hd__clkbuf_2
X_12020_ _15905_/A vssd1 vssd1 vccd1 vccd1 _12020_/X sky130_fd_sc_hd__buf_2
XFILLER_183_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21218_ _21319_/A _21218_/B _21218_/C vssd1 vssd1 vccd1 vccd1 _21218_/X sky130_fd_sc_hd__and3_1
XANTENNA__18644__B1 _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22198_ _22166_/A _22166_/B _22166_/C _22176_/A vssd1 vssd1 vccd1 vccd1 _22199_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_160_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17625__A _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21149_ _21125_/A _21125_/B _21134_/B _21236_/A vssd1 vssd1 vccd1 vccd1 _21149_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_24_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19543__C _19811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13971_ _13890_/A _13890_/B _15084_/A vssd1 vssd1 vccd1 vccd1 _13971_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12769__A _23452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15710_ _15908_/A _15908_/B _15721_/A vssd1 vssd1 vccd1 vccd1 _15719_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__19840__A _19840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12922_ _13138_/C _13138_/D _12923_/C vssd1 vssd1 vccd1 vccd1 _12962_/A sky130_fd_sc_hd__a21o_1
XFILLER_74_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16690_ _16360_/A _15655_/X _15902_/B _16202_/Y vssd1 vssd1 vccd1 vccd1 _16690_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15641_ _11871_/A _15797_/A _15640_/Y vssd1 vssd1 vccd1 vccd1 _15641_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_92_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12853_ _12633_/A _12862_/A _12851_/Y _12648_/A _12852_/Y vssd1 vssd1 vccd1 vccd1
+ _12859_/B sky130_fd_sc_hd__o221ai_2
XFILLER_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19357__D1 _17581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _18403_/A _18403_/B _23535_/Q vssd1 vssd1 vccd1 vccd1 _18370_/B sky130_fd_sc_hd__and3_1
X_11804_ _11799_/X _11801_/X _19123_/C _11788_/Y _11803_/X vssd1 vssd1 vccd1 vccd1
+ _11805_/C sky130_fd_sc_hd__o2111ai_2
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15572_ _15577_/A _23508_/Q _15569_/B vssd1 vssd1 vccd1 vccd1 _15573_/B sky130_fd_sc_hd__o21ai_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12784_/A vssd1 vssd1 vccd1 vccd1 _12815_/B sky130_fd_sc_hd__buf_2
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19372__A1 _12243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17311_ _17140_/B _17305_/Y _17888_/A _17307_/Y _16529_/C vssd1 vssd1 vccd1 vccd1
+ _17313_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__23512__D input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14523_ input3/X vssd1 vssd1 vccd1 vccd1 _14538_/C sky130_fd_sc_hd__clkbuf_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _18322_/A _18349_/A _18349_/B vssd1 vssd1 vccd1 vccd1 _18292_/B sky130_fd_sc_hd__o21ai_1
XFILLER_15_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _16364_/A _16364_/B vssd1 vssd1 vccd1 vccd1 _11736_/A sky130_fd_sc_hd__nand2_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17242_ _19334_/A vssd1 vssd1 vccd1 vccd1 _19674_/B sky130_fd_sc_hd__clkbuf_4
X_14454_ _14441_/Y _14445_/Y _14453_/Y vssd1 vssd1 vccd1 vccd1 _14454_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_186_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11666_ _11980_/A _11980_/B _11983_/A _11665_/Y vssd1 vssd1 vccd1 vccd1 _12024_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13405_ _21793_/C _22035_/C _21793_/B vssd1 vssd1 vccd1 vccd1 _13446_/B sky130_fd_sc_hd__and3_1
X_17173_ _17173_/A _17173_/B vssd1 vssd1 vccd1 vccd1 _17181_/A sky130_fd_sc_hd__nand2_1
X_14385_ _14149_/A _14751_/B _14246_/A _14458_/A vssd1 vssd1 vccd1 vccd1 _14385_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_128_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11597_ _23382_/Q vssd1 vssd1 vccd1 vccd1 _11618_/C sky130_fd_sc_hd__buf_2
XFILLER_183_862 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16124_ _11971_/X _11972_/X _15821_/A _16047_/A vssd1 vssd1 vccd1 vccd1 _16124_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_128_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13336_ _13377_/C vssd1 vssd1 vccd1 vccd1 _13354_/B sky130_fd_sc_hd__buf_2
XFILLER_170_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16423__B _16423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_574 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15697__B1 _14569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16055_ _16055_/A vssd1 vssd1 vccd1 vccd1 _16055_/X sky130_fd_sc_hd__buf_2
X_13267_ _13495_/A _13279_/A vssd1 vssd1 vccd1 vccd1 _13268_/C sky130_fd_sc_hd__nor2_1
XFILLER_170_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15006_ _15124_/A _15124_/B _15013_/C _15013_/D vssd1 vssd1 vccd1 vccd1 _15006_/Y
+ sky130_fd_sc_hd__nand4_1
X_12218_ _12159_/X _12160_/Y _12162_/Y vssd1 vssd1 vccd1 vccd1 _12218_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_155_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15039__B _15075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13198_ _13175_/X _13195_/X _13196_/Y _13197_/X vssd1 vssd1 vccd1 vccd1 _13199_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12380__C1 _19082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19814_ _20061_/A _20055_/C _20055_/D vssd1 vssd1 vccd1 vccd1 _19815_/B sky130_fd_sc_hd__and3_1
XANTENNA__17535__A _17535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12149_ _12149_/A vssd1 vssd1 vccd1 vccd1 _12149_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_2_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__23256__B _23256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19745_ _19733_/Y _19743_/X _19744_/X vssd1 vssd1 vccd1 vccd1 _19745_/Y sky130_fd_sc_hd__a21boi_2
X_16957_ _16957_/A _16957_/B vssd1 vssd1 vccd1 vccd1 _16961_/C sky130_fd_sc_hd__nand2_2
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15055__A _15353_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15908_ _15908_/A _15908_/B vssd1 vssd1 vccd1 vccd1 _15908_/Y sky130_fd_sc_hd__nor2_1
X_19676_ _19859_/A _19674_/Y _19675_/X _19667_/A vssd1 vssd1 vccd1 vccd1 _19676_/X
+ sky130_fd_sc_hd__o211a_1
X_16888_ _16888_/A _16888_/B _16888_/C vssd1 vssd1 vccd1 vccd1 _16953_/A sky130_fd_sc_hd__nand3_2
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16413__A2 _17406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18627_ _18464_/B _18464_/C _18464_/A vssd1 vssd1 vccd1 vccd1 _18627_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15839_ _16022_/A _15894_/A _15895_/A vssd1 vssd1 vccd1 vccd1 _16078_/A sky130_fd_sc_hd__a21o_1
XFILLER_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19900__D _19900_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21092__B1_N _20984_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18558_ _12540_/A _12540_/B _18565_/A vssd1 vssd1 vccd1 vccd1 _18564_/B sky130_fd_sc_hd__a21boi_1
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17509_ _16480_/X _12379_/X _18376_/B _18376_/D _17361_/B vssd1 vssd1 vccd1 vccd1
+ _17514_/D sky130_fd_sc_hd__o41ai_2
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18489_ _18473_/X _18480_/Y _18481_/X vssd1 vssd1 vccd1 vccd1 _18670_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__17420__D _17860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21170__B2 _12674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12845__C _12845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20520_ _20509_/A _20509_/B _20506_/X vssd1 vssd1 vccd1 vccd1 _20520_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_166_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15924__A1 _11864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19115__A1 _19116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20451_ _20455_/A _20451_/B _20451_/C vssd1 vssd1 vccd1 vccd1 _20457_/A sky130_fd_sc_hd__nor3_1
XFILLER_159_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20382_ _20327_/A _20329_/B _20331_/B _20331_/A _20381_/A vssd1 vssd1 vccd1 vccd1
+ _20383_/B sky130_fd_sc_hd__o221ai_2
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23170_ _23407_/Q input24/X _23178_/S vssd1 vssd1 vccd1 vccd1 _23171_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22121_ _22121_/A vssd1 vssd1 vccd1 vccd1 _22644_/A sky130_fd_sc_hd__buf_2
XFILLER_134_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15152__A2 _14184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22052_ _22025_/Y _22032_/Y _22051_/X vssd1 vssd1 vccd1 vccd1 _22052_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_161_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21003_ _21130_/A _21001_/Y _21002_/Y vssd1 vssd1 vccd1 vccd1 _21003_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17445__A _17445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19363__C _19363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12269__A3 _16523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19082__D _20368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22954_ _23311_/Q input24/X _22962_/S vssd1 vssd1 vccd1 vccd1 _22955_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21905_ _21905_/A _21905_/B _22031_/A vssd1 vssd1 vccd1 vccd1 _22037_/A sky130_fd_sc_hd__nand3_2
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22885_ _22885_/A _22885_/B vssd1 vssd1 vccd1 vccd1 _23574_/D sky130_fd_sc_hd__nor2_4
XFILLER_44_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23588__CLK _23588_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21836_ _21844_/B vssd1 vssd1 vccd1 vccd1 _21836_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16508__B _16558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21767_ _21767_/A vssd1 vssd1 vccd1 vccd1 _22508_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23506_ _23510_/CLK hold23/X vssd1 vssd1 vccd1 vccd1 _23506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20718_ _20718_/A _20718_/B vssd1 vssd1 vccd1 vccd1 _20718_/Y sky130_fd_sc_hd__nand2_1
X_21698_ _21698_/A _21698_/B _21698_/C _21704_/D vssd1 vssd1 vccd1 vccd1 _21716_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_134_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12729__A1 _12709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21430__A _21432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23437_ _23437_/CLK _23437_/D vssd1 vssd1 vccd1 vccd1 _23437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20649_ _20962_/A _20801_/C _20962_/C vssd1 vssd1 vccd1 vccd1 _20649_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__19657__A2 _19307_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14170_ _14818_/B _14821_/A _14818_/A vssd1 vssd1 vccd1 vccd1 _14227_/B sky130_fd_sc_hd__a21oi_2
XFILLER_137_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23368_ _23433_/CLK _23368_/D vssd1 vssd1 vccd1 vccd1 _23368_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__20046__A _20046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11668__A _19363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__A2 _11951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ _13121_/A _13121_/B _13121_/C _20905_/C vssd1 vssd1 vccd1 vccd1 _13124_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_180_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22319_ _22197_/A _22197_/B _22290_/A _22318_/Y vssd1 vssd1 vccd1 vccd1 _22319_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_178_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23299_ _23300_/CLK _23299_/D vssd1 vssd1 vccd1 vccd1 _23299_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18617__B1 _11915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_718 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ _13052_/A _23453_/Q _13052_/C vssd1 vssd1 vccd1 vccd1 _13058_/B sky130_fd_sc_hd__nand3_1
XFILLER_127_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12003_ _11625_/A _11711_/B _11916_/A _11647_/B vssd1 vssd1 vccd1 vccd1 _16032_/A
+ sky130_fd_sc_hd__a211oi_4
X_17860_ _17860_/A _20142_/A vssd1 vssd1 vccd1 vccd1 _17860_/Y sky130_fd_sc_hd__nand2_2
XFILLER_120_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23507__D input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16811_ _15742_/X _15766_/X _17742_/A _17741_/A _17055_/A vssd1 vssd1 vccd1 vccd1
+ _16811_/X sky130_fd_sc_hd__o221a_1
X_17791_ _17791_/A vssd1 vssd1 vccd1 vccd1 _17798_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12499__A _16141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1024 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19530_ _19530_/A _19694_/A _19799_/C _19530_/D vssd1 vssd1 vccd1 vccd1 _19534_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16742_ _16742_/A vssd1 vssd1 vccd1 vccd1 _18276_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13954_ _14058_/A _13943_/X _13953_/Y vssd1 vssd1 vccd1 vccd1 _13954_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__15306__C _15415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12905_ _12901_/A _12901_/B _12901_/C _12901_/D vssd1 vssd1 vccd1 vccd1 _12905_/Y
+ sky130_fd_sc_hd__a22oi_4
X_19461_ _19461_/A vssd1 vssd1 vccd1 vccd1 _19636_/A sky130_fd_sc_hd__inv_2
X_16673_ _16662_/A _16662_/B _17388_/A _16318_/C _16704_/B vssd1 vssd1 vccd1 vccd1
+ _16939_/B sky130_fd_sc_hd__o2111ai_2
X_13885_ _23365_/Q vssd1 vssd1 vccd1 vccd1 _14024_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21267__A_N _21207_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18412_ _18277_/D _20317_/C _20317_/B _18376_/C _18376_/D vssd1 vssd1 vccd1 vccd1
+ _18413_/B sky130_fd_sc_hd__a311o_1
XFILLER_59_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12836_ _12836_/A _12836_/B vssd1 vssd1 vccd1 vccd1 _12837_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15624_ _15624_/A vssd1 vssd1 vccd1 vccd1 _15637_/D sky130_fd_sc_hd__buf_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _19392_/A vssd1 vssd1 vccd1 vccd1 _19601_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18343_ _18384_/B _18343_/B vssd1 vssd1 vccd1 vccd1 _18344_/B sky130_fd_sc_hd__and2b_1
XANTENNA__22139__C _22139_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15555_ _15540_/A _15539_/A _15539_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _15564_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12770_/B _12770_/C _13122_/B _12766_/X vssd1 vssd1 vccd1 vccd1 _12845_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_790 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14506_ _16821_/A vssd1 vssd1 vccd1 vccd1 _15964_/B sky130_fd_sc_hd__clkbuf_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18274_ _18330_/A _20265_/A _18328_/A _18276_/C vssd1 vssd1 vccd1 vccd1 _18274_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11718_ _12323_/A _11670_/X _11682_/Y _12297_/A vssd1 vssd1 vccd1 vccd1 _11908_/A
+ sky130_fd_sc_hd__o31a_2
XANTENNA__16137__C _16308_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15486_ _15486_/A vssd1 vssd1 vccd1 vccd1 _15486_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15906__A1 _16054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15906__B2 _15621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12698_ _20645_/C vssd1 vssd1 vccd1 vccd1 _20663_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_159_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17225_ _18506_/A vssd1 vssd1 vccd1 vccd1 _19664_/B sky130_fd_sc_hd__buf_4
X_14437_ _14465_/A _14435_/X _14465_/B vssd1 vssd1 vccd1 vccd1 _14446_/A sky130_fd_sc_hd__a21boi_1
XFILLER_30_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput11 wb_dat_i[13] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_4
X_11649_ _11809_/A vssd1 vssd1 vccd1 vccd1 _11649_/X sky130_fd_sc_hd__buf_2
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 wb_dat_i[23] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__22101__B1 _22102_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput33 wb_dat_i[4] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_4
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17156_ _17156_/A _17156_/B vssd1 vssd1 vccd1 vccd1 _17161_/B sky130_fd_sc_hd__nor2_1
Xinput44 x[1] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_2
XFILLER_128_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14368_ _14365_/C _14368_/B _14368_/C vssd1 vssd1 vccd1 vccd1 _14422_/C sky130_fd_sc_hd__nand3b_1
XFILLER_196_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16107_ _15650_/Y _15772_/X _15641_/Y vssd1 vssd1 vccd1 vccd1 _16276_/A sky130_fd_sc_hd__a21boi_4
XFILLER_157_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11943__A2 _15882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11578__A _23589_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13319_ _13279_/A _13491_/A _13630_/A vssd1 vssd1 vccd1 vccd1 _13320_/A sky130_fd_sc_hd__o21ai_1
XFILLER_182_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17087_ _19123_/B vssd1 vssd1 vccd1 vccd1 _20049_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14299_ _14936_/B vssd1 vssd1 vccd1 vccd1 _15075_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_143_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16038_ _16300_/A _16038_/B vssd1 vssd1 vccd1 vccd1 _16039_/A sky130_fd_sc_hd__nand2_1
XFILLER_192_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18623__A3 _18778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_1_0_bq_clk_i clkbuf_4_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _23499_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17989_ _17962_/X _17970_/Y _17984_/Y _17988_/Y vssd1 vssd1 vccd1 vccd1 _17999_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__21218__C _21218_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14645__A1 _23396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14645__B2 _23428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19728_ _19555_/Y _19556_/X _19546_/Y vssd1 vssd1 vccd1 vccd1 _19728_/X sky130_fd_sc_hd__o21a_1
XANTENNA__19480__A _19480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21915__B1 _22269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13999__A3 _14331_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19659_ _20046_/A _20047_/A _19659_/C vssd1 vssd1 vccd1 vccd1 _19659_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__17712__B _17712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18096__A _18096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22670_ _22670_/A _22725_/A _22670_/C _22670_/D vssd1 vssd1 vccd1 vccd1 _22671_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19336__A1 _18993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12959__A1 _21276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21621_ _21577_/B _21611_/B _21608_/Y _21568_/A vssd1 vssd1 vccd1 vccd1 _21621_/Y
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__11760__B _11760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18824__A _19011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21552_ _21552_/A _21633_/A vssd1 vssd1 vccd1 vccd1 _21556_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20503_ _12748_/X _20479_/A _12875_/C vssd1 vssd1 vccd1 vccd1 _20504_/A sky130_fd_sc_hd__o21a_1
XFILLER_193_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21483_ _21484_/C _21484_/A _23568_/Q vssd1 vssd1 vccd1 vccd1 _21485_/A sky130_fd_sc_hd__a21o_1
XFILLER_14_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23222_ _23430_/Q input14/X _23228_/S vssd1 vssd1 vccd1 vccd1 _23223_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13384__A1 _13304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20434_ _20414_/B _20414_/A _20205_/X _20120_/X vssd1 vssd1 vccd1 vccd1 _20446_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13687__B _22663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11934__A2 _11926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23153_ _23153_/A vssd1 vssd1 vccd1 vccd1 _23399_/D sky130_fd_sc_hd__clkbuf_1
X_20365_ _20365_/A vssd1 vssd1 vccd1 vccd1 _20368_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22104_ _22117_/D _22106_/B _22101_/Y _22103_/Y vssd1 vssd1 vccd1 vccd1 _22348_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_164_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20296_ _20183_/B _20183_/A _20243_/Y _20247_/B vssd1 vssd1 vccd1 vccd1 _20296_/Y
+ sky130_fd_sc_hd__o211ai_1
X_23084_ _23369_/Q input17/X _23084_/S vssd1 vssd1 vccd1 vccd1 _23085_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22035_ _22391_/A _22392_/B _22035_/C vssd1 vssd1 vccd1 vccd1 _22035_/X sky130_fd_sc_hd__and3_1
XFILLER_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16510__C _16510_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12111__A2 _12110_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22937_ _22937_/A vssd1 vssd1 vccd1 vccd1 _23303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ _13674_/A _13672_/C vssd1 vssd1 vccd1 vccd1 _13671_/C sky130_fd_sc_hd__xnor2_2
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22868_ _22868_/A _22868_/B vssd1 vssd1 vccd1 vccd1 _22868_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_71_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12621_ _12667_/B _12788_/B _12915_/A _13019_/B _20894_/A vssd1 vssd1 vccd1 vccd1
+ _12687_/A sky130_fd_sc_hd__o311ai_2
XFILLER_169_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21819_ _21817_/Y _21819_/B vssd1 vssd1 vccd1 vccd1 _21820_/B sky130_fd_sc_hd__and2b_1
XFILLER_19_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22799_ _22829_/A vssd1 vssd1 vccd1 vccd1 _22799_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15340_ _15402_/B _15402_/A vssd1 vssd1 vccd1 vccd1 _15442_/B sky130_fd_sc_hd__nor2_1
XFILLER_157_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17889__A1 _16665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12552_ _12227_/C _12080_/B _18565_/A _12540_/A vssd1 vssd1 vccd1 vccd1 _12552_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_185_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14981__B _15353_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15271_ _15271_/A _15326_/B vssd1 vssd1 vccd1 vccd1 _15271_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_968 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12483_ _12483_/A vssd1 vssd1 vccd1 vccd1 _12483_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12782__A _23453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17010_ _17010_/A _17010_/B _17010_/C _17026_/D vssd1 vssd1 vccd1 vccd1 _17012_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_172_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14222_ _14222_/A _14222_/B vssd1 vssd1 vccd1 vccd1 _14222_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18838__B1 _19029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14153_ _14150_/Y _14151_/Y _13997_/Y vssd1 vssd1 vccd1 vccd1 _14153_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_164_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13104_ _20464_/D _20464_/A _13103_/Y vssd1 vssd1 vccd1 vccd1 _13201_/A sky130_fd_sc_hd__a21oi_1
XFILLER_140_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18961_ _18951_/Y _18956_/X _18964_/A vssd1 vssd1 vccd1 vccd1 _18969_/C sky130_fd_sc_hd__o21bai_1
X_14084_ _15253_/A _14252_/D _15253_/C _14163_/B vssd1 vssd1 vccd1 vccd1 _14084_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_770 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ _17916_/A _17916_/B _17916_/C vssd1 vssd1 vccd1 vccd1 _17912_/X sky130_fd_sc_hd__and3_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13035_ _13122_/B _12936_/X _13041_/A vssd1 vssd1 vccd1 vccd1 _13035_/X sky130_fd_sc_hd__o21a_1
XFILLER_152_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18892_ _18892_/A _18892_/B vssd1 vssd1 vccd1 vccd1 _18893_/C sky130_fd_sc_hd__nand2_2
XFILLER_117_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16616__A2 _16370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1055 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17843_ _16804_/A _16804_/B _16819_/X _17050_/A vssd1 vssd1 vccd1 vccd1 _17972_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_121_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1099 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17774_ _17768_/Y _17773_/Y _17771_/Y vssd1 vssd1 vccd1 vccd1 _17782_/C sky130_fd_sc_hd__a21o_1
X_14986_ _15082_/B vssd1 vssd1 vccd1 vccd1 _15262_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19513_ _16437_/X _19858_/A _19656_/A vssd1 vssd1 vccd1 vccd1 _19514_/C sky130_fd_sc_hd__o21ai_1
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16725_ _16725_/A vssd1 vssd1 vccd1 vccd1 _16725_/Y sky130_fd_sc_hd__inv_2
X_13937_ _14044_/B vssd1 vssd1 vccd1 vccd1 _13937_/X sky130_fd_sc_hd__buf_2
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17577__B1 _20133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21373__A1 _20957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13850__A2 _21987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19444_ _19427_/X _19433_/Y _19439_/Y _19275_/Y vssd1 vssd1 vccd1 vccd1 _19444_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__21054__B _21054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16656_ _16723_/A _16723_/B _16723_/C vssd1 vssd1 vccd1 vccd1 _16950_/A sky130_fd_sc_hd__nand3_2
X_13868_ _21856_/A _21856_/B vssd1 vssd1 vccd1 vccd1 _13870_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12819_ _12975_/A _12819_/B vssd1 vssd1 vccd1 vccd1 _12908_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15607_ _23429_/Q vssd1 vssd1 vccd1 vccd1 _15729_/A sky130_fd_sc_hd__inv_2
X_19375_ _19568_/A _19569_/A vssd1 vssd1 vccd1 vccd1 _19387_/A sky130_fd_sc_hd__nand2_1
X_13799_ _13799_/A vssd1 vssd1 vccd1 vccd1 _13799_/X sky130_fd_sc_hd__clkbuf_2
X_16587_ _16586_/Y _16266_/C _16275_/A vssd1 vssd1 vccd1 vccd1 _16587_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18326_ _20368_/A vssd1 vssd1 vccd1 vccd1 _20366_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15538_ _15538_/A _15538_/B _15538_/C _15538_/D vssd1 vssd1 vccd1 vccd1 _15539_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16001__B1 _15878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18257_ _18254_/Y _18417_/D _18302_/B vssd1 vssd1 vccd1 vccd1 _18364_/B sky130_fd_sc_hd__a21o_1
XFILLER_148_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15469_ _15468_/X _15413_/B _15409_/A _15412_/B vssd1 vssd1 vccd1 vccd1 _15471_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__16552__A1 _16054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17208_ _17524_/C _17524_/D vssd1 vssd1 vccd1 vccd1 _17208_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18188_ _18242_/B _18242_/A vssd1 vssd1 vccd1 vccd1 _18209_/A sky130_fd_sc_hd__xnor2_1
XFILLER_155_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16314__D _17133_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17139_ _12004_/X _12006_/X _15936_/A _15937_/A vssd1 vssd1 vccd1 vccd1 _17140_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16304__B2 _16447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20150_ _20135_/X _20136_/X _20158_/A _20158_/B vssd1 vssd1 vccd1 vccd1 _20150_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__16855__A2 _11921_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14866__A1 _14879_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20081_ _20081_/A _20081_/B _20365_/A _20081_/D vssd1 vssd1 vccd1 vccd1 _20083_/A
+ sky130_fd_sc_hd__or4_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20133__B _20133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14618__A1 _14614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14618__B2 _14615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17723__A _17723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19557__A1 _12053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19557__B2 _17600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17568__B1 _16056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20983_ _20843_/B _20842_/A _20842_/B vssd1 vssd1 vccd1 vccd1 _20987_/B sky130_fd_sc_hd__a21bo_1
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22722_ _22722_/A _22722_/B _22722_/C vssd1 vssd1 vccd1 vccd1 _22723_/B sky130_fd_sc_hd__and3_1
XFILLER_26_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15043__A1 _15208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22653_ _13547_/X _22461_/X _22703_/A _22650_/B vssd1 vssd1 vccd1 vccd1 _22712_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__21116__A1 _21159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21604_ _21564_/A _21564_/B _21564_/C vssd1 vssd1 vccd1 vccd1 _21605_/C sky130_fd_sc_hd__a21boi_1
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22584_ _22556_/X _22584_/B _22584_/C vssd1 vssd1 vccd1 vccd1 _22589_/B sky130_fd_sc_hd__nand3b_1
XFILLER_167_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20875__B1 _21542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21535_ _21418_/B _21418_/C _21418_/A vssd1 vssd1 vccd1 vccd1 _21535_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16543__A1 _16530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14554__B1 _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21466_ _21465_/A _21465_/B _21465_/C vssd1 vssd1 vccd1 vccd1 _21467_/B sky130_fd_sc_hd__a21o_1
XFILLER_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23205_ _23205_/A vssd1 vssd1 vccd1 vccd1 _23422_/D sky130_fd_sc_hd__clkbuf_1
X_20417_ _20452_/C _20417_/B vssd1 vssd1 vccd1 vccd1 _20419_/B sky130_fd_sc_hd__nand2_1
XFILLER_135_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21397_ _21397_/A _21397_/B vssd1 vssd1 vccd1 vccd1 _21399_/C sky130_fd_sc_hd__and2_1
XANTENNA__16802__A _16802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23136_ _23182_/S vssd1 vssd1 vccd1 vccd1 _23145_/S sky130_fd_sc_hd__clkbuf_2
X_20348_ _20343_/Y _20344_/X _20384_/B _20340_/Y _20341_/X vssd1 vssd1 vccd1 vccd1
+ _20356_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_190_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23067_ _14879_/C input9/X _23073_/S vssd1 vssd1 vccd1 vccd1 _23068_/A sky130_fd_sc_hd__mux2_1
X_20279_ _20328_/A _20328_/B _20328_/C vssd1 vssd1 vccd1 vccd1 _20279_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16059__B1 _16464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22018_ _22018_/A _23330_/Q vssd1 vssd1 vccd1 vccd1 _22144_/C sky130_fd_sc_hd__nand2_4
XFILLER_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14609__A1 _15605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17633__A _17723_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_348 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14840_ _14836_/Y _14840_/B _14840_/C vssd1 vssd1 vccd1 vccd1 _14844_/B sky130_fd_sc_hd__nand3b_1
XFILLER_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14085__A2 _14068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14771_ _14878_/A _14883_/A _14091_/A _23361_/Q vssd1 vssd1 vccd1 vccd1 _14774_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA_input17_A wb_dat_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11983_ _11983_/A _12282_/A _18469_/D vssd1 vssd1 vccd1 vccd1 _18812_/B sky130_fd_sc_hd__nand3_4
XFILLER_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16510_ _16539_/A _16539_/B _16510_/C _18017_/D vssd1 vssd1 vccd1 vccd1 _16532_/C
+ sky130_fd_sc_hd__nand4_1
X_13722_ _13569_/Y _13720_/Y _13575_/Y vssd1 vssd1 vccd1 vccd1 _13723_/C sky130_fd_sc_hd__a21bo_1
XFILLER_147_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17490_ _17663_/A _17663_/B _17497_/C _17497_/D vssd1 vssd1 vccd1 vccd1 _17490_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_186_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16441_ _16436_/X _16438_/Y _16440_/Y vssd1 vssd1 vccd1 vccd1 _16441_/Y sky130_fd_sc_hd__o21ai_1
X_13653_ _13645_/A _13645_/B _13651_/X _13652_/X vssd1 vssd1 vccd1 vccd1 _13653_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_108_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14388__A3 _13985_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _12571_/X _12766_/A _12652_/A vssd1 vssd1 vccd1 vccd1 _12604_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_169_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _16372_/A vssd1 vssd1 vccd1 vccd1 _16457_/D sky130_fd_sc_hd__clkbuf_2
X_19160_ _19308_/C vssd1 vssd1 vccd1 vccd1 _19651_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13584_ _13756_/A _13756_/B _13585_/A _22700_/D vssd1 vssd1 vccd1 vccd1 _13698_/B
+ sky130_fd_sc_hd__o211a_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19720__A1 _12324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18111_ _18022_/B _18028_/B _18109_/Y _18110_/X vssd1 vssd1 vccd1 vccd1 _18156_/A
+ sky130_fd_sc_hd__a211o_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _15245_/B _15315_/X _15321_/X vssd1 vssd1 vccd1 vccd1 _15323_/X sky130_fd_sc_hd__a21o_1
XFILLER_158_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _18557_/B _12523_/B _12528_/A _12528_/B vssd1 vssd1 vccd1 vccd1 _12535_/Y
+ sky130_fd_sc_hd__o211ai_2
X_19091_ _19091_/A _19091_/B _19091_/C vssd1 vssd1 vccd1 vccd1 _19091_/Y sky130_fd_sc_hd__nand3_1
XFILLER_9_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18042_ _18043_/C _18043_/B _18043_/A vssd1 vssd1 vccd1 vccd1 _18132_/A sky130_fd_sc_hd__a21oi_1
XFILLER_172_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15254_ _15254_/A _15254_/B _15254_/C vssd1 vssd1 vccd1 vccd1 _15255_/B sky130_fd_sc_hd__nand3_1
X_12466_ _12461_/Y _12463_/Y _12465_/X vssd1 vssd1 vccd1 vccd1 _12469_/B sky130_fd_sc_hd__a21o_1
XFILLER_166_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14205_ _14934_/A _14800_/B _14800_/A vssd1 vssd1 vccd1 vccd1 _14219_/C sky130_fd_sc_hd__a21o_1
X_15185_ _15185_/A _15185_/B _15185_/C vssd1 vssd1 vccd1 vccd1 _15190_/A sky130_fd_sc_hd__nand3_1
X_12397_ _12396_/A _12396_/B _12396_/C vssd1 vssd1 vccd1 vccd1 _12546_/A sky130_fd_sc_hd__a21o_1
XFILLER_193_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16298__B1 _15862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14136_ _14181_/A _14115_/Y _14116_/X _14118_/X _14121_/Y vssd1 vssd1 vccd1 vccd1
+ _14137_/C sky130_fd_sc_hd__o221ai_1
XANTENNA_output85_A _14603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19993_ _19822_/A _19823_/A _19992_/X vssd1 vssd1 vccd1 vccd1 _19993_/X sky130_fd_sc_hd__a21o_1
XFILLER_152_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18944_ _18944_/A _18944_/B _18944_/C vssd1 vssd1 vccd1 vccd1 _18944_/Y sky130_fd_sc_hd__nand3_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23032__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ _14777_/B vssd1 vssd1 vccd1 vccd1 _14980_/A sky130_fd_sc_hd__clkbuf_2
X_13018_ _20628_/B _23447_/Q vssd1 vssd1 vccd1 vccd1 _13018_/Y sky130_fd_sc_hd__nand2_2
XFILLER_95_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18875_ _18875_/A _18875_/B _18875_/C vssd1 vssd1 vccd1 vccd1 _18875_/X sky130_fd_sc_hd__and3_1
XFILLER_94_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_955 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17826_ _17935_/D _17703_/B _17703_/C _17943_/A _18253_/A vssd1 vssd1 vccd1 vccd1
+ _17828_/A sky130_fd_sc_hd__a311o_1
XFILLER_95_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13790__B _22064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21065__A _21065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17757_ _17710_/X _17760_/B _17754_/Y _17969_/D _20217_/D vssd1 vssd1 vccd1 vccd1
+ _17773_/D sky130_fd_sc_hd__o2111ai_2
XFILLER_81_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14969_ _23361_/Q _14864_/Y _14970_/B vssd1 vssd1 vccd1 vccd1 _15115_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__19180__D _19180_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16708_ _16708_/A _16708_/B vssd1 vssd1 vccd1 vccd1 _16709_/C sky130_fd_sc_hd__nand2_1
XFILLER_35_543 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17688_ _23527_/Q vssd1 vssd1 vccd1 vccd1 _17693_/A sky130_fd_sc_hd__inv_2
XFILLER_62_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19427_ _19428_/A _19616_/A _19427_/C vssd1 vssd1 vccd1 vccd1 _19427_/X sky130_fd_sc_hd__and3_1
XANTENNA__15998__A _15998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16639_ _16639_/A vssd1 vssd1 vccd1 vccd1 _16639_/X sky130_fd_sc_hd__buf_2
XANTENNA__18374__A _20368_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19358_ _17742_/X _17741_/X _12185_/X _12184_/X _17443_/A vssd1 vssd1 vccd1 vccd1
+ _19358_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15981__C1 _12207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18093__B _19967_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19711__A1 _12053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18309_ _18309_/A _18362_/A _18362_/B vssd1 vssd1 vccd1 vccd1 _18319_/C sky130_fd_sc_hd__nand3_1
XFILLER_175_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19289_ _18926_/A _19289_/B _19289_/C vssd1 vssd1 vccd1 vccd1 _19290_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__16525__B2 _17248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21320_ _21317_/Y _21318_/X _21319_/Y vssd1 vssd1 vccd1 vccd1 _21320_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12215__A2_N _12110_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21251_ _21123_/X _21129_/Y _21135_/Y _21151_/Y _21241_/A vssd1 vssd1 vccd1 vccd1
+ _21251_/Y sky130_fd_sc_hd__o2111ai_2
XFILLER_172_960 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20202_ _20310_/C _20310_/B vssd1 vssd1 vccd1 vccd1 _20203_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_515 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21182_ _21500_/A _21279_/D _21440_/C _21182_/D vssd1 vssd1 vccd1 vccd1 _21184_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_144_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11766__A _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20133_ _20268_/C _20133_/B _20212_/A _20133_/D vssd1 vssd1 vccd1 vccd1 _20134_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__23023__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20064_ _12113_/X _18660_/X _11686_/Y _11849_/C _19800_/C vssd1 vssd1 vccd1 vccd1
+ _20066_/B sky130_fd_sc_hd__o311a_2
XFILLER_135_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A wb_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1072 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17789__B1 _18163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18450__A1 _12311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20966_ _20966_/A _20966_/B _20966_/C vssd1 vssd1 vccd1 vccd1 _20967_/B sky130_fd_sc_hd__and3_1
XFILLER_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_159 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19950__A1 _16408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17410__C1 _18503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22705_ _22707_/A _22702_/X _22707_/B vssd1 vssd1 vccd1 vccd1 _22709_/A sky130_fd_sc_hd__a21oi_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _20479_/X _21047_/C _20897_/C _20897_/D vssd1 vssd1 vccd1 vccd1 _20902_/A
+ sky130_fd_sc_hd__nand4b_1
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22636_ _22637_/A _22637_/B _22636_/C vssd1 vssd1 vccd1 vccd1 _22646_/A sky130_fd_sc_hd__nand3_1
XFILLER_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18505__A2 _16604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12250__A1 _12090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22567_ _22567_/A _22567_/B vssd1 vssd1 vccd1 vccd1 _22567_/Y sky130_fd_sc_hd__nor2_2
XFILLER_127_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12320_ _11799_/X _11801_/X _12260_/Y _19534_/C _12273_/B vssd1 vssd1 vccd1 vccd1
+ _12321_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_21_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21518_ _21516_/Y _21566_/B vssd1 vssd1 vccd1 vccd1 _21521_/B sky130_fd_sc_hd__and2b_1
XFILLER_5_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22498_ _22501_/C _22501_/D _22500_/A vssd1 vssd1 vccd1 vccd1 _22499_/C sky130_fd_sc_hd__a21o_1
XFILLER_182_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12251_ _12251_/A _12251_/B vssd1 vssd1 vccd1 vccd1 _12251_/X sky130_fd_sc_hd__or2_1
XANTENNA__12002__A1 _12184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21449_ _21506_/A vssd1 vssd1 vccd1 vccd1 _21510_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12182_ _12426_/B vssd1 vssd1 vccd1 vccd1 _19539_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_162_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23119_ _11677_/X input29/X _23123_/S vssd1 vssd1 vccd1 vccd1 _23120_/A sky130_fd_sc_hd__mux2_1
XANTENNA__19843__A _19949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17066__C _17066_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16990_ _16988_/Y _16989_/Y _16777_/Y _16998_/C vssd1 vssd1 vccd1 vccd1 _16994_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_62_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13502__A1 _22280_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15941_ _15941_/A _15943_/A _15943_/B vssd1 vssd1 vccd1 vccd1 _15948_/C sky130_fd_sc_hd__and3_1
XANTENNA__13502__B2 _22381_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17244__A2 _18093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18441__A1 _18439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18660_ _12245_/X _11784_/C _11999_/B _14646_/A vssd1 vssd1 vccd1 vccd1 _18660_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _18755_/C vssd1 vssd1 vccd1 vccd1 _19700_/C sky130_fd_sc_hd__buf_2
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23515__D input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17611_ _17644_/A vssd1 vssd1 vccd1 vccd1 _17611_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14823_ _14855_/A _14855_/B vssd1 vssd1 vccd1 vccd1 _14825_/C sky130_fd_sc_hd__xor2_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _23539_/Q _18733_/A _18589_/Y _18590_/X vssd1 vssd1 vccd1 vccd1 _18593_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14463__C1 _13972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _17498_/B _17498_/C _17498_/A _17502_/C _17502_/A vssd1 vssd1 vccd1 vccd1
+ _17673_/A sky130_fd_sc_hd__a32oi_2
XFILLER_63_148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11966_ _11966_/A _11966_/B _12066_/A _19334_/A vssd1 vssd1 vccd1 vccd1 _11967_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11816__B2 _11815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14754_ _14764_/A _14764_/B _14181_/A vssd1 vssd1 vccd1 vccd1 _14754_/X sky130_fd_sc_hd__a21o_1
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17547__A3 _17391_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13705_ _13736_/A _13720_/A _13705_/C _13705_/D vssd1 vssd1 vccd1 vccd1 _13711_/B
+ sky130_fd_sc_hd__nand4_1
X_17473_ _17473_/A _17473_/B _17473_/C _17473_/D vssd1 vssd1 vccd1 vccd1 _17475_/B
+ sky130_fd_sc_hd__nand4_2
X_14685_ _23340_/Q _14668_/X _14673_/X _23308_/Q _14678_/X vssd1 vssd1 vccd1 vccd1
+ _14685_/X sky130_fd_sc_hd__a221o_1
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11897_ _12130_/A vssd1 vssd1 vccd1 vccd1 _18461_/A sky130_fd_sc_hd__clkbuf_4
X_19212_ _19221_/B _19221_/C _19221_/A vssd1 vssd1 vccd1 vccd1 _19212_/Y sky130_fd_sc_hd__a21oi_1
X_16424_ _16424_/A _16424_/B _16424_/C vssd1 vssd1 vccd1 vccd1 _16424_/Y sky130_fd_sc_hd__nand3_1
X_13636_ _21921_/C _21793_/B _21793_/C _21764_/B _22172_/C vssd1 vssd1 vccd1 vccd1
+ _13636_/X sky130_fd_sc_hd__a32o_2
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12954__B _13181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19154__C1 _19502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16609__A1_N _16123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19143_ _19135_/Y _19410_/C _19142_/Y vssd1 vssd1 vccd1 vccd1 _19147_/A sky130_fd_sc_hd__a21o_1
XFILLER_157_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16355_ _16355_/A vssd1 vssd1 vccd1 vccd1 _16356_/A sky130_fd_sc_hd__clkbuf_4
X_13567_ _13566_/Y _13482_/Y _13479_/X vssd1 vssd1 vccd1 vccd1 _13569_/B sky130_fd_sc_hd__a21bo_1
XFILLER_157_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13131__A _13131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12518_ _17456_/A vssd1 vssd1 vccd1 vccd1 _12518_/X sky130_fd_sc_hd__buf_2
XFILLER_9_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15306_ _15363_/A _15416_/A _15415_/A _15358_/A vssd1 vssd1 vccd1 vccd1 _15308_/D
+ sky130_fd_sc_hd__nand4_2
X_19074_ _19069_/Y _19071_/X _19072_/Y _19073_/Y vssd1 vssd1 vccd1 vccd1 _19075_/C
+ sky130_fd_sc_hd__o2bb2ai_2
X_16286_ _16860_/B vssd1 vssd1 vccd1 vccd1 _17108_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13498_ _13498_/A _13498_/B vssd1 vssd1 vccd1 vccd1 _13663_/C sky130_fd_sc_hd__nand2_1
XFILLER_185_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18025_ _17902_/B _17881_/Y _18024_/X vssd1 vssd1 vccd1 vccd1 _18026_/B sky130_fd_sc_hd__a21boi_1
XFILLER_172_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15237_ _15237_/A _15237_/B vssd1 vssd1 vccd1 vccd1 _15245_/A sky130_fd_sc_hd__nand2_1
X_12449_ _12444_/A _18497_/A _12447_/Y _12448_/X vssd1 vssd1 vccd1 vccd1 _12449_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__18360__C _23535_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15168_ _15233_/B vssd1 vssd1 vccd1 vccd1 _15369_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1012 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11586__A _19017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14119_ _14262_/A vssd1 vssd1 vccd1 vccd1 _14384_/A sky130_fd_sc_hd__buf_2
XANTENNA__18680__A1 _12184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15058__A _15408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19976_ _19668_/X _17763_/X _19980_/C _20058_/A vssd1 vssd1 vccd1 vccd1 _19977_/B
+ sky130_fd_sc_hd__o211ai_1
X_15099_ _15099_/A _15099_/B vssd1 vssd1 vccd1 vccd1 _15099_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20899__A _21174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18927_ _18927_/A _18927_/B vssd1 vssd1 vccd1 vccd1 _23522_/D sky130_fd_sc_hd__xor2_1
XFILLER_80_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18858_ _18858_/A _18858_/B _18858_/C vssd1 vssd1 vccd1 vccd1 _18862_/B sky130_fd_sc_hd__nand3_1
XFILLER_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17640__C1 _17898_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17809_ _17708_/Y _17805_/Y _17808_/Y vssd1 vssd1 vccd1 vccd1 _17814_/B sky130_fd_sc_hd__o21ai_2
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18789_ _15904_/A _15905_/A _18476_/A _18484_/A _18479_/A vssd1 vssd1 vccd1 vccd1
+ _18984_/A sky130_fd_sc_hd__o221ai_2
XFILLER_48_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20820_ _20820_/A _20820_/B _20820_/C vssd1 vssd1 vccd1 vccd1 _20837_/A sky130_fd_sc_hd__nand3_1
XFILLER_39_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20751_ _20751_/A _20751_/B vssd1 vssd1 vccd1 vccd1 _20751_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23470_ _23571_/CLK _23482_/Q vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_196_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20682_ _12706_/Y _20681_/Y _20506_/X vssd1 vssd1 vccd1 vccd1 _20682_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22421_ _22405_/A _22418_/X _22420_/X vssd1 vssd1 vccd1 vccd1 _22421_/X sky130_fd_sc_hd__a21o_1
XFILLER_149_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22352_ _23275_/Q _22353_/B vssd1 vssd1 vccd1 vccd1 _22354_/A sky130_fd_sc_hd__and2_1
XFILLER_164_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21303_ _21365_/A _21314_/A _21295_/Y _21293_/Y vssd1 vssd1 vccd1 vccd1 _21303_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23244__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22283_ _22283_/A vssd1 vssd1 vccd1 vccd1 _22283_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21966__B1_N _21842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21234_ _21333_/B _21229_/Y _21231_/Y _21233_/X vssd1 vssd1 vccd1 vccd1 _21402_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16071__B _16075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21165_ _21493_/C _20966_/A _20966_/B _21164_/X vssd1 vssd1 vccd1 vccd1 _21165_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_132_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_719 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20116_ _20116_/A _20116_/B vssd1 vssd1 vccd1 vccd1 _20207_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23185__A _23241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13496__B1 _13495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21096_ _21094_/X _21095_/Y _21083_/Y vssd1 vssd1 vccd1 vccd1 _21096_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12104__B _16365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15118__D _15233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20047_ _20047_/A vssd1 vssd1 vccd1 vccd1 _20215_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_100_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_487 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18974__A2 _18490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22507__B1 _22505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11820_/A vssd1 vssd1 vccd1 vccd1 _12353_/A sky130_fd_sc_hd__buf_4
XFILLER_22_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13216__A _23479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _21997_/X _22420_/B _22420_/C _21881_/Y vssd1 vssd1 vccd1 vccd1 _21998_/Y
+ sky130_fd_sc_hd__o31ai_2
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14_0_bq_clk_i clkbuf_3_7_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _23558_/CLK
+ sky130_fd_sc_hd__clkbuf_8
X_11751_ _11820_/A _16360_/A _11766_/C vssd1 vssd1 vccd1 vccd1 _12265_/B sky130_fd_sc_hd__o21ai_2
XFILLER_54_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20949_ _20810_/B _20819_/B _20819_/A vssd1 vssd1 vccd1 vccd1 _20950_/C sky130_fd_sc_hd__a21boi_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_855 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14470_ _14819_/A vssd1 vssd1 vccd1 vccd1 _14933_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11682_ _11851_/A _11852_/A _18657_/C vssd1 vssd1 vccd1 vccd1 _11682_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_42_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20049__A _20049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_78 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13421_ _13620_/A vssd1 vssd1 vccd1 vccd1 _13453_/A sky130_fd_sc_hd__buf_2
XFILLER_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22619_ _22619_/A _22619_/B vssd1 vssd1 vccd1 vccd1 _22629_/C sky130_fd_sc_hd__nand2_1
XANTENNA__19838__A _19838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_730 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23599_ input39/X vssd1 vssd1 vccd1 vccd1 _23599_/X sky130_fd_sc_hd__clkbuf_1
X_16140_ _16140_/A _16815_/C vssd1 vssd1 vccd1 vccd1 _17741_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21494__B1 _21495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _21901_/D vssd1 vssd1 vccd1 vccd1 _13354_/C sky130_fd_sc_hd__buf_2
XFILLER_155_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17162__B2 _17155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12294__A1_N _12297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12303_ _12300_/C _12303_/B _12303_/C vssd1 vssd1 vccd1 vccd1 _12303_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_6_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16071_ _16075_/B _16075_/C vssd1 vssd1 vccd1 vccd1 _16071_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13283_ _13814_/B vssd1 vssd1 vccd1 vccd1 _22280_/B sky130_fd_sc_hd__buf_2
XANTENNA__23235__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12790__A _23454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15022_ _15022_/A _15081_/B _15022_/C vssd1 vssd1 vccd1 vccd1 _15023_/A sky130_fd_sc_hd__nand3_1
X_12234_ _12546_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12563_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17077__B _17077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19830_ _19830_/A vssd1 vssd1 vccd1 vccd1 _19876_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12165_ _11814_/A _18500_/A _11996_/Y vssd1 vssd1 vccd1 vccd1 _12166_/B sky130_fd_sc_hd__o21ai_1
XFILLER_2_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16673__B1 _17388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19761_ _19554_/X _19534_/D _19532_/X vssd1 vssd1 vccd1 vccd1 _19762_/B sky130_fd_sc_hd__a21bo_1
XFILLER_123_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16973_ _16663_/X _16704_/A _16970_/Y _16972_/X vssd1 vssd1 vccd1 vccd1 _16975_/A
+ sky130_fd_sc_hd__o22ai_1
X_12096_ _12432_/A _12099_/D _12095_/Y _12121_/A vssd1 vssd1 vccd1 vccd1 _18445_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_122_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18712_ _18712_/A vssd1 vssd1 vccd1 vccd1 _18904_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15924_ _11864_/X _11865_/X _15610_/X _15918_/C _15660_/A vssd1 vssd1 vccd1 vccd1
+ _16194_/C sky130_fd_sc_hd__o221ai_4
X_19692_ _19486_/A _19486_/B _19492_/C vssd1 vssd1 vccd1 vccd1 _19692_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_77_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput9 wb_dat_i[11] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_4
XFILLER_92_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18643_ _19180_/B vssd1 vssd1 vccd1 vccd1 _20146_/B sky130_fd_sc_hd__buf_4
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _15686_/A _15686_/B _14569_/X _15931_/A vssd1 vssd1 vccd1 vccd1 _15855_/Y
+ sky130_fd_sc_hd__a211oi_4
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21046__C _23299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17243__D _17243_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14806_ _14806_/A _14911_/C _14806_/C _15254_/B vssd1 vssd1 vccd1 vccd1 _14806_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_36_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18574_ _18576_/A _18570_/Y _18573_/Y vssd1 vssd1 vccd1 vccd1 _18574_/X sky130_fd_sc_hd__o21a_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15044__C _15044_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15786_ _15782_/Y _15785_/Y _15946_/A vssd1 vssd1 vccd1 vccd1 _15786_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _12571_/A _12722_/A _20625_/A vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__o21ai_2
XFILLER_80_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17525_ _17537_/A _17537_/B _17934_/B _18059_/B vssd1 vssd1 vccd1 vccd1 _17528_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14737_ _16800_/D _16807_/B _14736_/X _18435_/B vssd1 vssd1 vccd1 vccd1 _14738_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11949_ _16140_/A vssd1 vssd1 vccd1 vccd1 _18434_/B sky130_fd_sc_hd__buf_4
XANTENNA__16437__A _16437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14883__C _14883_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15341__A _15442_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17456_ _17456_/A vssd1 vssd1 vccd1 vccd1 _17600_/A sky130_fd_sc_hd__buf_2
XFILLER_60_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14668_ _22968_/D vssd1 vssd1 vccd1 vccd1 _14668_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16156__B _19363_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16407_ _16407_/A _16407_/B _16407_/C vssd1 vssd1 vccd1 vccd1 _16517_/C sky130_fd_sc_hd__nand3_2
XFILLER_38_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _13619_/A _13619_/B _13619_/C vssd1 vssd1 vccd1 vccd1 _13645_/A sky130_fd_sc_hd__nand3_2
XFILLER_32_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17387_ _17299_/A _17299_/B _17299_/C _17331_/A _17331_/B vssd1 vssd1 vccd1 vccd1
+ _17387_/Y sky130_fd_sc_hd__a311oi_2
XFILLER_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14599_ _15639_/C vssd1 vssd1 vccd1 vccd1 _14599_/X sky130_fd_sc_hd__buf_2
XFILLER_158_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19126_ _12184_/X _12185_/X _18607_/C _18607_/A vssd1 vssd1 vccd1 vccd1 _19126_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16338_ _16340_/B _16297_/Y _16104_/A _16337_/X vssd1 vssd1 vccd1 vccd1 _16338_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11973__B1 _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19057_ _19059_/A _19059_/B _19058_/A _19057_/D vssd1 vssd1 vccd1 vccd1 _19063_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__23226__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16269_ _16347_/C _16018_/A _16009_/A vssd1 vssd1 vccd1 vccd1 _16270_/C sky130_fd_sc_hd__a21boi_1
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ _18016_/C _17323_/X _17324_/X _18007_/Y vssd1 vssd1 vccd1 vccd1 _18008_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_142_941 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19959_ _19957_/X _19958_/X _19952_/A _20043_/B vssd1 vssd1 vccd1 vccd1 _20072_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22970_ _23038_/S vssd1 vssd1 vccd1 vccd1 _22979_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21921_ _22292_/A _22293_/A _21921_/C vssd1 vssd1 vccd1 vccd1 _21922_/B sky130_fd_sc_hd__nand3_2
XFILLER_68_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21852_ _21852_/A _23482_/Q vssd1 vssd1 vccd1 vccd1 _21854_/A sky130_fd_sc_hd__nor2_2
XFILLER_71_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_800 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20803_ _21036_/A _20802_/Y _12674_/A _21061_/A vssd1 vssd1 vccd1 vccd1 _20973_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21783_ _21783_/A _21783_/B vssd1 vssd1 vccd1 vccd1 _21783_/X sky130_fd_sc_hd__xor2_2
XFILLER_23_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23522_ _23575_/CLK _23522_/D vssd1 vssd1 vccd1 vccd1 _23522_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18684__A1_N _12184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15251__A _15251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20734_ _20862_/B _20727_/X _20730_/Y _20733_/Y vssd1 vssd1 vccd1 vccd1 _20737_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19118__C1 _19363_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16066__B _16523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23453_ _23462_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _23453_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19669__B1 _20209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20665_ _20647_/Y _20663_/Y _20664_/X vssd1 vssd1 vccd1 vccd1 _20666_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22404_ _22405_/A _22405_/B _22405_/C vssd1 vssd1 vccd1 vccd1 _22406_/A sky130_fd_sc_hd__a21o_1
XFILLER_136_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17144__A1 _16360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23384_ _23385_/CLK _23384_/D vssd1 vssd1 vccd1 vccd1 _23384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20596_ _13205_/B _13205_/A _20594_/Y _20595_/X vssd1 vssd1 vccd1 vccd1 _20597_/C
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_109_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22335_ _22670_/D vssd1 vssd1 vccd1 vccd1 _22716_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__23217__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22266_ _22263_/X _22264_/Y _22265_/Y vssd1 vssd1 vccd1 vccd1 _22332_/C sky130_fd_sc_hd__a21oi_2
XFILLER_191_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21217_ _21217_/A vssd1 vssd1 vccd1 vccd1 _21319_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18644__A1 _19859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22197_ _22197_/A _22197_/B vssd1 vssd1 vccd1 vccd1 _22200_/B sky130_fd_sc_hd__nand2_1
XFILLER_183_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21148_ _21132_/A _21132_/B _21126_/Y _21134_/C vssd1 vssd1 vccd1 vccd1 _21148_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__21428__A _21455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17625__B _17625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19543__D _19709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21079_ _21079_/A vssd1 vssd1 vccd1 vccd1 _21430_/C sky130_fd_sc_hd__clkbuf_2
X_13970_ _14797_/B vssd1 vssd1 vccd1 vccd1 _15084_/A sky130_fd_sc_hd__clkinv_2
XFILLER_59_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14681__A2 _14672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _12921_/A _13203_/A vssd1 vssd1 vccd1 vccd1 _13088_/B sky130_fd_sc_hd__xor2_4
XANTENNA__18801__D1 _15928_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19840__B _20046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15640_ _11864_/X _11865_/X _16677_/B _16677_/C vssd1 vssd1 vccd1 vccd1 _15640_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12852_ _12932_/A _12722_/A _12725_/A vssd1 vssd1 vccd1 vccd1 _12852_/Y sky130_fd_sc_hd__o21ai_2
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19357__C1 _11747_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11803_ _11803_/A vssd1 vssd1 vccd1 vccd1 _11803_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15571_ _15571_/A _15571_/B vssd1 vssd1 vccd1 vccd1 _23496_/D sky130_fd_sc_hd__nand2_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _20528_/C vssd1 vssd1 vccd1 vccd1 _12784_/A sky130_fd_sc_hd__inv_2
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12785__A _12815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1071 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17310_ _17388_/A vssd1 vssd1 vccd1 vccd1 _17888_/A sky130_fd_sc_hd__buf_2
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ input4/X vssd1 vssd1 vccd1 vccd1 _14538_/B sky130_fd_sc_hd__clkbuf_2
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11723_/A _11741_/A _11860_/A _11733_/Y vssd1 vssd1 vccd1 vccd1 _16364_/B
+ sky130_fd_sc_hd__o211ai_4
X_18290_ _18322_/A _18349_/A _18349_/B vssd1 vssd1 vccd1 vccd1 _18292_/A sky130_fd_sc_hd__or3_1
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _19840_/A vssd1 vssd1 vccd1 vccd1 _19949_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19568__A _19568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14453_ _14446_/Y _14441_/Y _14452_/X vssd1 vssd1 vccd1 vccd1 _14453_/Y sky130_fd_sc_hd__a21oi_1
X_11665_ _11665_/A _11758_/A vssd1 vssd1 vccd1 vccd1 _11665_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15933__A2 _15605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19124__A2 _17586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13404_ _21882_/C vssd1 vssd1 vccd1 vccd1 _21793_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17172_ _17172_/A _17172_/B _17172_/C vssd1 vssd1 vccd1 vccd1 _17187_/A sky130_fd_sc_hd__nand3_2
X_14384_ _14384_/A vssd1 vssd1 vccd1 vccd1 _14458_/A sky130_fd_sc_hd__buf_2
XFILLER_31_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11596_ _19327_/B vssd1 vssd1 vccd1 vccd1 _15991_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_195_690 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16123_ _16123_/A _16123_/B vssd1 vssd1 vccd1 vccd1 _16610_/A sky130_fd_sc_hd__nand2_2
X_13335_ _23323_/Q vssd1 vssd1 vccd1 vccd1 _13377_/C sky130_fd_sc_hd__inv_2
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15146__B1 _15286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_874 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14505__A _16798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266_ _23475_/Q vssd1 vssd1 vccd1 vccd1 _13279_/A sky130_fd_sc_hd__inv_2
XFILLER_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16054_ _16054_/A vssd1 vssd1 vccd1 vccd1 _16054_/X sky130_fd_sc_hd__buf_2
XFILLER_124_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12217_ _12217_/A _12217_/B _12217_/C vssd1 vssd1 vccd1 vccd1 _12217_/X sky130_fd_sc_hd__and3_1
X_15005_ _15004_/A _15004_/B _15004_/C _15004_/D vssd1 vssd1 vccd1 vccd1 _15013_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22431__A2 _21892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ _13196_/C _13196_/A _13196_/B vssd1 vssd1 vccd1 vccd1 _13197_/X sky130_fd_sc_hd__a21o_1
XFILLER_194_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12380__B1 _12379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19813_ _19701_/B _19807_/X _19975_/A vssd1 vssd1 vccd1 vccd1 _19815_/A sky130_fd_sc_hd__o21ai_1
XFILLER_124_996 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ _15704_/B vssd1 vssd1 vccd1 vccd1 _12149_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20242__A _20290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19744_ _19572_/X _19573_/X _19588_/Y _19747_/A vssd1 vssd1 vccd1 vccd1 _19744_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12079_ _20217_/D vssd1 vssd1 vccd1 vccd1 _18163_/A sky130_fd_sc_hd__clkbuf_4
X_16956_ _16956_/A _16956_/B vssd1 vssd1 vccd1 vccd1 _16957_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11885__A2_N _11883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15907_ _15907_/A _15907_/B vssd1 vssd1 vccd1 vccd1 _16236_/A sky130_fd_sc_hd__nand2_1
X_19675_ _19675_/A _19868_/A _19675_/C vssd1 vssd1 vccd1 vccd1 _19675_/X sky130_fd_sc_hd__and3_1
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16887_ _16655_/B _16655_/C _16655_/D _16650_/Y vssd1 vssd1 vccd1 vccd1 _16888_/C
+ sky130_fd_sc_hd__a31oi_2
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18626_ _18712_/A _18721_/B _18715_/B vssd1 vssd1 vccd1 vccd1 _18707_/B sky130_fd_sc_hd__and3_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16413__A3 _17406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15838_ _15810_/X _15837_/Y _16062_/B vssd1 vssd1 vccd1 vccd1 _15895_/A sky130_fd_sc_hd__o21ai_1
XFILLER_65_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18557_ _18557_/A _18557_/B vssd1 vssd1 vccd1 vccd1 _18584_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15769_ _16447_/A _15766_/X _16126_/A _17092_/A vssd1 vssd1 vccd1 vccd1 _15843_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_75_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17508_ _18211_/D vssd1 vssd1 vccd1 vccd1 _18376_/D sky130_fd_sc_hd__buf_2
X_18488_ _18458_/Y _18465_/X _18482_/Y _18487_/X vssd1 vssd1 vccd1 vccd1 _18495_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_21_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17439_ _17439_/A _17566_/A vssd1 vssd1 vccd1 vccd1 _17440_/A sky130_fd_sc_hd__nand2_1
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15924__A2 _11865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20450_ _23557_/Q _20449_/Y _20440_/Y _20419_/X vssd1 vssd1 vccd1 vccd1 _20451_/C
+ sky130_fd_sc_hd__a22oi_1
X_19109_ _19109_/A vssd1 vssd1 vccd1 vccd1 _19442_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20381_ _20381_/A _20381_/B vssd1 vssd1 vccd1 vccd1 _20411_/A sky130_fd_sc_hd__or2_2
XANTENNA__18532__D _18945_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22120_ _21919_/Y _22167_/C _22062_/X vssd1 vssd1 vccd1 vccd1 _22130_/B sky130_fd_sc_hd__o21ai_1
XFILLER_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22051_ _22047_/B _21740_/B _13453_/A _21747_/Y vssd1 vssd1 vccd1 vccd1 _22051_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17726__A _19674_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21002_ _20885_/A _20851_/Y _21001_/Y _21130_/A vssd1 vssd1 vccd1 vccd1 _21002_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_99_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17445__B _17581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19363__D _19363_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12589__B _20532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22953_ _22953_/A vssd1 vssd1 vccd1 vccd1 _22962_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_29_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13871__B1 _13870_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21904_ _21777_/A _21777_/B _13620_/A vssd1 vssd1 vccd1 vccd1 _21913_/B sky130_fd_sc_hd__a21o_1
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22884_ _22882_/X _22873_/Y _22891_/A _22881_/Y vssd1 vssd1 vccd1 vccd1 _22885_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21835_ _21826_/X _21827_/Y _21834_/Y vssd1 vssd1 vccd1 vccd1 _21835_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21766_ _21766_/A vssd1 vssd1 vccd1 vccd1 _22508_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20717_ _20717_/A _20853_/A vssd1 vssd1 vccd1 vccd1 _20724_/A sky130_fd_sc_hd__nand2_1
X_23505_ _23518_/CLK _23505_/D vssd1 vssd1 vccd1 vccd1 _23505_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21697_ _21698_/A _21698_/C _21696_/Y vssd1 vssd1 vccd1 vccd1 _21716_/B sky130_fd_sc_hd__a21bo_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23436_ _23437_/CLK _23436_/D vssd1 vssd1 vccd1 vccd1 _23436_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12729__A2 _12722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21430__B _21432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20648_ _12765_/A _12722_/X _12754_/A _20645_/Y _20647_/Y vssd1 vssd1 vccd1 vccd1
+ _20653_/A sky130_fd_sc_hd__o221ai_1
XFILLER_109_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11949__A _16140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23367_ _23431_/CLK _23367_/D vssd1 vssd1 vccd1 vccd1 _23367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20579_ _20579_/A _20579_/B vssd1 vssd1 vccd1 vccd1 _20736_/B sky130_fd_sc_hd__nand2_1
XFILLER_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _13121_/A _13121_/B _20905_/C _13121_/C vssd1 vssd1 vccd1 vccd1 _13133_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_164_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22318_ _22184_/Y _22193_/Y _22290_/B vssd1 vssd1 vccd1 vccd1 _22318_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__20672__A1 _21431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11668__B _19363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23298_ _23298_/CLK _23298_/D vssd1 vssd1 vccd1 vccd1 _23298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12490__D _18524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ _13051_/A _23455_/Q _13051_/C vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__and3_1
XFILLER_152_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18617__A1 _16638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22249_ _22249_/A _22249_/B vssd1 vssd1 vccd1 vccd1 _22445_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12002_ _12184_/A _12185_/A _16198_/C vssd1 vssd1 vccd1 vccd1 _12002_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_127_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13883__B _23505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input47_A x[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16810_ _16810_/A vssd1 vssd1 vccd1 vccd1 _17039_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17790_ _17792_/A _17792_/B _17792_/C vssd1 vssd1 vccd1 vccd1 _17790_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12114__B1 _12113_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16741_ _16741_/A vssd1 vssd1 vccd1 vccd1 _16742_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13953_ _14396_/A _14777_/B vssd1 vssd1 vccd1 vccd1 _13953_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15306__D _15358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19460_ _19460_/A vssd1 vssd1 vccd1 vccd1 _23525_/D sky130_fd_sc_hd__clkbuf_1
X_12904_ _12904_/A _12988_/A _12988_/B vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__and3_1
XFILLER_19_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23532__CLK _23538_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16672_ _17133_/C _15936_/A _17137_/C _16745_/A _19161_/A vssd1 vssd1 vccd1 vccd1
+ _16704_/B sky130_fd_sc_hd__a32o_1
XFILLER_62_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13884_ _23351_/Q vssd1 vssd1 vccd1 vccd1 _14863_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__23126__A0 _12245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_714 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14406__A2 _15120_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18411_ _18411_/A _18411_/B _18392_/A _18410_/X vssd1 vssd1 vccd1 vccd1 _18411_/X
+ sky130_fd_sc_hd__or4bb_1
XFILLER_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15623_ _15712_/C vssd1 vssd1 vccd1 vccd1 _16187_/C sky130_fd_sc_hd__buf_2
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ _19391_/A vssd1 vssd1 vccd1 vccd1 _19601_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12835_ _12835_/A _20966_/C _12835_/C _12835_/D vssd1 vssd1 vccd1 vccd1 _12836_/B
+ sky130_fd_sc_hd__and4_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _18343_/B _18384_/B vssd1 vssd1 vccd1 vccd1 _18344_/A sky130_fd_sc_hd__and2b_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15468_/X _15538_/D _15538_/A _15564_/A vssd1 vssd1 vccd1 vccd1 _15556_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16159__A2 _15884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12766_/A vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14505_ _16798_/B vssd1 vssd1 vccd1 vccd1 _16821_/A sky130_fd_sc_hd__buf_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _20210_/A vssd1 vssd1 vccd1 vccd1 _20265_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16137__D _16634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ _18945_/C _11717_/B _11717_/C _19648_/A vssd1 vssd1 vccd1 vccd1 _12297_/A
+ sky130_fd_sc_hd__nand4_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15485_ _15483_/X _15486_/A _15511_/C _15485_/D vssd1 vssd1 vccd1 vccd1 _15493_/A
+ sky130_fd_sc_hd__and4b_1
X_12697_ _23451_/Q vssd1 vssd1 vccd1 vccd1 _20645_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__15906__A2 _16055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_638 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17224_ _19662_/C vssd1 vssd1 vccd1 vccd1 _19840_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11648_ _11648_/A _11918_/B vssd1 vssd1 vccd1 vccd1 _11809_/A sky130_fd_sc_hd__nand2_1
X_14436_ _14436_/A _14436_/B _14436_/C vssd1 vssd1 vccd1 vccd1 _14465_/B sky130_fd_sc_hd__nand3_1
Xinput12 wb_dat_i[14] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_4
XFILLER_156_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput23 wb_dat_i[24] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
Xinput34 wb_dat_i[5] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_8
XFILLER_128_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17155_ _17150_/A _17146_/X _17151_/A vssd1 vssd1 vccd1 vccd1 _17155_/X sky130_fd_sc_hd__a21o_1
XANTENNA__14590__A1 _13349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput45 x[2] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_2
XFILLER_156_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11579_ _12071_/A _16815_/A vssd1 vssd1 vccd1 vccd1 _12173_/A sky130_fd_sc_hd__nand2_2
XANTENNA__14590__B2 _15713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14367_ _14367_/A _14367_/B _14367_/C vssd1 vssd1 vccd1 vccd1 _14368_/C sky130_fd_sc_hd__nand3_1
XANTENNA__22652__A2 _13470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16106_ _16108_/B _16108_/C _16108_/A vssd1 vssd1 vccd1 vccd1 _16106_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13318_ _13318_/A _13814_/B _13318_/C vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__nand3_2
XFILLER_182_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17086_ _19703_/C vssd1 vssd1 vccd1 vccd1 _19123_/B sky130_fd_sc_hd__clkbuf_2
X_14298_ _14298_/A _14834_/A _14298_/C vssd1 vssd1 vccd1 vccd1 _14307_/A sky130_fd_sc_hd__nand3_1
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16037_ _15761_/X _15762_/Y _15763_/Y _15704_/A _12149_/A vssd1 vssd1 vccd1 vccd1
+ _16038_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13249_ _13249_/A _13680_/B vssd1 vssd1 vccd1 vccd1 _13287_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17988_ _17988_/A _17992_/C _17992_/B _17988_/D vssd1 vssd1 vccd1 vccd1 _17988_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_42_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19727_ _19719_/Y _19893_/A _19726_/X vssd1 vssd1 vccd1 vccd1 _19730_/A sky130_fd_sc_hd__a21oi_1
X_16939_ _16939_/A _16939_/B vssd1 vssd1 vccd1 vccd1 _16939_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__21915__A1 _22045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19658_ _19684_/B vssd1 vssd1 vccd1 vccd1 _19658_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23117__A0 _11604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13017__C _23451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17712__C _17960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18609_ _18599_/Y _18603_/X _18606_/Y _18608_/Y vssd1 vssd1 vccd1 vccd1 _18620_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19589_ _19572_/X _19376_/A _19573_/C _19588_/Y vssd1 vssd1 vccd1 vccd1 _19589_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13605__B1 _13603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19336__A2 _19173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21620_ _21615_/X _21618_/Y _21619_/Y vssd1 vssd1 vccd1 vccd1 _21624_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__13314__A _23476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12959__A2 _13181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21551_ _21551_/A _21592_/B vssd1 vssd1 vccd1 vccd1 _21590_/A sky130_fd_sc_hd__nand2_1
XFILLER_194_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20502_ _12601_/C _20481_/B _14615_/X vssd1 vssd1 vccd1 vccd1 _20502_/X sky130_fd_sc_hd__a21o_4
XFILLER_194_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21482_ _21482_/A _21482_/B _21482_/C vssd1 vssd1 vccd1 vccd1 _21484_/A sky130_fd_sc_hd__nand3_1
XFILLER_147_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23221_ _23221_/A vssd1 vssd1 vccd1 vccd1 _23429_/D sky130_fd_sc_hd__clkbuf_1
X_20433_ _20409_/A _20432_/Y _20431_/C vssd1 vssd1 vccd1 vccd1 _20446_/C sky130_fd_sc_hd__o21bai_2
XFILLER_181_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11769__A _15928_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18847__A1 _11822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23152_ _23399_/Q input15/X _23156_/S vssd1 vssd1 vccd1 vccd1 _23153_/A sky130_fd_sc_hd__mux2_1
X_20364_ _20364_/A vssd1 vssd1 vccd1 vccd1 _20384_/A sky130_fd_sc_hd__inv_2
XFILLER_101_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22103_ _22118_/B vssd1 vssd1 vccd1 vccd1 _22103_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17456__A _17456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_719 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23083_ _23083_/A vssd1 vssd1 vccd1 vccd1 _23368_/D sky130_fd_sc_hd__clkbuf_1
X_20295_ _20295_/A _20295_/B vssd1 vssd1 vccd1 vccd1 _20295_/X sky130_fd_sc_hd__xor2_1
XFILLER_161_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16360__A _16360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14884__A2 _14108_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22034_ _22034_/A vssd1 vssd1 vccd1 vccd1 _22392_/B sky130_fd_sc_hd__buf_2
XFILLER_114_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16510__D _18017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12647__A1 _12637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15704__A _15704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22936_ _23303_/Q input15/X _22940_/S vssd1 vssd1 vccd1 vccd1 _22937_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22867_ _22812_/A _22866_/X _22843_/A vssd1 vssd1 vccd1 vccd1 _22868_/B sky130_fd_sc_hd__a21boi_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12620_ _14655_/A vssd1 vssd1 vccd1 vccd1 _20894_/A sky130_fd_sc_hd__buf_2
XFILLER_189_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21818_ _22420_/A _13659_/Y _13777_/Y _13776_/Y vssd1 vssd1 vccd1 vccd1 _21819_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22798_ _22798_/A _22834_/A vssd1 vssd1 vccd1 vccd1 _22829_/B sky130_fd_sc_hd__or2_1
XFILLER_145_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12551_ _12563_/C vssd1 vssd1 vccd1 vccd1 _12565_/B sky130_fd_sc_hd__inv_2
XANTENNA__17889__A2 _17029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12280__C1 _12279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21749_ _22168_/A _22057_/A _21905_/B vssd1 vssd1 vccd1 vccd1 _21749_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_169_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12482_ _12447_/Y _12448_/X _12445_/C _18497_/A vssd1 vssd1 vccd1 vccd1 _12483_/A
+ sky130_fd_sc_hd__o211ai_1
X_15270_ _15270_/A _15270_/B _15326_/A vssd1 vssd1 vccd1 vccd1 _15326_/B sky130_fd_sc_hd__nand3_1
XFILLER_156_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16254__B _16254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11679__A _23583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14572__A1 _23266_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14221_ _14221_/A _14221_/B vssd1 vssd1 vccd1 vccd1 _14224_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18172__D _18172_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19846__A _19846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23419_ _23425_/CLK _23419_/D vssd1 vssd1 vccd1 vccd1 _23419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152_ _13933_/Y _13954_/Y _14150_/Y _14151_/Y vssd1 vssd1 vccd1 vccd1 _14152_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13103_ _20464_/A _12985_/Y _13102_/Y vssd1 vssd1 vccd1 vccd1 _13103_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18960_ _18862_/B _18862_/C _18958_/X _18959_/Y vssd1 vssd1 vccd1 vccd1 _18964_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_14083_ _15253_/C _14163_/B _15253_/A _14448_/A vssd1 vssd1 vccd1 vccd1 _14083_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17911_ _17911_/A _18038_/C vssd1 vssd1 vccd1 vccd1 _17916_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_782 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23518__D input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ _13034_/A _13034_/B vssd1 vssd1 vccd1 vccd1 _20557_/A sky130_fd_sc_hd__nand2_2
XFILLER_79_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18891_ _18707_/A _18707_/B _18706_/A vssd1 vssd1 vccd1 vccd1 _18892_/B sky130_fd_sc_hd__o21ai_1
XFILLER_152_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16077__A1 _16326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17842_ _17575_/X _17734_/Y _17841_/Y vssd1 vssd1 vccd1 vccd1 _17842_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14088__B1 _14863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17773_ _17773_/A _17773_/B _17773_/C _17773_/D vssd1 vssd1 vccd1 vccd1 _17773_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14985_ _15316_/A _15317_/A _15118_/A _15263_/A _14975_/C vssd1 vssd1 vccd1 vccd1
+ _14985_/X sky130_fd_sc_hd__a32o_1
XFILLER_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19512_ _19868_/A _20142_/C _19512_/C _19512_/D vssd1 vssd1 vccd1 vccd1 _19514_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16724_ _16950_/B _16723_/X _16715_/Y _16720_/Y vssd1 vssd1 vccd1 vccd1 _16724_/X
+ sky130_fd_sc_hd__o211a_1
X_13936_ _14011_/B vssd1 vssd1 vccd1 vccd1 _14044_/B sky130_fd_sc_hd__inv_2
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19443_ _19443_/A _19443_/B vssd1 vssd1 vccd1 vccd1 _19443_/Y sky130_fd_sc_hd__nor2_2
X_16655_ _16655_/A _16655_/B _16655_/C _16655_/D vssd1 vssd1 vccd1 vccd1 _16723_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13867_ _21856_/C _21856_/D _21856_/A _21856_/B vssd1 vssd1 vccd1 vccd1 _13867_/Y
+ sky130_fd_sc_hd__a22oi_4
XANTENNA__21054__C _21054_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15606_ _15599_/X _15604_/X _15920_/D _16657_/B vssd1 vssd1 vccd1 vccd1 _15612_/A
+ sky130_fd_sc_hd__o211ai_4
X_19374_ _19374_/A _19374_/B _19374_/C vssd1 vssd1 vccd1 vccd1 _19569_/A sky130_fd_sc_hd__nand3_2
X_12818_ _12975_/B _12975_/C vssd1 vssd1 vccd1 vccd1 _12819_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16586_ _16586_/A _16586_/B vssd1 vssd1 vccd1 vccd1 _16586_/Y sky130_fd_sc_hd__nand2_1
X_13798_ _13625_/X _13781_/X _13794_/Y _13797_/Y vssd1 vssd1 vccd1 vccd1 _13799_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_16_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18325_ _20265_/C vssd1 vssd1 vccd1 vccd1 _20368_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15537_ _15468_/X _15538_/D _15538_/A _15538_/B vssd1 vssd1 vccd1 vccd1 _15539_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12601_/A _12748_/X _12688_/B _23294_/Q vssd1 vssd1 vccd1 vccd1 _12997_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_72_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14891__C _15175_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_452 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18256_ _18256_/A vssd1 vssd1 vccd1 vccd1 _18417_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_175_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15468_ _15538_/C vssd1 vssd1 vccd1 vccd1 _15468_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16552__A2 _16055_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17207_ _16969_/X _16975_/Y _17365_/D _16994_/D vssd1 vssd1 vccd1 vccd1 _17524_/D
+ sky130_fd_sc_hd__o211ai_4
XFILLER_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14419_ _14492_/B _14492_/C vssd1 vssd1 vccd1 vccd1 _14495_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14563__A1 _23265_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18829__A1 _18455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18187_ _18187_/A _18187_/B vssd1 vssd1 vccd1 vccd1 _18242_/A sky130_fd_sc_hd__xor2_1
XANTENNA__14563__B2 _12678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15399_ _15391_/Y _15397_/X _15437_/B vssd1 vssd1 vccd1 vccd1 _15442_/C sky130_fd_sc_hd__o21ai_4
XFILLER_144_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17138_ _17138_/A vssd1 vssd1 vccd1 vccd1 _17307_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17069_ _17069_/A vssd1 vssd1 vccd1 vccd1 _17069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20080_ _20080_/A vssd1 vssd1 vccd1 vccd1 _20365_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19491__A _19491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14079__B1 _14188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19006__A1 _19210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17723__B _17723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19557__A2 _12509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20982_ _20984_/B _20984_/C _20984_/A vssd1 vssd1 vccd1 vccd1 _21111_/B sky130_fd_sc_hd__a21o_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22721_ _22718_/X _22722_/C _22722_/A vssd1 vssd1 vccd1 vccd1 _22723_/A sky130_fd_sc_hd__a21oi_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15043__A2 _15075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22652_ _22830_/C _13470_/X _22650_/Y _22651_/X vssd1 vssd1 vccd1 vccd1 _22661_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18517__B1 _12463_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21603_ _21601_/X _21645_/A _21599_/X vssd1 vssd1 vccd1 vccd1 _21605_/B sky130_fd_sc_hd__o21a_1
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22583_ _22580_/Y _22581_/X _22582_/X vssd1 vssd1 vccd1 vccd1 _22584_/C sky130_fd_sc_hd__o21ai_1
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22076__B _22076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21534_ _21540_/A _21540_/B vssd1 vssd1 vccd1 vccd1 _21539_/A sky130_fd_sc_hd__nor2_1
XFILLER_139_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13357__A2 _22186_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14554__A1 _23263_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21465_ _21465_/A _21465_/B _21465_/C vssd1 vssd1 vccd1 vccd1 _21465_/X sky130_fd_sc_hd__and3_1
XANTENNA__15751__B1 _15736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14554__B2 _14553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20627__A1 _20502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23204_ _15664_/C input37/X _23206_/S vssd1 vssd1 vccd1 vccd1 _23205_/A sky130_fd_sc_hd__mux2_1
X_20416_ _20362_/Y _20415_/X _20412_/B _20431_/B vssd1 vssd1 vccd1 vccd1 _20417_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_153_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21396_ _21270_/A _21270_/B _21270_/C _21274_/A vssd1 vssd1 vccd1 vccd1 _21397_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13210__C _13210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23135_ _23135_/A vssd1 vssd1 vccd1 vccd1 _23391_/D sky130_fd_sc_hd__clkbuf_1
X_20347_ _20337_/Y _20384_/B _20340_/Y _20341_/X vssd1 vssd1 vccd1 vccd1 _20356_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12317__B1 _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23066_ _23066_/A vssd1 vssd1 vccd1 vccd1 _23360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20278_ _20219_/X _20277_/Y _20220_/Y vssd1 vssd1 vccd1 vccd1 _20328_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14322__B _15017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17256__B1 _19694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16059__B2 _16479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22017_ _21744_/A _23328_/Q _13358_/X _22018_/A vssd1 vssd1 vccd1 vccd1 _22144_/A
+ sky130_fd_sc_hd__o31ai_4
XFILLER_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17633__B _17960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14085__A3 _14069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14770_ _14774_/A vssd1 vssd1 vccd1 vccd1 _14990_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22966__S _22966_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11982_ _11980_/Y _18798_/B _18468_/A vssd1 vssd1 vccd1 vccd1 _11982_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_44_511 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13721_ _13756_/B _13575_/B _13569_/Y _13720_/Y vssd1 vssd1 vccd1 vccd1 _13723_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_95_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22919_ _22919_/A vssd1 vssd1 vccd1 vccd1 _23295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16440_ _19512_/C _16436_/X _16462_/D _16523_/D _16389_/X vssd1 vssd1 vccd1 vccd1
+ _16440_/Y sky130_fd_sc_hd__a311oi_4
X_13652_ _13470_/A _13553_/A _13630_/A _13630_/B _13636_/X vssd1 vssd1 vccd1 vccd1
+ _13652_/X sky130_fd_sc_hd__o221a_1
XFILLER_182_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18508__B1 _18503_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _12929_/A _21036_/C _12930_/A vssd1 vssd1 vccd1 vccd1 _12652_/A sky130_fd_sc_hd__nand3_2
X_16371_ _17066_/C vssd1 vssd1 vccd1 vccd1 _17454_/B sky130_fd_sc_hd__clkbuf_4
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13583_ _21891_/A vssd1 vssd1 vccd1 vccd1 _22700_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_197_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18110_ _18110_/A _18110_/B vssd1 vssd1 vccd1 vccd1 _18110_/X sky130_fd_sc_hd__and2_1
XANTENNA__19181__B1 _19332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _15237_/B _15237_/A _15315_/X _15321_/X vssd1 vssd1 vccd1 vccd1 _15380_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_9_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19090_ _19090_/A _19090_/B _19090_/C _19090_/D vssd1 vssd1 vccd1 vccd1 _19090_/Y
+ sky130_fd_sc_hd__nand4_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12534_/A vssd1 vssd1 vccd1 vccd1 _18557_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18041_ _17919_/C _18040_/Y _17919_/D vssd1 vssd1 vccd1 vccd1 _18043_/A sky130_fd_sc_hd__a21bo_1
XFILLER_129_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15253_ _15253_/A _15253_/B _15253_/C vssd1 vssd1 vccd1 vccd1 _15255_/A sky130_fd_sc_hd__nand3_1
XFILLER_138_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12465_ _11931_/A _11931_/B _12464_/Y _11961_/Y vssd1 vssd1 vccd1 vccd1 _12465_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14204_ _14793_/C _14246_/B vssd1 vssd1 vccd1 vccd1 _14800_/A sky130_fd_sc_hd__nand2_2
XFILLER_193_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12396_ _12396_/A _12396_/B _12396_/C vssd1 vssd1 vccd1 vccd1 _12398_/C sky130_fd_sc_hd__nand3_4
X_15184_ _15250_/A _15187_/C _15249_/A vssd1 vssd1 vccd1 vccd1 _15185_/C sky130_fd_sc_hd__a21bo_1
XFILLER_67_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21291__A1 _20502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16298__B2 _15862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14135_ _14135_/A vssd1 vssd1 vccd1 vccd1 _14181_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19992_ _19992_/A _19992_/B _19992_/C vssd1 vssd1 vccd1 vccd1 _19992_/X sky130_fd_sc_hd__and3_1
XFILLER_152_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13505__C1 _13495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18943_ _18500_/X _18604_/X _18755_/Y _18934_/Y _18938_/X vssd1 vssd1 vccd1 vccd1
+ _18944_/B sky130_fd_sc_hd__o221ai_1
XFILLER_113_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output78_A _14720_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14066_ _14285_/B _14292_/A vssd1 vssd1 vccd1 vccd1 _14141_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17247__B1 _15884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13017_ _20628_/A _20628_/B _23451_/Q vssd1 vssd1 vccd1 vccd1 _13025_/A sky130_fd_sc_hd__nand3_1
X_18874_ _18830_/Y _18833_/Y _18871_/Y _18872_/Y _18873_/X vssd1 vssd1 vccd1 vccd1
+ _18875_/A sky130_fd_sc_hd__o221ai_4
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17825_ _17823_/Y _18139_/A _23528_/Q vssd1 vssd1 vccd1 vccd1 _17825_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_95_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13808__B1 _13603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17756_ _12088_/X _17752_/X _17876_/A vssd1 vssd1 vccd1 vccd1 _17773_/C sky130_fd_sc_hd__o21ai_1
X_14968_ _14968_/A _14968_/B _14968_/C vssd1 vssd1 vccd1 vccd1 _14968_/X sky130_fd_sc_hd__and3_1
XFILLER_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22543__A1 _13547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16707_ _16707_/A _16707_/B vssd1 vssd1 vccd1 vccd1 _16708_/B sky130_fd_sc_hd__nand2_1
X_13919_ _14193_/A vssd1 vssd1 vccd1 vccd1 _14078_/A sky130_fd_sc_hd__clkbuf_2
X_17687_ _17541_/Y _17686_/X _17682_/A vssd1 vssd1 vccd1 vccd1 _17945_/B sky130_fd_sc_hd__o21a_1
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14899_ _14899_/A _14899_/B _14908_/C _14968_/C vssd1 vssd1 vccd1 vccd1 _14900_/C
+ sky130_fd_sc_hd__nand4_1
X_19426_ _12508_/A _19116_/A _19903_/B _19425_/X vssd1 vssd1 vccd1 vccd1 _19427_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_90_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16638_ _16638_/A vssd1 vssd1 vccd1 vccd1 _16638_/X sky130_fd_sc_hd__buf_2
XANTENNA__15998__B _15998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19357_ _17742_/X _17741_/X _11749_/X _11747_/X _17581_/A vssd1 vssd1 vccd1 vccd1
+ _19357_/Y sky130_fd_sc_hd__o2111ai_4
X_16569_ _16490_/X _16052_/X _16433_/X _16757_/D vssd1 vssd1 vccd1 vccd1 _16570_/B
+ sky130_fd_sc_hd__o211ai_1
X_18308_ _18304_/Y _18306_/Y _18154_/X _18307_/Y vssd1 vssd1 vccd1 vccd1 _18362_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_188_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19288_ _19288_/A _19288_/B _19288_/C vssd1 vssd1 vccd1 vccd1 _19289_/C sky130_fd_sc_hd__nand3_1
XFILLER_148_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18239_ _18239_/A _18322_/A _18239_/C vssd1 vssd1 vccd1 vccd1 _18349_/A sky130_fd_sc_hd__nor3_2
XFILLER_148_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21250_ _21154_/Y _21158_/Y _21237_/Y vssd1 vssd1 vccd1 vccd1 _21342_/B sky130_fd_sc_hd__a21o_1
XFILLER_198_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20201_ _20201_/A _20201_/B _20201_/C vssd1 vssd1 vccd1 vccd1 _20310_/B sky130_fd_sc_hd__nand3_1
XFILLER_172_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21181_ _21181_/A vssd1 vssd1 vccd1 vccd1 _21440_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_131_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20132_ _20133_/D _20055_/B _20055_/A _20212_/A _18172_/C vssd1 vssd1 vccd1 vccd1
+ _20151_/B sky130_fd_sc_hd__a32o_1
XFILLER_104_549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11766__B _11766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20063_ _19803_/X _20210_/A _17565_/X _19668_/X vssd1 vssd1 vccd1 vccd1 _20066_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_112_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_16 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17789__A1 _16523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1084 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20798__C _20798_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18450__A2 _19859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14796__C _15195_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_831 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20965_ _20959_/X _20960_/Y _20963_/Y vssd1 vssd1 vccd1 vccd1 _20967_/A sky130_fd_sc_hd__o21ai_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17410__B1 _18503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19950__A2 _19838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22704_ _22638_/Y _22756_/B _22701_/C _22703_/Y vssd1 vssd1 vccd1 vccd1 _22707_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20896_ _20902_/C _21046_/A _21046_/B _20901_/C vssd1 vssd1 vccd1 vccd1 _21174_/A
+ sky130_fd_sc_hd__nand4_4
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22635_ _22635_/A vssd1 vssd1 vccd1 vccd1 _22703_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16085__A _19363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22566_ _22566_/A _22566_/B _22566_/C vssd1 vssd1 vccd1 vccd1 _22567_/B sky130_fd_sc_hd__nand3_1
XANTENNA__17713__A1 _19670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12250__A2 _12238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21517_ _21517_/A _21517_/B vssd1 vssd1 vccd1 vccd1 _21566_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14527__A1 _23262_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14527__B2 _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22497_ _22501_/A _22501_/B vssd1 vssd1 vccd1 vccd1 _22500_/A sky130_fd_sc_hd__nand2_1
XFILLER_142_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12250_ _12090_/A _12238_/X _12244_/X _12271_/A vssd1 vssd1 vccd1 vccd1 _12289_/B
+ sky130_fd_sc_hd__o31a_1
X_21448_ _21448_/A _21448_/B _21668_/A _21561_/B vssd1 vssd1 vccd1 vccd1 _21506_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12002__A2 _12185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20335__A _20335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _12181_/A _12181_/B _12181_/C vssd1 vssd1 vccd1 vccd1 _12211_/A sky130_fd_sc_hd__nand3_1
XFILLER_150_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21379_ _21376_/A _21376_/B _21378_/C _21378_/A vssd1 vssd1 vccd1 vccd1 _21383_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_107_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_78 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16251__C _16281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23118_ _23118_/A vssd1 vssd1 vccd1 vccd1 _23383_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__19843__B _20142_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17229__B1 _17228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23049_ _14188_/C input32/X _23051_/S vssd1 vssd1 vccd1 vccd1 _23050_/A sky130_fd_sc_hd__mux2_1
X_15940_ _15948_/B vssd1 vssd1 vccd1 vccd1 _16246_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12171__D1 _16122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18977__B1 _19505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ _18600_/A vssd1 vssd1 vccd1 vccd1 _18755_/C sky130_fd_sc_hd__buf_2
XFILLER_130_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18441__A2 _18440_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12788__A _20894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _17610_/A vssd1 vssd1 vccd1 vccd1 _17610_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11692__A _23586_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14822_ _14822_/A _14822_/B vssd1 vssd1 vccd1 vccd1 _14855_/B sky130_fd_sc_hd__nand2_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _18589_/A _18589_/B _23540_/Q vssd1 vssd1 vccd1 vccd1 _18590_/X sky130_fd_sc_hd__a21o_1
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14463__B1 _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _17699_/A _17519_/B _17540_/X vssd1 vssd1 vccd1 vccd1 _17541_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__23273__CLK _23492_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _14105_/A _14115_/Y _14756_/B vssd1 vssd1 vccd1 vccd1 _14753_/Y sky130_fd_sc_hd__o21ai_2
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _18506_/A vssd1 vssd1 vccd1 vccd1 _19334_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16204__A1 _14599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _22388_/B vssd1 vssd1 vccd1 vccd1 _13705_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_17472_ _17270_/Y _17273_/Y _17268_/C _17276_/B vssd1 vssd1 vccd1 vccd1 _17475_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14684_ _23403_/Q _14672_/X _14677_/X _23435_/Q _14683_/X vssd1 vssd1 vccd1 vccd1
+ _14684_/X sky130_fd_sc_hd__a221o_1
XANTENNA__13115__C _21174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11896_ _11896_/A _11896_/B vssd1 vssd1 vccd1 vccd1 _12130_/A sky130_fd_sc_hd__nor2_4
X_19211_ _19012_/B _19210_/Y _19013_/X vssd1 vssd1 vccd1 vccd1 _19221_/A sky130_fd_sc_hd__o21ai_1
XFILLER_189_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16423_ _16423_/A _16423_/B vssd1 vssd1 vccd1 vccd1 _16424_/C sky130_fd_sc_hd__and2_1
XFILLER_32_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13635_ _13814_/B vssd1 vssd1 vccd1 vccd1 _22172_/C sky130_fd_sc_hd__buf_2
XFILLER_13_761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19154__B1 _19505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19142_ _18944_/C _19141_/Y _19410_/B vssd1 vssd1 vccd1 vccd1 _19142_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13412__A _22270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16354_ _16575_/A _16575_/B _16576_/B vssd1 vssd1 vccd1 vccd1 _16435_/B sky130_fd_sc_hd__nand3_1
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_732 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13566_ _13650_/A _21793_/B _21793_/C _13566_/D vssd1 vssd1 vccd1 vccd1 _13566_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17825__B1_N _23528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15305_ _15305_/A vssd1 vssd1 vccd1 vccd1 _15416_/A sky130_fd_sc_hd__clkbuf_2
X_19073_ _19073_/A vssd1 vssd1 vccd1 vccd1 _19073_/Y sky130_fd_sc_hd__inv_2
X_12517_ _17592_/A _17590_/A _19364_/C vssd1 vssd1 vccd1 vccd1 _17456_/A sky130_fd_sc_hd__o21ai_4
XFILLER_121_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16285_ _16284_/Y _15716_/C _16856_/C vssd1 vssd1 vccd1 vccd1 _16860_/B sky130_fd_sc_hd__a21boi_2
XFILLER_157_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13497_ _13497_/A vssd1 vssd1 vccd1 vccd1 _13712_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18024_ _17881_/C _17881_/A _17881_/B vssd1 vssd1 vccd1 vccd1 _18024_/X sky130_fd_sc_hd__a21o_1
XFILLER_172_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15236_ _15172_/Y _15175_/X _15095_/X _15170_/Y vssd1 vssd1 vccd1 vccd1 _15237_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ _11822_/X _19040_/A _12455_/C _12422_/D vssd1 vssd1 vccd1 vccd1 _12448_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15167_ _15233_/A vssd1 vssd1 vccd1 vccd1 _15369_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12379_ _12379_/A vssd1 vssd1 vccd1 vccd1 _12379_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_181_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1024 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19209__A1 _12053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14118_ _14174_/A vssd1 vssd1 vccd1 vccd1 _14118_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19975_ _19975_/A _19975_/B vssd1 vssd1 vccd1 vccd1 _19977_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18680__A2 _12185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15098_ _14181_/X _15488_/C _15097_/Y vssd1 vssd1 vccd1 vccd1 _15107_/B sky130_fd_sc_hd__o21ai_1
XFILLER_141_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20899__B _20905_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16691__A1 _11766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18926_ _18926_/A _19288_/C vssd1 vssd1 vccd1 vccd1 _18927_/B sky130_fd_sc_hd__or2b_1
XFILLER_140_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14049_ _14054_/A _14054_/B vssd1 vssd1 vccd1 vccd1 _14049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18857_ _11926_/A _18675_/B _18958_/C _18958_/B vssd1 vssd1 vccd1 vccd1 _18858_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17640__B1 _19957_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17808_ _17662_/A _17669_/X _17807_/Y vssd1 vssd1 vccd1 vccd1 _17808_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18788_ _18788_/A _18973_/C _19804_/A vssd1 vssd1 vccd1 vccd1 _18796_/A sky130_fd_sc_hd__nand3_1
XFILLER_36_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_639 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17739_ _17285_/X _17980_/A _17750_/A vssd1 vssd1 vccd1 vccd1 _17759_/A sky130_fd_sc_hd__o21ai_1
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20750_ _21157_/A _21157_/B vssd1 vssd1 vccd1 vccd1 _20751_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15802__A _15802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14206__B1 _14089_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19409_ _19409_/A _19409_/B _19409_/C vssd1 vssd1 vccd1 vccd1 _19409_/X sky130_fd_sc_hd__and3_1
XFILLER_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14757__B2 _14876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20681_ _21431_/A _21431_/B _20681_/C vssd1 vssd1 vccd1 vccd1 _20681_/Y sky130_fd_sc_hd__nand3_1
X_22420_ _22420_/A _22420_/B _22420_/C vssd1 vssd1 vccd1 vccd1 _22420_/X sky130_fd_sc_hd__or3_1
XFILLER_149_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22351_ _22351_/A _22351_/B vssd1 vssd1 vccd1 vccd1 _22353_/B sky130_fd_sc_hd__nand2_1
XFILLER_109_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16903__C1 _15682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21302_ _21302_/A vssd1 vssd1 vccd1 vccd1 _21314_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22282_ _22656_/B _22479_/A _22279_/Y _22281_/X vssd1 vssd1 vccd1 vccd1 _22289_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__15182__A1 _14212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21233_ _21232_/Y _21333_/A _21223_/Y vssd1 vssd1 vccd1 vccd1 _21233_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__22073__C _22073_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18656__C1 _20047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16131__B1 _15998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21164_ _21069_/C _21163_/Y _21083_/B _21161_/Y vssd1 vssd1 vccd1 vccd1 _21164_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18671__A2 _18627_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20115_ _20023_/Y _20114_/Y _20185_/B vssd1 vssd1 vccd1 vccd1 _20116_/B sky130_fd_sc_hd__o21bai_1
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13496__A1 _13498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21095_ _21095_/A _21212_/B vssd1 vssd1 vccd1 vccd1 _21095_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12104__C _15682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20046_ _20046_/A vssd1 vssd1 vccd1 vccd1 _20215_/B sky130_fd_sc_hd__clkbuf_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_76 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23180__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21997_ _21997_/A vssd1 vssd1 vccd1 vccd1 _21997_/X sky130_fd_sc_hd__buf_2
XFILLER_57_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11738_/X _11740_/X _11741_/Y _11747_/X _11749_/X vssd1 vssd1 vccd1 vccd1
+ _11766_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_183_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12471__A2 _18675_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21191__B1 _13131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20948_/A _21057_/A vssd1 vssd1 vccd1 vccd1 _20950_/B sky130_fd_sc_hd__nand2_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _12105_/C vssd1 vssd1 vccd1 vccd1 _18657_/C sky130_fd_sc_hd__clkbuf_4
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20879_ _20878_/A _20878_/B _23562_/Q vssd1 vssd1 vccd1 vccd1 _21031_/A sky130_fd_sc_hd__a21o_1
X_13420_ _23473_/Q vssd1 vssd1 vccd1 vccd1 _13620_/A sky130_fd_sc_hd__inv_2
XFILLER_197_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22618_ _22619_/A _22619_/B _22616_/Y _22858_/A vssd1 vssd1 vccd1 vccd1 _22623_/B
+ sky130_fd_sc_hd__a22o_1
X_23598_ _23598_/CLK _23598_/D vssd1 vssd1 vccd1 vccd1 _23598_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20297__A2 _20243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13351_ _13348_/X _13483_/C _13349_/X _13416_/A vssd1 vssd1 vccd1 vccd1 _13351_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_194_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22549_ _22549_/A _22549_/B vssd1 vssd1 vccd1 vccd1 _22599_/B sky130_fd_sc_hd__nor2_1
XFILLER_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22264__B _22264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ _12393_/A _12393_/B _12392_/C vssd1 vssd1 vccd1 vccd1 _12303_/C sky130_fd_sc_hd__nand3_1
XANTENNA__18461__C _18461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16070_ _17248_/C _16070_/B _16070_/C _19199_/D vssd1 vssd1 vccd1 vccd1 _16075_/C
+ sky130_fd_sc_hd__nand4_2
X_13282_ _23474_/Q vssd1 vssd1 vccd1 vccd1 _13814_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15021_ _15019_/A _15195_/C _15195_/A _15081_/A _15020_/C vssd1 vssd1 vccd1 vccd1
+ _15022_/C sky130_fd_sc_hd__a32o_1
XANTENNA__11687__A _23397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ _12061_/Y _11719_/X _12391_/C _12230_/Y _12232_/X vssd1 vssd1 vccd1 vccd1
+ _12546_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_120_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11734__A1 _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ _12199_/A _12199_/B vssd1 vssd1 vccd1 vccd1 _12198_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_655 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19760_ _19745_/Y _19752_/Y _19757_/Y vssd1 vssd1 vccd1 vccd1 _19762_/A sky130_fd_sc_hd__o21ai_1
X_16972_ _16724_/X _16971_/Y _16964_/B _16964_/A vssd1 vssd1 vccd1 vccd1 _16972_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12095_ _12100_/B vssd1 vssd1 vccd1 vccd1 _12095_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23526__D _23526_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18711_ _18707_/A _18707_/B _18708_/A vssd1 vssd1 vccd1 vccd1 _18717_/A sky130_fd_sc_hd__o21ai_1
XFILLER_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15923_ _17137_/C _16198_/C _15936_/A vssd1 vssd1 vccd1 vccd1 _15923_/X sky130_fd_sc_hd__and3_1
X_19691_ _19740_/A _19880_/A vssd1 vssd1 vccd1 vccd1 _19731_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18642_ _18476_/A _18484_/X _18479_/A vssd1 vssd1 vccd1 vccd1 _19180_/B sky130_fd_sc_hd__o21a_1
XANTENNA__12949__C _20966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _12208_/A _16370_/A _15753_/B _15975_/A _15993_/A vssd1 vssd1 vccd1 vccd1
+ _15859_/B sky130_fd_sc_hd__o221ai_1
XFILLER_49_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12311__A _12311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _14805_/A _14805_/B vssd1 vssd1 vccd1 vccd1 _14928_/A sky130_fd_sc_hd__nand2_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _18571_/Y _18572_/X _19089_/A _12545_/Y vssd1 vssd1 vccd1 vccd1 _18573_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _15785_/A _15785_/B _15785_/C vssd1 vssd1 vccd1 vccd1 _15785_/Y sky130_fd_sc_hd__nand3_2
XFILLER_18_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12997_ _12997_/A _20620_/C _12997_/C vssd1 vssd1 vccd1 vccd1 _20625_/A sky130_fd_sc_hd__nand3_2
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _17524_/A _17524_/B _17524_/C _17524_/D vssd1 vssd1 vccd1 vccd1 _17934_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_33_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _23595_/Q _23596_/Q vssd1 vssd1 vccd1 vccd1 _14736_/X sky130_fd_sc_hd__or2_1
X_11948_ _11948_/A vssd1 vssd1 vccd1 vccd1 _11948_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _17845_/C _17586_/A _17587_/A vssd1 vssd1 vccd1 vccd1 _17597_/A sky130_fd_sc_hd__nand3_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _14688_/A vssd1 vssd1 vccd1 vccd1 _14667_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11879_ _12183_/A vssd1 vssd1 vccd1 vccd1 _18952_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__16156__C _17057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16406_ _16383_/X _16386_/X _16396_/A _16396_/B vssd1 vssd1 vccd1 vccd1 _16407_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__15400__A2 _15442_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13618_ _13610_/Y _13609_/X _22269_/C _13616_/Y _13816_/A vssd1 vssd1 vccd1 vccd1
+ _13619_/C sky130_fd_sc_hd__o2111ai_2
X_17386_ _17221_/X _17222_/Y _17289_/Y _17292_/Y vssd1 vssd1 vccd1 vccd1 _17386_/X
+ sky130_fd_sc_hd__o211a_1
X_14598_ _23423_/Q vssd1 vssd1 vccd1 vccd1 _15639_/C sky130_fd_sc_hd__buf_2
XFILLER_125_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19125_ _19125_/A _19125_/B _19125_/C vssd1 vssd1 vccd1 vccd1 _19391_/A sky130_fd_sc_hd__nand3_4
XFILLER_146_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16337_ _16422_/B _16336_/X _16425_/A _16099_/Y vssd1 vssd1 vccd1 vccd1 _16337_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_185_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13962__A2 _13945_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13549_ _13531_/X _13507_/A _13548_/X _13540_/Y _13543_/Y vssd1 vssd1 vccd1 vccd1
+ _13697_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_72_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11973__A1 _11971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19056_ _19058_/B vssd1 vssd1 vccd1 vccd1 _19057_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16268_ _16268_/A _16268_/B _16268_/C _16268_/D vssd1 vssd1 vccd1 vccd1 _16586_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_161_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16172__B _17445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18007_ _16665_/X _17029_/X _17712_/B _17712_/A _17723_/B vssd1 vssd1 vccd1 vccd1
+ _18007_/Y sky130_fd_sc_hd__o2111ai_2
X_15219_ _15219_/A _15219_/B vssd1 vssd1 vccd1 vccd1 _23275_/D sky130_fd_sc_hd__xnor2_1
XFILLER_160_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18638__C1 _18479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18102__A1 _17766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16199_ _16183_/A _16194_/Y _16198_/X vssd1 vssd1 vccd1 vccd1 _16199_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_160_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16664__A1 _16458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16664__B2 _16663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19958_ _12237_/A _19953_/A _20079_/A _19848_/Y _19847_/X vssd1 vssd1 vccd1 vccd1
+ _19958_/X sky130_fd_sc_hd__o311a_1
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18909_ _19090_/B _19091_/A _18909_/C vssd1 vssd1 vccd1 vccd1 _18910_/C sky130_fd_sc_hd__nand3_1
XFILLER_132_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19889_ _19889_/A _19889_/B _19889_/C vssd1 vssd1 vccd1 vccd1 _19897_/B sky130_fd_sc_hd__nand3_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21920_ _13465_/A _13410_/A _21919_/Y vssd1 vssd1 vccd1 vccd1 _21920_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13317__A _13766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21851_ _22107_/D _21981_/A _21858_/D _21972_/A vssd1 vssd1 vccd1 vccd1 _21861_/B
+ sky130_fd_sc_hd__nand4b_1
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20802_ _21047_/A _20800_/B _13151_/B vssd1 vssd1 vccd1 vccd1 _20802_/Y sky130_fd_sc_hd__a21oi_1
X_21782_ _21782_/A _21782_/B _21782_/C vssd1 vssd1 vccd1 vccd1 _21805_/C sky130_fd_sc_hd__nand3_1
XANTENNA__17450__C _17450_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12875__B _12875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23521_ _23582_/CLK _23521_/D vssd1 vssd1 vccd1 vccd1 _23521_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20733_ _20714_/A _20714_/B _20715_/C _20731_/Y _20732_/Y vssd1 vssd1 vccd1 vccd1
+ _20733_/Y sky130_fd_sc_hd__a221oi_4
XFILLER_168_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19118__B1 _19363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13052__A _13052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16066__C _16066_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19669__A1 _19670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23452_ _23559_/CLK hold13/X vssd1 vssd1 vccd1 vccd1 _23452_/Q sky130_fd_sc_hd__dfxtp_2
X_20664_ _20639_/C _12689_/X _12640_/X _12692_/Y _12792_/A vssd1 vssd1 vccd1 vccd1
+ _20664_/X sky130_fd_sc_hd__a311o_1
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19669__B2 _16066_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22403_ _22403_/A vssd1 vssd1 vccd1 vccd1 _22405_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_183_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17459__A _20049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23383_ _23385_/CLK _23383_/D vssd1 vssd1 vccd1 vccd1 _23383_/Q sky130_fd_sc_hd__dfxtp_1
X_20595_ _20595_/A _20595_/B _20595_/C vssd1 vssd1 vccd1 vccd1 _20595_/X sky130_fd_sc_hd__and3_1
XFILLER_13_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17144__A2 _17635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22334_ _22221_/B _22226_/X _22357_/A _22357_/B vssd1 vssd1 vccd1 vccd1 _22341_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__17695__A3 _23526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22265_ _22510_/B _22263_/B _22264_/Y _22434_/A vssd1 vssd1 vccd1 vccd1 _22265_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__14902__A1 _14588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21216_ _21216_/A vssd1 vssd1 vccd1 vccd1 _21221_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22196_ _22158_/A _22166_/Y _22176_/A vssd1 vssd1 vccd1 vccd1 _22200_/A sky130_fd_sc_hd__a21bo_1
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21147_ _21147_/A _21147_/B vssd1 vssd1 vccd1 vccd1 _23544_/D sky130_fd_sc_hd__xor2_1
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17625__C _17625_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21078_ _21078_/A _21163_/A _21163_/B vssd1 vssd1 vccd1 vccd1 _21082_/B sky130_fd_sc_hd__nand3_4
XFILLER_150_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20029_ _20196_/C vssd1 vssd1 vccd1 vccd1 _20029_/Y sky130_fd_sc_hd__inv_2
X_12920_ _12812_/A _12812_/B _12810_/Y _12817_/B vssd1 vssd1 vccd1 vccd1 _13203_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_24_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19840__C _20047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12851_ _12851_/A _23450_/Q _12851_/C _20620_/C vssd1 vssd1 vccd1 vccd1 _12851_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_74_778 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19357__B1 _11749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _12419_/A vssd1 vssd1 vccd1 vccd1 _19123_/C sky130_fd_sc_hd__buf_2
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _23507_/Q _15569_/B _23508_/Q vssd1 vssd1 vccd1 vccd1 _15571_/B sky130_fd_sc_hd__a21bo_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _23453_/Q vssd1 vssd1 vccd1 vccd1 _20528_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_54_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ input1/X vssd1 vssd1 vccd1 vccd1 _14535_/A sky130_fd_sc_hd__clkbuf_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _23586_/Q vssd1 vssd1 vccd1 vccd1 _11733_/Y sky130_fd_sc_hd__clkinv_2
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16040__C1 _15682_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17240_ _19949_/D vssd1 vssd1 vccd1 vccd1 _19957_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_30_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _15208_/A _14472_/D _15310_/B _14469_/D vssd1 vssd1 vccd1 vccd1 _14452_/X
+ sky130_fd_sc_hd__and4_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11664_ _11823_/B vssd1 vssd1 vccd1 vccd1 _11980_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13403_ _21909_/C vssd1 vssd1 vccd1 vccd1 _22035_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_186_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19124__A3 _17587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17171_ _17334_/A _17335_/A _17169_/Y _17170_/X vssd1 vssd1 vccd1 vccd1 _17172_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__22664__B1 _21829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14383_ _14334_/Y _14381_/Y _14457_/A _14806_/A vssd1 vssd1 vccd1 vccd1 _14390_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_70_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11595_ _12474_/A vssd1 vssd1 vccd1 vccd1 _19327_/B sky130_fd_sc_hd__buf_2
XFILLER_167_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16122_ _16122_/A _16122_/B _16314_/B _16314_/C vssd1 vssd1 vccd1 vccd1 _16123_/B
+ sky130_fd_sc_hd__nand4_2
X_13334_ _21902_/C vssd1 vssd1 vccd1 vccd1 _22028_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23461__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21219__A1 _21218_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16053_ _12040_/X _16035_/X _16039_/A _16310_/B vssd1 vssd1 vccd1 vccd1 _16060_/A
+ sky130_fd_sc_hd__a22o_1
X_13265_ _23474_/Q vssd1 vssd1 vccd1 vccd1 _13495_/A sky130_fd_sc_hd__inv_2
XANTENNA__12306__A _12306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20427__C1 _20371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15004_ _15004_/A _15004_/B _15004_/C _15004_/D vssd1 vssd1 vccd1 vccd1 _15013_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_170_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12216_ _12216_/A _12216_/B vssd1 vssd1 vccd1 vccd1 _12217_/A sky130_fd_sc_hd__nand2_1
XANTENNA__21619__A _23571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13196_ _13196_/A _13196_/B _13196_/C vssd1 vssd1 vccd1 vccd1 _13196_/Y sky130_fd_sc_hd__nand3_1
XFILLER_151_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19812_ _19190_/A _12518_/X _19811_/Y vssd1 vssd1 vccd1 vccd1 _19975_/A sky130_fd_sc_hd__o21ai_2
XFILLER_123_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12147_ _12147_/A vssd1 vssd1 vccd1 vccd1 _12147_/X sky130_fd_sc_hd__buf_2
XANTENNA__14521__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20242__B _20242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19743_ _19743_/A vssd1 vssd1 vccd1 vccd1 _19743_/X sky130_fd_sc_hd__clkbuf_2
X_12078_ _20142_/D vssd1 vssd1 vccd1 vccd1 _20217_/D sky130_fd_sc_hd__clkbuf_2
X_16955_ _17173_/B _16954_/Y _16951_/A _16944_/A vssd1 vssd1 vccd1 vccd1 _16955_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15906_ _16054_/A _16055_/A _15618_/X _15621_/X _16866_/A vssd1 vssd1 vccd1 vccd1
+ _15907_/B sky130_fd_sc_hd__o221a_1
X_19674_ _19674_/A _19674_/B _19674_/C vssd1 vssd1 vccd1 vccd1 _19674_/Y sky130_fd_sc_hd__nand3_1
X_16886_ _16877_/X _16878_/Y _16884_/Y _16894_/A vssd1 vssd1 vccd1 vccd1 _16888_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__12041__A _12475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18625_ _18715_/B _18712_/A _18721_/B vssd1 vssd1 vccd1 vccd1 _18707_/A sky130_fd_sc_hd__a21oi_1
XFILLER_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15837_ _16062_/B _16073_/B vssd1 vssd1 vccd1 vccd1 _15837_/Y sky130_fd_sc_hd__nand2_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18556_ _18545_/Y _18548_/Y _18560_/A vssd1 vssd1 vccd1 vccd1 _18557_/A sky130_fd_sc_hd__o21ai_1
X_15768_ _15841_/B vssd1 vssd1 vccd1 vccd1 _17092_/A sky130_fd_sc_hd__buf_2
XFILLER_46_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17507_ _18211_/C vssd1 vssd1 vccd1 vccd1 _18376_/B sky130_fd_sc_hd__buf_2
X_14719_ _23381_/Q _14635_/A _14718_/X vssd1 vssd1 vccd1 vccd1 _14719_/X sky130_fd_sc_hd__o21a_1
X_18487_ _11670_/X _12279_/A _18474_/X _19491_/A _18473_/X vssd1 vssd1 vccd1 vccd1
+ _18487_/X sky130_fd_sc_hd__o221a_1
XFILLER_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15699_ _15699_/A _16027_/B _15983_/A _15831_/A vssd1 vssd1 vccd1 vccd1 _15699_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_36_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17438_ _17249_/X _17250_/X _16027_/D _17569_/A vssd1 vssd1 vccd1 vccd1 _17566_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_177_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17369_ _17369_/A _17369_/B _17369_/C _17369_/D vssd1 vssd1 vccd1 vccd1 _17522_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_118_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19108_ _19108_/A vssd1 vssd1 vccd1 vccd1 _19293_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20380_ _20327_/A _20329_/B _20331_/A _20331_/B vssd1 vssd1 vccd1 vccd1 _20381_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__16334__B1 _16071_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19039_ _18875_/B _18875_/C _18840_/Y _18828_/Y vssd1 vssd1 vccd1 vccd1 _19066_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19494__A _19840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22958__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22050_ _22037_/X _22153_/A _22270_/C _22479_/B _22040_/Y vssd1 vssd1 vccd1 vccd1
+ _22050_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_86_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21001_ _21132_/A _21131_/B vssd1 vssd1 vccd1 vccd1 _21001_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15527__A _15527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17445__C _18778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12123__A1 _12117_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22952_ _22952_/A vssd1 vssd1 vccd1 vccd1 _23310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21903_ _22562_/A _22024_/C _22031_/A vssd1 vssd1 vccd1 vccd1 _22040_/A sky130_fd_sc_hd__nand3_2
XFILLER_44_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22883_ _22891_/A _22881_/Y _22882_/X _22873_/Y vssd1 vssd1 vccd1 vccd1 _22885_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18276__C _18276_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21834_ _13848_/A _13848_/B _21833_/X vssd1 vssd1 vccd1 vccd1 _21834_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_70_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18011__B1 _20164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21765_ _13392_/A _13392_/B _13469_/A vssd1 vssd1 vccd1 vccd1 _21783_/A sky130_fd_sc_hd__a21o_1
XFILLER_169_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23504_ _23510_/CLK _23504_/D vssd1 vssd1 vccd1 vccd1 _23504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20716_ _20716_/A _20716_/B _20716_/C vssd1 vssd1 vccd1 vccd1 _20853_/A sky130_fd_sc_hd__nand3_1
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21696_ _21698_/B _21704_/D vssd1 vssd1 vccd1 vccd1 _21696_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22095__A _22754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23435_ _23435_/CLK _23435_/D vssd1 vssd1 vccd1 vccd1 _23435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20647_ _12674_/A _12849_/A _20646_/Y vssd1 vssd1 vccd1 vccd1 _20647_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16093__A _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11937__A1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__B2 _11936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20578_ _20578_/A _20578_/B _20578_/C vssd1 vssd1 vccd1 vccd1 _20578_/X sky130_fd_sc_hd__and3_1
X_23366_ _23431_/CLK _23366_/D vssd1 vssd1 vccd1 vccd1 _23366_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18865__A2 _18840_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22317_ _22291_/Y _22312_/Y _22315_/Y _22316_/Y vssd1 vssd1 vccd1 vccd1 _22332_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__20672__A2 _21431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12771__D _12845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16821__A _16821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23297_ _23297_/CLK _23297_/D vssd1 vssd1 vccd1 vccd1 _23297_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12126__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22949__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23071__A0 _14632_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13050_ _13052_/A _23454_/Q _13052_/C vssd1 vssd1 vccd1 vccd1 _20529_/A sky130_fd_sc_hd__nand3_1
XANTENNA__18617__A2 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22248_ _22348_/B _22348_/C vssd1 vssd1 vccd1 vccd1 _22249_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12001_ _19000_/B vssd1 vssd1 vccd1 vccd1 _16198_/C sky130_fd_sc_hd__buf_2
XANTENNA__11965__A _18506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22179_ _22037_/X _22474_/C _22051_/X vssd1 vssd1 vccd1 vccd1 _22179_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16740_ _16740_/A vssd1 vssd1 vccd1 vccd1 _16744_/B sky130_fd_sc_hd__clkbuf_2
X_13952_ _14246_/B vssd1 vssd1 vccd1 vccd1 _14777_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _12991_/A _12988_/A _12988_/B vssd1 vssd1 vccd1 vccd1 _12903_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__21174__A _21174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16671_ _16671_/A _16671_/B vssd1 vssd1 vccd1 vccd1 _16745_/A sky130_fd_sc_hd__nand2_1
X_13883_ _14469_/D _23505_/Q vssd1 vssd1 vccd1 vccd1 _14007_/A sky130_fd_sc_hd__nand2_1
XANTENNA__23126__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18410_ _18410_/A _18382_/C vssd1 vssd1 vccd1 vccd1 _18410_/X sky130_fd_sc_hd__or2b_1
XFILLER_98_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15622_ _15622_/A vssd1 vssd1 vccd1 vccd1 _15761_/A sky130_fd_sc_hd__buf_2
X_19390_ _19355_/Y _19468_/A _19600_/A vssd1 vssd1 vccd1 vccd1 _19390_/X sky130_fd_sc_hd__and3b_1
X_12834_ _20966_/C _13157_/B _12835_/C _12835_/A vssd1 vssd1 vccd1 vccd1 _12836_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_34_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _18341_/A _18341_/B vssd1 vssd1 vccd1 vccd1 _18384_/B sky130_fd_sc_hd__nand2_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15468_/X _15446_/A _15538_/B vssd1 vssd1 vccd1 vccd1 _15564_/A sky130_fd_sc_hd__a21boi_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12765_/A vssd1 vssd1 vccd1 vccd1 _13122_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12968__A3 _21358_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14504_ _15735_/C vssd1 vssd1 vccd1 vccd1 _16798_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_187_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18272_ _18272_/A _18279_/B _19425_/C _20268_/D vssd1 vssd1 vccd1 vccd1 _18272_/X
+ sky130_fd_sc_hd__and4_1
X_11716_ _19323_/A vssd1 vssd1 vccd1 vccd1 _19648_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15455_/A _15096_/A _15096_/B _15483_/C vssd1 vssd1 vccd1 vccd1 _15486_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12696_ _12696_/A vssd1 vssd1 vccd1 vccd1 _20663_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17223_ _17077_/B _17070_/X _17069_/X _17068_/X vssd1 vssd1 vccd1 vccd1 _17232_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14435_ _14465_/C _14465_/D vssd1 vssd1 vccd1 vccd1 _14435_/X sky130_fd_sc_hd__and2_1
X_11647_ _11960_/B _11647_/B vssd1 vssd1 vccd1 vccd1 _12147_/A sky130_fd_sc_hd__nand2_4
XFILLER_168_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 wb_dat_i[15] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1042 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13420__A _23473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17154_ _12323_/X _17230_/A _17307_/A _17150_/B _17140_/Y vssd1 vssd1 vccd1 vccd1
+ _17154_/X sky130_fd_sc_hd__o311a_1
Xinput24 wb_dat_i[25] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_2
XANTENNA__16316__B1 _15972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput35 wb_dat_i[6] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_4
X_14366_ _14367_/C _14367_/B _14367_/A vssd1 vssd1 vccd1 vccd1 _14368_/B sky130_fd_sc_hd__a21o_1
XFILLER_156_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11578_ _23589_/Q vssd1 vssd1 vccd1 vccd1 _16815_/A sky130_fd_sc_hd__buf_2
XFILLER_122_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput46 x[3] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16867__A1 _18859_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16105_ _16077_/X _16340_/A _16340_/C vssd1 vssd1 vccd1 vccd1 _16108_/A sky130_fd_sc_hd__a21boi_2
XFILLER_122_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13317_ _13766_/A _13766_/B vssd1 vssd1 vccd1 vccd1 _13491_/A sky130_fd_sc_hd__nand2_1
X_17085_ _12509_/X _16377_/X _17077_/A vssd1 vssd1 vccd1 vccd1 _17089_/C sky130_fd_sc_hd__o21ai_2
XFILLER_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14297_ _14469_/D vssd1 vssd1 vccd1 vccd1 _14298_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__23062__A0 _14188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16036_ _16447_/A _15766_/X _15706_/A _15682_/B vssd1 vssd1 vccd1 vccd1 _16300_/A
+ sky130_fd_sc_hd__o211ai_2
X_13248_ _13656_/B vssd1 vssd1 vccd1 vccd1 _13680_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_171_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11875__A _11875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18683__A1_N _18474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13179_ _13179_/A vssd1 vssd1 vccd1 vccd1 _20775_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17987_ _17986_/D _17986_/B _17611_/X _20210_/D vssd1 vssd1 vccd1 vccd1 _17992_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_111_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19726_ _19560_/Y _19555_/Y _19556_/X _19546_/Y vssd1 vssd1 vccd1 vccd1 _19726_/X
+ sky130_fd_sc_hd__o31a_1
X_16938_ _16934_/X _16936_/Y _16937_/Y _16924_/Y vssd1 vssd1 vccd1 vccd1 _16948_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__21915__A2 _22045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17044__A1 _15742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19657_ _19304_/X _19307_/Y _19655_/X _19855_/C _19525_/D vssd1 vssd1 vccd1 vccd1
+ _19684_/B sky130_fd_sc_hd__o221ai_4
XFILLER_26_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16869_ _16635_/B _16614_/Y _16617_/X _16153_/B vssd1 vssd1 vccd1 vccd1 _16870_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_26_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17712__D _17712_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23117__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18608_ _18607_/X _18534_/Y _18537_/Y _18536_/X vssd1 vssd1 vccd1 vccd1 _18608_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_19588_ _19588_/A _19588_/B vssd1 vssd1 vccd1 vccd1 _19588_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14802__B1 _15301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18539_ _18540_/A _18540_/B _18540_/C vssd1 vssd1 vccd1 vccd1 _18721_/A sky130_fd_sc_hd__a21oi_2
XFILLER_178_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18824__C _19539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15810__A _16019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21550_ _21548_/X _21504_/A _21545_/X _21547_/X vssd1 vssd1 vccd1 vccd1 _21592_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_20_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20501_ _20501_/A vssd1 vssd1 vccd1 vccd1 _20501_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_166_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21481_ _21346_/X _21423_/Y _21576_/A vssd1 vssd1 vccd1 vccd1 _21482_/A sky130_fd_sc_hd__o21ai_1
XFILLER_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20432_ _20411_/A _20415_/A _20411_/C vssd1 vssd1 vccd1 vccd1 _20432_/Y sky130_fd_sc_hd__a21oi_1
X_23220_ _16780_/B input13/X _23228_/S vssd1 vssd1 vccd1 vccd1 _23221_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20363_ _20335_/A _20363_/B vssd1 vssd1 vccd1 vccd1 _20364_/A sky130_fd_sc_hd__and2b_1
XFILLER_106_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23151_ _23151_/A vssd1 vssd1 vccd1 vccd1 _23398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22102_ _22102_/A _22240_/B _22102_/C vssd1 vssd1 vccd1 vccd1 _22118_/B sky130_fd_sc_hd__nand3_2
XFILLER_134_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23082_ _23368_/Q input16/X _23084_/S vssd1 vssd1 vccd1 vccd1 _23083_/A sky130_fd_sc_hd__mux2_1
X_20294_ _20252_/A _20252_/B _20243_/A _20243_/B vssd1 vssd1 vccd1 vccd1 _20294_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__20163__A _20217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22033_ _22033_/A vssd1 vssd1 vccd1 vccd1 _22391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12647__A2 _12640_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22935_ _22935_/A vssd1 vssd1 vccd1 vccd1 _23302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16088__A _16423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23108__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22866_ _22788_/X _22805_/X _22789_/X _22843_/B vssd1 vssd1 vccd1 vccd1 _22866_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21817_ _13777_/Y _13776_/Y _21816_/X vssd1 vssd1 vccd1 vccd1 _21817_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_197_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22797_ _22797_/A _22797_/B _22797_/C vssd1 vssd1 vccd1 vccd1 _22834_/A sky130_fd_sc_hd__nor3_1
XFILLER_58_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _12370_/Y _12384_/Y _12398_/C _12549_/Y vssd1 vssd1 vccd1 vccd1 _12563_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_24_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15349__A1 _15298_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12280__B1 _11717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21748_ _22020_/B vssd1 vssd1 vccd1 vccd1 _22168_/A sky130_fd_sc_hd__buf_2
XFILLER_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16546__B1 _15731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17743__C1 _17243_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ _12481_/A _12481_/B vssd1 vssd1 vccd1 vccd1 _12487_/A sky130_fd_sc_hd__nand2_1
XFILLER_184_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21679_ _21694_/C vssd1 vssd1 vccd1 vccd1 _21679_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14220_ _14220_/A _14220_/B vssd1 vssd1 vccd1 vccd1 _14221_/A sky130_fd_sc_hd__nand2_1
X_23418_ _23428_/CLK _23418_/D vssd1 vssd1 vccd1 vccd1 _23418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18838__A2 _19656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_886 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14151_ _13985_/X _13989_/Y _13971_/X vssd1 vssd1 vccd1 vccd1 _14151_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23349_ _23349_/CLK _23349_/D vssd1 vssd1 vccd1 vccd1 _23349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ _12984_/A _12984_/B _13106_/B vssd1 vssd1 vccd1 vccd1 _13102_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_180_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14082_ _14774_/C vssd1 vssd1 vccd1 vccd1 _14448_/A sky130_fd_sc_hd__buf_2
X_17910_ _17911_/A _18038_/C _17916_/C _17916_/A vssd1 vssd1 vccd1 vccd1 _17915_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _12893_/Y _12894_/X _12860_/A vssd1 vssd1 vccd1 vccd1 _13034_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__19862__A _19862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18890_ _18884_/A _18884_/B _18889_/Y _19062_/A vssd1 vssd1 vccd1 vccd1 _18893_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_133_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17841_ _17742_/X _17741_/X _17414_/C _18778_/A _17414_/D vssd1 vssd1 vccd1 vccd1
+ _17841_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_117_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17772_ _17747_/X _17758_/Y _17768_/Y _17771_/Y vssd1 vssd1 vccd1 vccd1 _17782_/B
+ sky130_fd_sc_hd__o211ai_4
X_14984_ _14984_/A vssd1 vssd1 vccd1 vccd1 _15263_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19511_ _19511_/A vssd1 vssd1 vccd1 vccd1 _20142_/C sky130_fd_sc_hd__clkbuf_4
X_16723_ _16723_/A _16723_/B _16723_/C vssd1 vssd1 vccd1 vccd1 _16723_/X sky130_fd_sc_hd__and3_1
X_13935_ _14172_/A _14172_/B _14774_/C vssd1 vssd1 vccd1 vccd1 _14058_/A sky130_fd_sc_hd__nand3_1
XFILLER_93_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_704 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19442_ _19442_/A _19442_/B vssd1 vssd1 vccd1 vccd1 _19442_/Y sky130_fd_sc_hd__nand2_2
X_16654_ _16175_/B _16175_/C _16175_/A vssd1 vssd1 vccd1 vccd1 _16723_/B sky130_fd_sc_hd__a21oi_1
X_13866_ _21840_/A _21839_/B _21839_/A vssd1 vssd1 vccd1 vccd1 _21856_/B sky130_fd_sc_hd__nand3_2
XFILLER_179_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21054__D _21054_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15605_ _15605_/A vssd1 vssd1 vccd1 vccd1 _15920_/D sky130_fd_sc_hd__inv_2
X_12817_ _12817_/A _12817_/B vssd1 vssd1 vccd1 vccd1 _12975_/C sky130_fd_sc_hd__nor2_1
XFILLER_90_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19373_ _19126_/X _19121_/X _19123_/Y vssd1 vssd1 vccd1 vccd1 _19374_/C sky130_fd_sc_hd__a21boi_1
X_16585_ _16585_/A vssd1 vssd1 vccd1 vccd1 _16585_/Y sky130_fd_sc_hd__inv_2
X_13797_ _13797_/A _13797_/B vssd1 vssd1 vccd1 vccd1 _13797_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18324_ _18324_/A _18335_/C _18324_/C _18339_/A vssd1 vssd1 vccd1 vccd1 _18339_/B
+ sky130_fd_sc_hd__nand4_1
X_15536_ _15536_/A _15536_/B _15536_/C _15225_/B vssd1 vssd1 vccd1 vccd1 _15538_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_31_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12748_/A vssd1 vssd1 vccd1 vccd1 _12748_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17734__C1 _17845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18255_ _18207_/X _18208_/X _18302_/B _18254_/Y vssd1 vssd1 vccd1 vccd1 _18364_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_176_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15467_ _15467_/A _15467_/B _15467_/C vssd1 vssd1 vccd1 vccd1 _15501_/A sky130_fd_sc_hd__nand3_1
XFILLER_31_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12679_ _12577_/A _12678_/Y _13014_/A vssd1 vssd1 vccd1 vccd1 _12680_/A sky130_fd_sc_hd__a21oi_2
XFILLER_187_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17206_ _17024_/Y _17027_/Y _17365_/D vssd1 vssd1 vccd1 vccd1 _17524_/C sky130_fd_sc_hd__o21bai_4
XFILLER_147_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14418_ _14418_/A _14418_/B _14418_/C vssd1 vssd1 vccd1 vccd1 _14492_/B sky130_fd_sc_hd__nand3_1
XFILLER_191_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18186_ _18186_/A _18186_/B vssd1 vssd1 vccd1 vccd1 _18187_/B sky130_fd_sc_hd__or2_1
X_15398_ _15391_/Y _15396_/X _15335_/B _15395_/Y vssd1 vssd1 vccd1 vccd1 _15437_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__18829__A2 _18461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17137_ _19323_/A _17625_/B _17137_/C vssd1 vssd1 vccd1 vccd1 _17138_/A sky130_fd_sc_hd__nand3_1
XANTENNA__21833__A1 _22754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14349_ _14358_/C _14358_/B _14349_/C _14349_/D vssd1 vssd1 vccd1 vccd1 _14350_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_156_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17068_ _17068_/A vssd1 vssd1 vccd1 vccd1 _17068_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16019_ _16019_/A _16019_/B vssd1 vssd1 vccd1 vccd1 _16073_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20133__D _20133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_904 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19006__A2 _19191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17723__C _17723_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19709_ _19709_/A _19709_/B _19709_/C vssd1 vssd1 vccd1 vccd1 _19819_/B sky130_fd_sc_hd__and3_1
XANTENNA__11837__B1 _19180_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15524__B _15525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20981_ _20989_/A _20989_/B _20994_/C vssd1 vssd1 vccd1 vccd1 _20981_/Y sky130_fd_sc_hd__o21ai_1
X_22720_ _22720_/A _22720_/B vssd1 vssd1 vccd1 vccd1 _22722_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_523 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21542__A _21542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1097 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22651_ _22650_/A _22650_/B _22713_/D _22712_/A vssd1 vssd1 vccd1 vccd1 _22651_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14251__B2 _14867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21602_ _21602_/A _21602_/B vssd1 vssd1 vccd1 vccd1 _21645_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22582_ _21997_/X _22461_/X _22368_/Y _22489_/C vssd1 vssd1 vccd1 vccd1 _22582_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22076__C _22218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21533_ _21541_/A _23569_/Q _21541_/C vssd1 vssd1 vccd1 vccd1 _21540_/B sky130_fd_sc_hd__and3_1
XFILLER_166_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14156__A _14230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22077__A1 _22218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12014__B1 _11841_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21464_ _21464_/A _21464_/B vssd1 vssd1 vccd1 vccd1 _21465_/C sky130_fd_sc_hd__nand2_1
XANTENNA__15751__A1 _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15751__B2 _15738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23203_ _23203_/A vssd1 vssd1 vccd1 vccd1 _23421_/D sky130_fd_sc_hd__clkbuf_1
X_20415_ _20415_/A _20415_/B _20452_/B vssd1 vssd1 vccd1 vccd1 _20415_/X sky130_fd_sc_hd__and3_1
XFILLER_175_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20627__A2 _20504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21395_ _21399_/B vssd1 vssd1 vccd1 vccd1 _21424_/B sky130_fd_sc_hd__inv_2
XFILLER_190_940 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16371__A _17066_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23134_ _12100_/B input38/X _23134_/S vssd1 vssd1 vccd1 vccd1 _23135_/A sky130_fd_sc_hd__mux2_1
X_20346_ _20342_/Y _20345_/X _23554_/Q vssd1 vssd1 vccd1 vccd1 _20359_/C sky130_fd_sc_hd__o21bai_1
XANTENNA__16161__D1 _16499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12317__A1 _11747_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20277_ _20287_/B _20277_/B vssd1 vssd1 vccd1 vccd1 _20277_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23065_ _14883_/C input8/X _23073_/S vssd1 vssd1 vccd1 vccd1 _23066_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_47 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14322__C _15253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22016_ _22548_/A _22130_/A _22136_/A _22276_/A vssd1 vssd1 vccd1 vccd1 _22016_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15806__A2 _15621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17633__C _18016_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11981_ _23390_/Q vssd1 vssd1 vccd1 vccd1 _18468_/A sky130_fd_sc_hd__buf_2
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1029 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13235__A _13659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ _13720_/A _13720_/B _13720_/C _13720_/D vssd1 vssd1 vccd1 vccd1 _13720_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22918_ _12875_/B input38/X _22918_/S vssd1 vssd1 vccd1 vccd1 _22919_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22548__A _22548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13651_ _13632_/X _13630_/Y _22553_/C _22226_/C vssd1 vssd1 vccd1 vccd1 _13651_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22849_ _22849_/A _22849_/B vssd1 vssd1 vccd1 vccd1 _22849_/X sky130_fd_sc_hd__xor2_4
XFILLER_140_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18508__B2 _12460_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ _13052_/C vssd1 vssd1 vccd1 vccd1 _12930_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16370_ _16370_/A vssd1 vssd1 vccd1 vccd1 _16370_/X sky130_fd_sc_hd__buf_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13736_/A _13582_/B _22553_/D _22566_/C vssd1 vssd1 vccd1 vccd1 _13756_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_185_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15321_/A _15321_/B vssd1 vssd1 vccd1 vccd1 _15321_/X sky130_fd_sc_hd__xor2_1
XFILLER_157_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _12203_/A _12203_/B _12203_/C _12532_/Y vssd1 vssd1 vccd1 vccd1 _12533_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_13_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18040_ _17798_/A _17790_/Y _17798_/C vssd1 vssd1 vccd1 vccd1 _18040_/Y sky130_fd_sc_hd__o21ai_1
X_15252_ _15263_/A _15254_/C _15254_/A _15419_/A vssd1 vssd1 vccd1 vccd1 _15303_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12464_ _16815_/B _11582_/A _11947_/C _16140_/A vssd1 vssd1 vccd1 vccd1 _12464_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__18480__B _20320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14203_ _14203_/A _14203_/B vssd1 vssd1 vccd1 vccd1 _14793_/C sky130_fd_sc_hd__nand2_1
XFILLER_172_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15183_ _14212_/X _15166_/Y _15181_/X vssd1 vssd1 vccd1 vccd1 _15249_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__19484__A2 _19480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ _12547_/B _12547_/A _12392_/X _12394_/X vssd1 vssd1 vccd1 vccd1 _12396_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__16281__A _16281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ _15001_/A _14026_/X _14107_/A _14110_/X _14112_/Y vssd1 vssd1 vccd1 vccd1
+ _14137_/B sky130_fd_sc_hd__o32a_1
XANTENNA__21291__A2 _20504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19991_ _19991_/A _19991_/B _19991_/C vssd1 vssd1 vccd1 vccd1 _19991_/Y sky130_fd_sc_hd__nand3_2
XFILLER_180_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17527__D _18059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18942_ _18942_/A _18942_/B vssd1 vssd1 vccd1 vccd1 _18944_/A sky130_fd_sc_hd__nand2_1
X_14065_ _14284_/A _14284_/B _14285_/B _14285_/C vssd1 vssd1 vccd1 vccd1 _14292_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12314__A _12508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13016_ _20620_/B vssd1 vssd1 vccd1 vccd1 _20628_/B sky130_fd_sc_hd__clkbuf_2
X_18873_ _18841_/A _18841_/B _18844_/C _18872_/B vssd1 vssd1 vccd1 vccd1 _18873_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17824_ _17682_/A _17682_/B _17538_/X _17527_/C vssd1 vssd1 vccd1 vccd1 _18139_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_94_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20888__D _21268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18001__A _20081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17755_ _17760_/A _17760_/B _17754_/Y vssd1 vssd1 vccd1 vccd1 _17876_/A sky130_fd_sc_hd__o21ai_1
X_14967_ _15004_/B _14884_/X _14885_/Y _14891_/Y vssd1 vssd1 vccd1 vccd1 _14967_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16706_ _16706_/A _16706_/B vssd1 vssd1 vccd1 vccd1 _16708_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13918_ _23354_/Q _23353_/Q vssd1 vssd1 vccd1 vccd1 _14193_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17686_ _17686_/A vssd1 vssd1 vccd1 vccd1 _17686_/X sky130_fd_sc_hd__clkbuf_2
X_14898_ _14898_/A vssd1 vssd1 vccd1 vccd1 _14968_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_63_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19425_ _19534_/C _19900_/A _19425_/C _19614_/A vssd1 vssd1 vccd1 vccd1 _19425_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16637_ _16637_/A _16637_/B _16637_/C vssd1 vssd1 vccd1 vccd1 _16649_/B sky130_fd_sc_hd__nand3_2
X_13849_ _22220_/C _13582_/B _13674_/A _13680_/D _13846_/Y vssd1 vssd1 vccd1 vccd1
+ _13849_/Y sky130_fd_sc_hd__a221oi_2
XANTENNA__16456__A _17259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19356_ _12378_/A _12378_/B _17435_/X _17434_/X _17567_/X vssd1 vssd1 vccd1 vccd1
+ _19361_/A sky130_fd_sc_hd__o221a_2
XANTENNA__12244__B1 _16458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16568_ _16433_/X _16757_/D _16572_/B vssd1 vssd1 vccd1 vccd1 _16570_/A sky130_fd_sc_hd__a21bo_1
XFILLER_148_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18307_ _18251_/A _18251_/B _18254_/Y vssd1 vssd1 vccd1 vccd1 _18307_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18093__D _18172_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15519_ _15483_/X _15493_/A _15515_/Y _15516_/X _15518_/X vssd1 vssd1 vccd1 vccd1
+ _15520_/B sky130_fd_sc_hd__o41a_1
X_19287_ _19278_/X _19283_/X _19286_/Y vssd1 vssd1 vccd1 vccd1 _19290_/A sky130_fd_sc_hd__o21ai_1
X_16499_ _16499_/A vssd1 vssd1 vccd1 vccd1 _16536_/B sky130_fd_sc_hd__buf_2
XFILLER_176_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18238_ _18322_/A _18239_/C _18239_/A vssd1 vssd1 vccd1 vccd1 _18240_/A sky130_fd_sc_hd__o21a_1
XFILLER_164_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18169_ _18169_/A _20151_/C _18218_/A _18172_/A vssd1 vssd1 vccd1 vccd1 _18170_/D
+ sky130_fd_sc_hd__nand4_2
XANTENNA__16191__A _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20200_ _20311_/A _20200_/B vssd1 vssd1 vccd1 vccd1 _20203_/A sky130_fd_sc_hd__or2_1
XFILLER_144_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21180_ _21037_/A _21279_/C _21174_/Y vssd1 vssd1 vccd1 vccd1 _21184_/B sky130_fd_sc_hd__o21ai_1
X_20131_ _12237_/X _20081_/D _20164_/B _20043_/A vssd1 vssd1 vccd1 vccd1 _20131_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_131_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15238__C _15238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20062_ _20151_/A _20062_/B _20062_/C _20133_/B vssd1 vssd1 vccd1 vccd1 _20066_/C
+ sky130_fd_sc_hd__nand4_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17789__A2 _16523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18986__A1 _12051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15254__B _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18846__A _18846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20964_ _20969_/A _12648_/X _20959_/X _20960_/Y _20963_/Y vssd1 vssd1 vccd1 vccd1
+ _21101_/B sky130_fd_sc_hd__o221ai_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22368__A _22564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17410__A1 _16684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22703_ _22703_/A _22830_/D vssd1 vssd1 vccd1 vccd1 _22703_/Y sky130_fd_sc_hd__nor2_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_718 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12894__A _12899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20895_ _21047_/B _23299_/Q vssd1 vssd1 vccd1 vccd1 _20901_/C sky130_fd_sc_hd__nand2_1
XFILLER_110_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22634_ _22757_/B vssd1 vssd1 vccd1 vccd1 _22830_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1012 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22565_ _22650_/A _22563_/Y _22564_/X vssd1 vssd1 vccd1 vccd1 _22565_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_194_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17713__A2 _17635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21516_ _21517_/A _21517_/B vssd1 vssd1 vccd1 vccd1 _21516_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_1018 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22496_ _22496_/A _22496_/B _22545_/B _22544_/A vssd1 vssd1 vccd1 vccd1 _22501_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21447_ _21500_/A vssd1 vssd1 vccd1 vccd1 _21668_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20335__B _20363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18674__B1 _12214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12180_ _11926_/A _12281_/A _11935_/X _12171_/Y _12177_/Y vssd1 vssd1 vccd1 vccd1
+ _12181_/C sky130_fd_sc_hd__o221ai_4
XFILLER_107_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21378_ _21378_/A _21378_/B _21378_/C vssd1 vssd1 vccd1 vccd1 _21383_/B sky130_fd_sc_hd__nand3_1
XFILLER_119_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23117_ _11604_/X input18/X _23123_/S vssd1 vssd1 vccd1 vccd1 _23118_/A sky130_fd_sc_hd__mux2_1
X_20329_ _20329_/A _20329_/B vssd1 vssd1 vccd1 vccd1 _20376_/B sky130_fd_sc_hd__nor2_1
XFILLER_150_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23048_ _23048_/A vssd1 vssd1 vccd1 vccd1 _23352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12171__C1 _16122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12710__A1 _12709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18977__A1 _11864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18977__B2 _19504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15870_ _16526_/B vssd1 vssd1 vccd1 vccd1 _16549_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_77_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12788__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input22_A wb_dat_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ _14821_/A _14821_/B _14821_/C vssd1 vssd1 vccd1 vccd1 _14822_/B sky130_fd_sc_hd__nand3_1
XFILLER_36_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _17353_/Y _17357_/Y _17700_/B vssd1 vssd1 vccd1 vccd1 _17540_/X sky130_fd_sc_hd__o21a_1
X_14752_ _14752_/A _14886_/B _14752_/C vssd1 vssd1 vccd1 vccd1 _14756_/B sky130_fd_sc_hd__nand3_4
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _16860_/C vssd1 vssd1 vccd1 vccd1 _18506_/A sky130_fd_sc_hd__buf_2
XFILLER_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21733__B1 _13797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _13736_/A _22388_/B _13705_/C _13720_/A vssd1 vssd1 vccd1 vccd1 _13711_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _17463_/Y _17471_/B _17471_/C vssd1 vssd1 vccd1 vccd1 _17480_/A sky130_fd_sc_hd__nand3b_1
XFILLER_189_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14683_ _23371_/Q _14667_/X _14682_/X vssd1 vssd1 vccd1 vccd1 _14683_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11895_ _11788_/A _17149_/A _12343_/A _11803_/X _11880_/X vssd1 vssd1 vccd1 vccd1
+ _11902_/A sky130_fd_sc_hd__a32o_2
X_19210_ _19210_/A _19649_/A vssd1 vssd1 vccd1 vccd1 _19210_/Y sky130_fd_sc_hd__nor2_1
X_16422_ _16474_/B _16422_/B vssd1 vssd1 vccd1 vccd1 _16422_/Y sky130_fd_sc_hd__nor2_1
X_13634_ _13634_/A _13634_/B _21925_/B vssd1 vssd1 vccd1 vccd1 _13634_/X sky130_fd_sc_hd__and3_2
XANTENNA__15963__A1 _15862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19154__A1 _16054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19154__B2 _19504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19141_ _19141_/A _19141_/B vssd1 vssd1 vccd1 vccd1 _19141_/Y sky130_fd_sc_hd__nand2_1
X_16353_ _16343_/A _16575_/B _16576_/B vssd1 vssd1 vccd1 vccd1 _16435_/A sky130_fd_sc_hd__a21o_1
XFILLER_13_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13565_ _13720_/A _13720_/B vssd1 vssd1 vccd1 vccd1 _13569_/A sky130_fd_sc_hd__nand2_1
XFILLER_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15304_ _15358_/A _14990_/A _14990_/B _15301_/A _15415_/A vssd1 vssd1 vccd1 vccd1
+ _15308_/A sky130_fd_sc_hd__a32o_1
X_19072_ _18931_/A _18931_/B _18882_/B vssd1 vssd1 vccd1 vccd1 _19072_/Y sky130_fd_sc_hd__a21oi_1
X_12516_ _18756_/A vssd1 vssd1 vccd1 vccd1 _19364_/C sky130_fd_sc_hd__buf_4
XFILLER_160_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16284_ _15599_/X _15921_/B _15713_/C vssd1 vssd1 vccd1 vccd1 _16284_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13496_ _13498_/A _13498_/B _13495_/X vssd1 vssd1 vccd1 vccd1 _13496_/X sky130_fd_sc_hd__a21o_1
X_18023_ _18028_/A _18028_/B vssd1 vssd1 vccd1 vccd1 _18026_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15235_ _15001_/X _15171_/Y _15375_/A _15234_/Y vssd1 vssd1 vccd1 vccd1 _15237_/A
+ sky130_fd_sc_hd__o31a_1
X_12447_ _18511_/A _12422_/D _12446_/Y vssd1 vssd1 vccd1 vccd1 _12447_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output90_A _23264_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15166_ _15319_/C _15305_/A vssd1 vssd1 vccd1 vccd1 _15166_/Y sky130_fd_sc_hd__nand2_1
X_12378_ _12378_/A _12378_/B _16500_/D vssd1 vssd1 vccd1 vccd1 _12378_/X sky130_fd_sc_hd__or3_1
XFILLER_99_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _14120_/A _14120_/B _14261_/A vssd1 vssd1 vccd1 vccd1 _14174_/A sky130_fd_sc_hd__nand3_1
X_19974_ _19980_/C _20058_/A _19973_/X vssd1 vssd1 vccd1 vccd1 _19974_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__19209__A2 _17408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__A _18941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15097_ _15099_/A _15095_/X _15096_/Y _15000_/B vssd1 vssd1 vccd1 vccd1 _15097_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_125_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18925_ _18925_/A _18925_/B _23542_/Q vssd1 vssd1 vccd1 vccd1 _19288_/C sky130_fd_sc_hd__nand3_1
XANTENNA__21357__A _21358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14048_ _14068_/A _14069_/A _14429_/A vssd1 vssd1 vccd1 vccd1 _14054_/B sky130_fd_sc_hd__nand3_1
XANTENNA__20899__C _21174_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12979__A _12979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18856_ _18856_/A vssd1 vssd1 vccd1 vccd1 _18958_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17640__A1 _17410_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17807_ _17558_/X _17806_/Y _17805_/A _17805_/B vssd1 vssd1 vccd1 vccd1 _17807_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18787_ _18972_/B _18972_/C vssd1 vssd1 vccd1 vccd1 _19184_/A sky130_fd_sc_hd__nand2_4
X_15999_ _15999_/A _15999_/B _15999_/C vssd1 vssd1 vccd1 vccd1 _16010_/A sky130_fd_sc_hd__nand3_1
XFILLER_94_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17738_ _17575_/A _17734_/Y _17840_/B _17840_/A vssd1 vssd1 vccd1 vccd1 _17750_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__12465__B1 _12464_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2_0_bq_clk_i_A clkbuf_4_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17669_ _17670_/A _17670_/B _17670_/C _17668_/Y vssd1 vssd1 vccd1 vccd1 _17669_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_51_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19408_ _19408_/A _19420_/A vssd1 vssd1 vccd1 vccd1 _19413_/A sky130_fd_sc_hd__nand2_1
XFILLER_195_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20680_ _20672_/X _20520_/Y _20678_/Y _20679_/Y vssd1 vssd1 vccd1 vccd1 _20680_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19339_ _19340_/A _19341_/A _19339_/C vssd1 vssd1 vccd1 vccd1 _19339_/X sky130_fd_sc_hd__and3_1
XFILLER_176_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22350_ _21854_/A _21854_/B _22247_/Y _22348_/Y _22349_/Y vssd1 vssd1 vccd1 vccd1
+ _22351_/B sky130_fd_sc_hd__o221ai_1
XFILLER_149_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16903__B1 _16365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21301_ _21192_/Y _21292_/Y _21356_/A _21061_/X vssd1 vssd1 vccd1 vccd1 _21301_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13178__D1 _13181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11991__A2 _12121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22281_ _13465_/X _22059_/X _22283_/A vssd1 vssd1 vccd1 vccd1 _22281_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21232_ _21232_/A _21232_/B _21232_/C vssd1 vssd1 vccd1 vccd1 _21232_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__18656__B1 _20046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_675 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16131__A1 _16119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21163_ _21163_/A _21163_/B vssd1 vssd1 vccd1 vccd1 _21163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20114_ _20184_/A _20184_/B _20185_/A vssd1 vssd1 vccd1 vccd1 _20114_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_104_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21094_ _21057_/A _21057_/B _20941_/Y _20940_/X vssd1 vssd1 vccd1 vccd1 _21094_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13496__A2 _13498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18279__C _19900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20045_ _18476_/X _18484_/X _17414_/B _17414_/A _20320_/C vssd1 vssd1 vccd1 vccd1
+ _20045_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22755__A2 _22392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_88 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22507__A2 _13599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21996_ _22510_/A _22363_/A _22510_/C vssd1 vssd1 vccd1 vccd1 _21996_/Y sky130_fd_sc_hd__nand3_2
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _20947_/A _20947_/B vssd1 vssd1 vccd1 vccd1 _20948_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11680_ _11724_/A vssd1 vssd1 vccd1 vccd1 _12105_/C sky130_fd_sc_hd__clkbuf_4
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20878_ _20878_/A _20878_/B _23562_/Q vssd1 vssd1 vccd1 vccd1 _21030_/B sky130_fd_sc_hd__nand3_1
XFILLER_121_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22617_ _22617_/A vssd1 vssd1 vccd1 vccd1 _22858_/A sky130_fd_sc_hd__clkbuf_2
X_23597_ _23598_/CLK _23597_/D vssd1 vssd1 vccd1 vccd1 _23597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13350_ _23472_/Q vssd1 vssd1 vccd1 vccd1 _13416_/A sky130_fd_sc_hd__inv_2
X_22548_ _22548_/A _22677_/A _22548_/C _22667_/D vssd1 vssd1 vccd1 vccd1 _22549_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_195_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ _12391_/B _12251_/B _12393_/B _12393_/A vssd1 vssd1 vccd1 vccd1 _12303_/B
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__22264__C _22663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ _13766_/B vssd1 vssd1 vccd1 vccd1 _13634_/B sky130_fd_sc_hd__clkbuf_1
X_22479_ _22479_/A _22479_/B _22637_/C _22636_/C vssd1 vssd1 vccd1 vccd1 _22479_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_120_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15020_ _15075_/A _15081_/A _15020_/C _15265_/A vssd1 vssd1 vccd1 vccd1 _15081_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_182_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12232_ _12203_/Y _12220_/Y _12231_/Y vssd1 vssd1 vccd1 vccd1 _12232_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22561__A _22637_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _12159_/X _12160_/Y _12161_/Y _12162_/Y vssd1 vssd1 vccd1 vccd1 _12199_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_150_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22280__B _22280_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16673__A2 _16662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20081__A _20081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12094_ _23391_/Q vssd1 vssd1 vccd1 vccd1 _12100_/B sky130_fd_sc_hd__buf_2
X_16971_ _16725_/A _16737_/A _16721_/Y vssd1 vssd1 vccd1 vccd1 _16971_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18710_ _18902_/A vssd1 vssd1 vccd1 vccd1 _18914_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15922_ _15922_/A vssd1 vssd1 vccd1 vccd1 _15936_/A sky130_fd_sc_hd__buf_2
X_19690_ _19740_/B vssd1 vssd1 vccd1 vccd1 _19880_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17083__C1 _17077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18641_ _12311_/A _19670_/B _18639_/A vssd1 vssd1 vccd1 vccd1 _18647_/A sky130_fd_sc_hd__o21ai_2
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _15852_/X _15843_/A _15759_/X _15754_/X vssd1 vssd1 vccd1 vccd1 _15859_/A
+ sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__12949__D _20966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804_ _14207_/Y _14212_/X _14800_/A _14802_/Y _14803_/Y vssd1 vssd1 vccd1 vccd1
+ _14805_/B sky130_fd_sc_hd__o221ai_4
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18572_ _12542_/A _18437_/D _12542_/B _12398_/C _12543_/Y vssd1 vssd1 vccd1 vccd1
+ _18572_/X sky130_fd_sc_hd__a311o_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12996_ _20907_/A _20906_/A _20908_/A vssd1 vssd1 vccd1 vccd1 _21061_/A sky130_fd_sc_hd__o21ai_4
X_15784_ _15908_/A _15908_/B _15721_/X _15719_/B vssd1 vssd1 vccd1 vccd1 _15785_/C
+ sky130_fd_sc_hd__o211ai_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _17523_/A _17523_/B vssd1 vssd1 vccd1 vccd1 _17524_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11947_ _11947_/A _16140_/A _11947_/C vssd1 vssd1 vccd1 vccd1 _11948_/A sky130_fd_sc_hd__and3_1
X_14735_ _14735_/A vssd1 vssd1 vccd1 vccd1 _16749_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _19543_/B _17454_/B vssd1 vssd1 vccd1 vccd1 _17454_/Y sky130_fd_sc_hd__nand2_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _23399_/Q _14640_/X _14647_/X _23431_/Q _14665_/X vssd1 vssd1 vccd1 vccd1
+ _14666_/X sky130_fd_sc_hd__a221o_1
XANTENNA__14739__A2 _16749_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ _12262_/B vssd1 vssd1 vccd1 vccd1 _16462_/B sky130_fd_sc_hd__buf_4
X_16405_ _16405_/A _16405_/B vssd1 vssd1 vccd1 vccd1 _16407_/B sky130_fd_sc_hd__nand2_1
X_13617_ _13348_/X _13366_/Y _13620_/C vssd1 vssd1 vccd1 vccd1 _13816_/A sky130_fd_sc_hd__a21oi_4
X_17385_ _17362_/C _17362_/A _17362_/B vssd1 vssd1 vccd1 vccd1 _17385_/Y sky130_fd_sc_hd__a21oi_1
X_14597_ _15664_/C _14516_/X _14594_/X _14596_/X vssd1 vssd1 vccd1 vccd1 _14597_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12039__A _15682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19124_ _19530_/A _17586_/A _17587_/A _19121_/X _19123_/Y vssd1 vssd1 vccd1 vccd1
+ _19125_/C sky130_fd_sc_hd__a32o_1
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16336_ _16475_/B _16418_/A vssd1 vssd1 vccd1 vccd1 _16336_/X sky130_fd_sc_hd__and2_1
X_13548_ _13547_/X _21815_/B _21815_/C _13525_/C _13544_/B vssd1 vssd1 vccd1 vccd1
+ _13548_/X sky130_fd_sc_hd__o41a_1
XFILLER_185_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11973__A2 _11972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16897__C1 _15937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11878__A _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19055_ _19055_/A _19055_/B _19055_/C vssd1 vssd1 vccd1 vccd1 _19058_/B sky130_fd_sc_hd__nand3_1
X_16267_ _15949_/X _16004_/X _16260_/Y _16261_/Y vssd1 vssd1 vccd1 vccd1 _16586_/A
+ sky130_fd_sc_hd__o22ai_1
X_13479_ _13701_/A _22035_/C _13701_/C vssd1 vssd1 vccd1 vccd1 _13479_/X sky130_fd_sc_hd__and3_1
XFILLER_195_1016 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18006_ _17899_/B _17712_/B _17712_/A _20081_/A _18211_/D vssd1 vssd1 vccd1 vccd1
+ _18006_/X sky130_fd_sc_hd__a311o_1
XANTENNA__16172__C _17235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15218_ _15218_/A _15218_/B vssd1 vssd1 vccd1 vccd1 _15219_/B sky130_fd_sc_hd__xnor2_4
XFILLER_127_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18638__B1 _18476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16198_ _17631_/A _17148_/A _16198_/C vssd1 vssd1 vccd1 vccd1 _16198_/X sky130_fd_sc_hd__and3_1
XFILLER_160_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20445__B1 _20031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17565__A _17565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15149_ _15220_/A _15220_/B _15220_/C _15439_/C vssd1 vssd1 vccd1 vccd1 _15219_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_141_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19957_ _19957_/A _20142_/B _20371_/C _19957_/D vssd1 vssd1 vccd1 vccd1 _19957_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_142_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18908_ _19091_/B _19091_/C vssd1 vssd1 vccd1 vccd1 _18910_/B sky130_fd_sc_hd__nand2_1
XANTENNA__15085__A _15488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19888_ _19888_/A _19888_/B _20003_/A _19888_/D vssd1 vssd1 vccd1 vccd1 _19889_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_132_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18839_ _18841_/A _18841_/B _18844_/C _18872_/B vssd1 vssd1 vccd1 vccd1 _18839_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13317__B _13766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21815__A _22236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14427__B2 _15094_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21850_ _21850_/A _21850_/B vssd1 vssd1 vccd1 vccd1 _21972_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20801_ _21036_/A _21036_/B _20801_/C vssd1 vssd1 vccd1 vccd1 _20814_/A sky130_fd_sc_hd__nand3_1
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21781_ _21780_/Y _13812_/A _13799_/A _13819_/Y vssd1 vssd1 vccd1 vccd1 _21782_/C
+ sky130_fd_sc_hd__a22oi_4
XANTENNA__17450__D _20317_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23520_ _23566_/CLK _23520_/D vssd1 vssd1 vccd1 vccd1 _23520_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_169_818 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20732_ _20715_/A _20715_/B _20715_/C _20718_/A vssd1 vssd1 vccd1 vccd1 _20732_/Y
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__19118__A1 _12246_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13938__B1 _13911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16066__D _19670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23451_ _23462_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _23451_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13052__B _23453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20663_ _21277_/A _21065_/A _20663_/C _20663_/D vssd1 vssd1 vccd1 vccd1 _20663_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19669__A2 _18455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22402_ _22402_/A vssd1 vssd1 vccd1 vccd1 _22516_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23382_ _23385_/CLK _23382_/D vssd1 vssd1 vccd1 vccd1 _23382_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_164_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17459__B _17605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20594_ _20594_/A _20594_/B vssd1 vssd1 vccd1 vccd1 _20594_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22333_ _22333_/A _22333_/B _22333_/C vssd1 vssd1 vccd1 vccd1 _22357_/B sky130_fd_sc_hd__nand3_2
XFILLER_87_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22264_ _22261_/Y _22264_/B _22663_/D vssd1 vssd1 vccd1 vccd1 _22264_/Y sky130_fd_sc_hd__nand3b_1
XANTENNA__14902__A2 _14050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19674__B _19674_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23263__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21215_ _21215_/A _21319_/B _21215_/C vssd1 vssd1 vccd1 vccd1 _21216_/A sky130_fd_sc_hd__nand3_1
X_22195_ _22197_/A _22197_/B _22214_/C vssd1 vssd1 vccd1 vccd1 _22195_/Y sky130_fd_sc_hd__nand3_2
XFILLER_133_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21146_ _21144_/Y _21146_/B vssd1 vssd1 vccd1 vccd1 _21147_/B sky130_fd_sc_hd__and2b_1
XFILLER_120_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22189__B1 _23331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21077_ _20962_/Y _21194_/A _21302_/A _21271_/B _21063_/Y vssd1 vssd1 vccd1 vccd1
+ _21163_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_58_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20028_ _20032_/A _20032_/B _20306_/A vssd1 vssd1 vccd1 vccd1 _20028_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12850_ _12850_/A _12850_/B vssd1 vssd1 vccd1 vccd1 _12851_/A sky130_fd_sc_hd__nand2_1
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19357__A1 _17742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _11896_/B vssd1 vssd1 vccd1 vccd1 _11801_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _13166_/A vssd1 vssd1 vccd1 vccd1 _13151_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ _21979_/A _21979_/B vssd1 vssd1 vccd1 vccd1 _23561_/D sky130_fd_sc_hd__xnor2_4
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ _14551_/A vssd1 vssd1 vccd1 vccd1 _14520_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11732_ _23584_/Q _11644_/C _11808_/A vssd1 vssd1 vccd1 vccd1 _11860_/A sky130_fd_sc_hd__o21ai_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11652__A1 _16802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16040__B1 _12018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14975_/C vssd1 vssd1 vccd1 vccd1 _15310_/B sky130_fd_sc_hd__buf_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11663_ _12024_/A vssd1 vssd1 vccd1 vccd1 _19363_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_186_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13402_ _21882_/A vssd1 vssd1 vccd1 vccd1 _21793_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17170_ _17350_/A _17170_/B _17170_/C vssd1 vssd1 vccd1 vccd1 _17170_/X sky130_fd_sc_hd__and3_1
XFILLER_41_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14382_ _14791_/C vssd1 vssd1 vccd1 vccd1 _14806_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11594_ _11971_/A _11972_/A vssd1 vssd1 vccd1 vccd1 _12474_/A sky130_fd_sc_hd__nand2_2
X_16121_ _16860_/A _17098_/C _16840_/A _16634_/C vssd1 vssd1 vccd1 vccd1 _16121_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_127_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13333_ _21739_/A vssd1 vssd1 vccd1 vccd1 _21902_/C sky130_fd_sc_hd__buf_2
XFILLER_155_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16052_ _16094_/B vssd1 vssd1 vccd1 vccd1 _16052_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13264_ _13483_/B _13264_/B _13264_/C vssd1 vssd1 vccd1 vccd1 _13766_/B sky130_fd_sc_hd__nand3_4
XFILLER_109_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15003_ _14181_/X _14999_/Y _15000_/Y _15002_/X vssd1 vssd1 vccd1 vccd1 _15004_/D
+ sky130_fd_sc_hd__o22ai_2
XFILLER_182_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12215_ _12107_/X _12110_/Y _12238_/A _12214_/X vssd1 vssd1 vccd1 vccd1 _12216_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_6_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13195_ _13189_/X _13191_/X _13192_/X _13193_/Y _13194_/Y vssd1 vssd1 vccd1 vccd1
+ _13195_/X sky130_fd_sc_hd__o2111a_1
XFILLER_68_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23537__D _23537_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19811_ _19811_/A _20055_/A _20055_/B vssd1 vssd1 vccd1 vccd1 _19811_/Y sky130_fd_sc_hd__nand3_1
XFILLER_2_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12146_ _16802_/A vssd1 vssd1 vccd1 vccd1 _12146_/X sky130_fd_sc_hd__buf_2
XFILLER_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19742_ _19742_/A _19742_/B _19742_/C vssd1 vssd1 vccd1 vccd1 _19743_/A sky130_fd_sc_hd__nand3_1
XFILLER_96_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12077_ _19811_/A vssd1 vssd1 vccd1 vccd1 _20142_/D sky130_fd_sc_hd__clkbuf_4
X_16954_ _16888_/A _16888_/B _16888_/C vssd1 vssd1 vccd1 vccd1 _16954_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15905_ _15905_/A vssd1 vssd1 vccd1 vccd1 _16055_/A sky130_fd_sc_hd__buf_2
X_19673_ _19675_/A _19667_/D _19667_/A _19665_/A vssd1 vssd1 vccd1 vccd1 _19673_/Y
+ sky130_fd_sc_hd__a22oi_4
X_16885_ _16885_/A vssd1 vssd1 vccd1 vccd1 _16894_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18624_ _18620_/Y _18931_/B _18622_/X _18623_/X vssd1 vssd1 vccd1 vccd1 _18712_/A
+ sky130_fd_sc_hd__o211ai_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _15836_/A _15836_/B _15836_/C vssd1 vssd1 vccd1 vccd1 _16073_/B sky130_fd_sc_hd__nand3_4
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18555_ _18555_/A _18555_/B _18555_/C vssd1 vssd1 vccd1 vccd1 _18560_/A sky130_fd_sc_hd__nand3_1
XFILLER_18_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _16808_/A _16800_/A _16619_/A vssd1 vssd1 vccd1 vccd1 _16126_/A sky130_fd_sc_hd__nand3_4
X_12979_ _12979_/A vssd1 vssd1 vccd1 vccd1 _13186_/C sky130_fd_sc_hd__clkbuf_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17506_ _17506_/A vssd1 vssd1 vccd1 vccd1 _18211_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__16167__C _16167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14718_ _23349_/Q _14531_/A _14546_/A _23317_/Q _14657_/A vssd1 vssd1 vccd1 vccd1
+ _14718_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18486_ _18486_/A vssd1 vssd1 vccd1 vccd1 _19491_/A sky130_fd_sc_hd__buf_2
XFILLER_178_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22466__A _22566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15698_ _15698_/A _15698_/B vssd1 vssd1 vccd1 vccd1 _15831_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17437_ _17571_/A vssd1 vssd1 vccd1 vccd1 _17437_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12992__A _23457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14649_ _15735_/B vssd1 vssd1 vccd1 vccd1 _15645_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16464__A _16464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17368_ _17036_/X _17195_/Y _17196_/Y vssd1 vssd1 vccd1 vccd1 _17369_/D sky130_fd_sc_hd__o21ai_1
XFILLER_158_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19107_ _19294_/B _19107_/B _19107_/C vssd1 vssd1 vccd1 vccd1 _19284_/C sky130_fd_sc_hd__nand3_1
XFILLER_118_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16319_ _16319_/A vssd1 vssd1 vccd1 vccd1 _16382_/A sky130_fd_sc_hd__buf_2
XFILLER_119_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16334__A1 _16066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17299_ _17299_/A _17299_/B _17299_/C vssd1 vssd1 vccd1 vccd1 _17337_/B sky130_fd_sc_hd__nand3_2
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19038_ _19148_/C _19148_/A _19148_/B vssd1 vssd1 vccd1 vccd1 _19038_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19494__B _19969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18087__B2 _20215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23080__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21000_ _21000_/A _21000_/B vssd1 vssd1 vccd1 vccd1 _21130_/A sky130_fd_sc_hd__and2_1
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15527__B _15527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21545__A _21545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22951_ _23310_/Q input23/X _22951_/S vssd1 vssd1 vccd1 vccd1 _22952_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20051__D1 _20215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13871__A2 _13867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21933__A3 _22045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21902_ _22028_/A _21902_/B _21902_/C vssd1 vssd1 vccd1 vccd1 _22031_/A sky130_fd_sc_hd__nand3_1
XFILLER_28_437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19015__A _19043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22882_ _22872_/B _23284_/Q vssd1 vssd1 vccd1 vccd1 _22882_/X sky130_fd_sc_hd__and2b_1
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12886__B _23452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21833_ _22754_/A _21815_/B _21815_/C _13848_/B _21832_/Y vssd1 vssd1 vccd1 vccd1
+ _21833_/X sky130_fd_sc_hd__o41a_1
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18276__D _18330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18011__A1 _18016_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21764_ _21783_/B _21764_/B _21764_/C vssd1 vssd1 vccd1 vccd1 _21764_/X sky130_fd_sc_hd__and3_1
XFILLER_196_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23503_ _23510_/CLK _23503_/D vssd1 vssd1 vccd1 vccd1 _23503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20715_ _20715_/A _20715_/B _20715_/C _20718_/A vssd1 vssd1 vccd1 vccd1 _20716_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_52_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21695_ _21695_/A _21695_/B vssd1 vssd1 vccd1 vccd1 _21704_/D sky130_fd_sc_hd__nor2_2
XFILLER_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19388__C _19568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23434_ _23434_/CLK _23434_/D vssd1 vssd1 vccd1 vccd1 _23434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20646_ _20921_/A _20921_/B _20681_/C vssd1 vssd1 vccd1 vccd1 _20646_/Y sky130_fd_sc_hd__nand3_2
XFILLER_177_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11937__A2 _11935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23365_ _23365_/CLK _23365_/D vssd1 vssd1 vccd1 vccd1 _23365_/Q sky130_fd_sc_hd__dfxtp_1
X_20577_ _20568_/Y _20575_/Y _20576_/Y vssd1 vssd1 vccd1 vccd1 _20577_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22316_ _22177_/Y _22195_/Y _22200_/Y _22215_/X vssd1 vssd1 vccd1 vccd1 _22316_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23296_ _23296_/CLK _23296_/D vssd1 vssd1 vccd1 vccd1 _23296_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_152_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23071__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22247_ _22117_/Y _22243_/Y _22246_/Y vssd1 vssd1 vccd1 vccd1 _22247_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__15718__A _15718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12898__B1 _12899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12000_ _11999_/B _18999_/C _11999_/A vssd1 vssd1 vccd1 vccd1 _12185_/A sky130_fd_sc_hd__a21oi_4
XFILLER_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22178_ _22211_/A _22211_/B _22061_/Y vssd1 vssd1 vccd1 vccd1 _22197_/B sky130_fd_sc_hd__o21ai_1
XFILLER_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14639__A1 _19156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14639__B2 _14631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20062__C _20062_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21129_ _21134_/C _21126_/Y _21127_/Y _21128_/Y vssd1 vssd1 vccd1 vccd1 _21129_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_78_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13951_ _13951_/A _13951_/B vssd1 vssd1 vccd1 vccd1 _14396_/A sky130_fd_sc_hd__nand2_2
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12902_ _12911_/A _12911_/B _12902_/C _12902_/D vssd1 vssd1 vccd1 vccd1 _12908_/B
+ sky130_fd_sc_hd__nand4_1
X_16670_ _17134_/C vssd1 vssd1 vccd1 vccd1 _17388_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13882_ _14377_/A vssd1 vssd1 vccd1 vccd1 _14469_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__21174__B _21174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ _15634_/C vssd1 vssd1 vccd1 vccd1 _15621_/X sky130_fd_sc_hd__clkbuf_4
X_12833_ _13115_/A _12833_/B _13115_/B _20962_/B vssd1 vssd1 vccd1 vccd1 _12835_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18538__C1 _18080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _18339_/A _18339_/B _18339_/C vssd1 vssd1 vccd1 vccd1 _18341_/B sky130_fd_sc_hd__a21o_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21902__B _21902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15552_ _15552_/A _15552_/B vssd1 vssd1 vccd1 vccd1 _23283_/D sky130_fd_sc_hd__xor2_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12792_/A vssd1 vssd1 vccd1 vccd1 _12765_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _16027_/B vssd1 vssd1 vccd1 vccd1 _19323_/A sky130_fd_sc_hd__buf_4
XFILLER_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14503_ _23414_/Q vssd1 vssd1 vccd1 vccd1 _15735_/C sky130_fd_sc_hd__buf_2
X_18271_ _20212_/D vssd1 vssd1 vccd1 vccd1 _20268_/D sky130_fd_sc_hd__clkbuf_2
X_15483_ _15508_/A _15511_/D _15483_/C vssd1 vssd1 vccd1 vccd1 _15483_/X sky130_fd_sc_hd__and3_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12695_/A vssd1 vssd1 vccd1 vccd1 _21271_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17222_ _17126_/A _17126_/B _17126_/C _17125_/B vssd1 vssd1 vccd1 vccd1 _17222_/Y
+ sky130_fd_sc_hd__a31oi_2
X_14434_ _14068_/X _14069_/X _14252_/D _14867_/C _14430_/D vssd1 vssd1 vccd1 vccd1
+ _14465_/D sky130_fd_sc_hd__a32o_1
X_11646_ _23587_/Q vssd1 vssd1 vccd1 vccd1 _11647_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_156_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 wb_dat_i[16] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17153_ _17156_/A _17359_/B _17161_/A vssd1 vssd1 vccd1 vccd1 _17220_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__16316__A1 _18461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 wb_dat_i[26] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_2
X_14365_ _14365_/A _14365_/B _14365_/C vssd1 vssd1 vccd1 vccd1 _14422_/B sky130_fd_sc_hd__nand3_1
XFILLER_122_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11577_ _12497_/A _12071_/A _16815_/B vssd1 vssd1 vccd1 vccd1 _11577_/Y sky130_fd_sc_hd__a21oi_1
Xinput36 wb_dat_i[7] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_4
XFILLER_10_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16316__B2 _16194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput47 x[4] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14327__B1 _14181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13316_ _21764_/C vssd1 vssd1 vccd1 vccd1 _22392_/C sky130_fd_sc_hd__clkbuf_4
X_16104_ _16104_/A _16297_/A _16297_/B vssd1 vssd1 vccd1 vccd1 _16340_/C sky130_fd_sc_hd__nand3_1
X_17084_ _17089_/A _17089_/B _17082_/X _17083_/X vssd1 vssd1 vccd1 vccd1 _17126_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_128_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16867__A2 _17605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14296_ _14936_/B vssd1 vssd1 vccd1 vccd1 _14834_/A sky130_fd_sc_hd__buf_2
XFILLER_155_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23062__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13247_ _13247_/A _22365_/C _13523_/A _13247_/D vssd1 vssd1 vccd1 vccd1 _13656_/B
+ sky130_fd_sc_hd__nand4_1
X_16035_ _16032_/X _16033_/X _16308_/C _16308_/D vssd1 vssd1 vccd1 vccd1 _16035_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19266__B1 _18373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17546__C _17546_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13178_ _13176_/X _13177_/X _13181_/A _13186_/C _13181_/B vssd1 vssd1 vccd1 vccd1
+ _13178_/X sky130_fd_sc_hd__o2111a_1
XFILLER_124_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12129_ _12399_/A _12399_/C vssd1 vssd1 vccd1 vccd1 _12129_/Y sky130_fd_sc_hd__nand2_1
X_17986_ _18172_/A _17986_/B _18100_/A _17986_/D vssd1 vssd1 vccd1 vccd1 _17992_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12052__A _12052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19725_ _19725_/A _19725_/B _19725_/C vssd1 vssd1 vccd1 vccd1 _19893_/A sky130_fd_sc_hd__nand3_2
XFILLER_111_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16937_ _16932_/Y _16647_/B _16647_/C vssd1 vssd1 vccd1 vccd1 _16937_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_111_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17044__A2 _16447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19656_ _19656_/A _19656_/B vssd1 vssd1 vccd1 vccd1 _19855_/C sky130_fd_sc_hd__nor2_2
XFILLER_93_852 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16868_ _16592_/B _17095_/A _15991_/A _17107_/A _17226_/D vssd1 vssd1 vccd1 vccd1
+ _16870_/B sky130_fd_sc_hd__o2111ai_1
X_18607_ _18607_/A _18947_/B _18607_/C vssd1 vssd1 vccd1 vccd1 _18607_/X sky130_fd_sc_hd__and3_1
XFILLER_77_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15819_ _17066_/C vssd1 vssd1 vccd1 vccd1 _17259_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19587_ _19587_/A _19747_/A _19587_/C vssd1 vssd1 vccd1 vccd1 _19587_/X sky130_fd_sc_hd__and3_1
X_16799_ _16799_/A vssd1 vssd1 vccd1 vccd1 _17569_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14802__B2 _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18538_ _18536_/X _18537_/Y _18534_/Y _18080_/A _12508_/D vssd1 vssd1 vccd1 vccd1
+ _18540_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_602 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_957 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16555__A1 _16531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18469_ _18649_/A _18469_/B _18469_/C _18469_/D vssd1 vssd1 vccd1 vccd1 _18470_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__16194__A _16194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20500_ _20496_/X _21431_/B _12696_/A _20645_/C _12695_/A vssd1 vssd1 vccd1 vccd1
+ _20501_/A sky130_fd_sc_hd__a32oi_2
XFILLER_166_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21480_ _21346_/X _21423_/Y _21528_/B _21576_/A vssd1 vssd1 vccd1 vccd1 _21484_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_140_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20431_ _20409_/A _20431_/B _20431_/C vssd1 vssd1 vccd1 vccd1 _20446_/B sky130_fd_sc_hd__nand3b_2
XFILLER_140_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23150_ _23398_/Q input14/X _23156_/S vssd1 vssd1 vccd1 vccd1 _23151_/A sky130_fd_sc_hd__mux2_1
X_20362_ _20031_/X _20301_/Y _20341_/X _20361_/Y vssd1 vssd1 vccd1 vccd1 _20362_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_107_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22101_ _22102_/A _22240_/B _22102_/C vssd1 vssd1 vccd1 vccd1 _22101_/Y sky130_fd_sc_hd__a21oi_1
X_23081_ _23081_/A vssd1 vssd1 vccd1 vccd1 _23367_/D sky130_fd_sc_hd__clkbuf_1
X_20293_ _20290_/B _20243_/B _20242_/B _20291_/X _20337_/A vssd1 vssd1 vccd1 vccd1
+ _20293_/X sky130_fd_sc_hd__a32o_2
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_751 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22032_ _22381_/A _22381_/B _13810_/B _22030_/Y _22562_/C vssd1 vssd1 vccd1 vccd1
+ _22032_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_88_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18849__A _19017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17753__A _17753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22934_ _23302_/Q input14/X _22940_/S vssd1 vssd1 vccd1 vccd1 _22935_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16088__B _16423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23451__CLK _23462_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22865_ _22865_/A _22865_/B vssd1 vssd1 vccd1 vccd1 _22868_/A sky130_fd_sc_hd__nor2_2
XFILLER_189_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21816_ _13741_/B _13741_/C _22420_/A vssd1 vssd1 vccd1 vccd1 _21816_/X sky130_fd_sc_hd__a21o_1
XFILLER_169_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22796_ _22797_/C _22797_/A _22797_/B vssd1 vssd1 vccd1 vccd1 _22798_/A sky130_fd_sc_hd__o21a_1
XANTENNA__18535__A2 _17586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12280__A1 _11611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21747_ _22047_/B _13355_/A _21745_/B vssd1 vssd1 vccd1 vccd1 _21747_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_185_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17743__B1 _18778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16546__B2 _15731_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13521__A _13732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12480_ _12480_/A _12480_/B vssd1 vssd1 vccd1 vccd1 _12481_/B sky130_fd_sc_hd__nor2_1
X_21678_ _21616_/X _21617_/X _21665_/Y _21694_/A _21698_/B vssd1 vssd1 vccd1 vccd1
+ _21691_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_132_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23417_ _23428_/CLK _23417_/D vssd1 vssd1 vccd1 vccd1 _23417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20629_ _20475_/B _20783_/A _20793_/A vssd1 vssd1 vccd1 vccd1 _20632_/A sky130_fd_sc_hd__o21ai_1
XFILLER_138_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22553__B _22554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14150_ _13985_/X _14162_/B _14407_/A _14150_/D vssd1 vssd1 vccd1 vccd1 _14150_/Y
+ sky130_fd_sc_hd__nand4b_1
XFILLER_193_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23348_ _23349_/CLK _23348_/D vssd1 vssd1 vccd1 vccd1 _23348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13101_ _13088_/B _13101_/B _13101_/C vssd1 vssd1 vccd1 vccd1 _20464_/A sky130_fd_sc_hd__nand3b_4
XFILLER_153_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14081_ _14178_/B vssd1 vssd1 vccd1 vccd1 _15253_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23279_ _23518_/CLK _23279_/D vssd1 vssd1 vccd1 vccd1 _23279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _13001_/X _13029_/Y _13030_/Y _13031_/Y vssd1 vssd1 vccd1 vccd1 _13032_/X
+ sky130_fd_sc_hd__o211a_2
XANTENNA__21055__B1 _13122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input52_A x[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11695__B _23587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15809__B1 _17465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20802__B1 _13151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17840_ _17840_/A _17840_/B vssd1 vssd1 vccd1 vccd1 _17840_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17771_ _17585_/C _17769_/Y _17770_/Y _17609_/A vssd1 vssd1 vccd1 vccd1 _17771_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_121_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14983_ _14983_/A vssd1 vssd1 vccd1 vccd1 _15422_/A sky130_fd_sc_hd__clkbuf_2
X_19510_ _16526_/D _19868_/A _19307_/Y vssd1 vssd1 vccd1 vccd1 _19514_/A sky130_fd_sc_hd__a21oi_1
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16722_ _16722_/A _16722_/B _16722_/C vssd1 vssd1 vccd1 vccd1 _16950_/B sky130_fd_sc_hd__nand3_2
X_13934_ _23495_/Q vssd1 vssd1 vccd1 vccd1 _14774_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__12600__A _20782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19971__A1 _12509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_72 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19441_ _19297_/X _19298_/Y _19268_/X _19299_/Y _19440_/Y vssd1 vssd1 vccd1 vccd1
+ _19447_/A sky130_fd_sc_hd__o221ai_4
X_16653_ _16655_/B _16655_/C _16655_/D _16655_/A vssd1 vssd1 vccd1 vccd1 _16723_/A
+ sky130_fd_sc_hd__a22o_1
X_13865_ _21839_/A _21840_/A _13863_/Y _13864_/Y vssd1 vssd1 vccd1 vccd1 _21856_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15604_ _16658_/B vssd1 vssd1 vccd1 vccd1 _15604_/X sky130_fd_sc_hd__clkbuf_4
X_19372_ _12243_/X _17763_/A _19363_/Y _19540_/A _19365_/Y vssd1 vssd1 vccd1 vccd1
+ _19374_/B sky130_fd_sc_hd__o221ai_1
X_12816_ _12816_/A _12816_/B _12816_/C vssd1 vssd1 vccd1 vccd1 _12817_/B sky130_fd_sc_hd__nor3_1
XANTENNA_clkbuf_4_7_0_bq_clk_i_A clkbuf_4_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16584_ _16584_/A vssd1 vssd1 vccd1 vccd1 _16989_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13796_ _13796_/A _13796_/B _21909_/C vssd1 vssd1 vccd1 vccd1 _13797_/B sky130_fd_sc_hd__and3_1
XFILLER_31_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18323_ _18285_/A _18284_/A _18284_/B _18286_/B _18286_/A vssd1 vssd1 vccd1 vccd1
+ _18343_/B sky130_fd_sc_hd__o32ai_2
XFILLER_72_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15535_ _15102_/A _15102_/B _15488_/B vssd1 vssd1 vccd1 vccd1 _15536_/C sky130_fd_sc_hd__a21o_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16537__A1 _16749_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12747_ _23447_/Q vssd1 vssd1 vccd1 vccd1 _20681_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_188_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17734__B1 _20317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _18302_/A _18254_/B _18254_/C vssd1 vssd1 vccd1 vccd1 _18254_/Y sky130_fd_sc_hd__nand3_2
XFILLER_148_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15466_ _15466_/A vssd1 vssd1 vccd1 vccd1 _15471_/A sky130_fd_sc_hd__inv_2
X_12678_ _23291_/Q _12873_/C _12678_/C vssd1 vssd1 vccd1 vccd1 _12678_/Y sky130_fd_sc_hd__nor3_2
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14246__B _14246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18941__B _18941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17205_ _17196_/Y _17200_/Y _17203_/Y _17204_/Y vssd1 vssd1 vccd1 vccd1 _17365_/D
+ sky130_fd_sc_hd__a22oi_4
X_11629_ _12207_/A vssd1 vssd1 vccd1 vccd1 _11935_/A sky130_fd_sc_hd__buf_4
X_14417_ _14420_/A _14352_/B _14414_/A _14414_/B vssd1 vssd1 vccd1 vccd1 _14418_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12023__A1 _12021_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18185_ _18185_/A _18185_/B _18185_/C vssd1 vssd1 vccd1 vccd1 _18186_/B sky130_fd_sc_hd__nor3_1
XFILLER_175_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15397_ _15335_/B _15395_/Y _15396_/X vssd1 vssd1 vccd1 vccd1 _15397_/X sky130_fd_sc_hd__a21o_1
XFILLER_129_876 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17136_ _16902_/Y _17140_/A _16913_/B _16904_/Y vssd1 vssd1 vccd1 vccd1 _17151_/A
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_184_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14348_ _14358_/C _14358_/B _14346_/Y _14347_/X vssd1 vssd1 vccd1 vccd1 _14350_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_183_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12292__A1_N _11717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15358__A _15358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17067_ _17077_/A _17077_/B vssd1 vssd1 vccd1 vccd1 _17067_/X sky130_fd_sc_hd__and2_1
X_14279_ _14279_/A _14279_/B _14279_/C vssd1 vssd1 vccd1 vccd1 _14358_/C sky130_fd_sc_hd__nand3_2
XFILLER_171_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16018_ _16018_/A vssd1 vssd1 vccd1 vccd1 _16347_/B sky130_fd_sc_hd__clkbuf_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17265__A2 _12518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _18077_/A _18079_/A _20146_/A _17969_/D vssd1 vssd1 vccd1 vccd1 _18157_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13826__A2 _13456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22546__B1 _22754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19708_ _19708_/A _19708_/B vssd1 vssd1 vccd1 vccd1 _19710_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11837__A1 _11849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20980_ _20980_/A _20980_/B _20980_/C vssd1 vssd1 vccd1 vccd1 _20994_/C sky130_fd_sc_hd__nand3_1
XANTENNA__11837__B2 _12475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19639_ _19613_/Y _19638_/Y _19467_/A vssd1 vssd1 vccd1 vccd1 _19772_/A sky130_fd_sc_hd__o21ai_2
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20572__A2 _20726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22650_ _22650_/A _22650_/B _22713_/D _22712_/A vssd1 vssd1 vccd1 vccd1 _22650_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_198_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15984__C1 _16840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23460__D _23472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21601_ _21590_/A _21590_/B _21602_/B vssd1 vssd1 vccd1 vccd1 _21601_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19012__B _19012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22581_ _22469_/X _22567_/Y _22468_/X _22579_/Y _22573_/A vssd1 vssd1 vccd1 vccd1
+ _22581_/X sky130_fd_sc_hd__o2111a_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21532_ _21541_/C _21541_/A _23569_/Q vssd1 vssd1 vccd1 vccd1 _21540_/A sky130_fd_sc_hd__a21oi_1
XFILLER_194_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21463_ _21463_/A _21463_/B _21463_/C _21463_/D vssd1 vssd1 vccd1 vccd1 _21464_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13211__B1 _13210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15751__A2 _11921_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23202_ _15713_/C input36/X _23206_/S vssd1 vssd1 vccd1 vccd1 _23203_/A sky130_fd_sc_hd__mux2_1
X_20414_ _20414_/A _20414_/B vssd1 vssd1 vccd1 vccd1 _20452_/C sky130_fd_sc_hd__nand2_1
XFILLER_181_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21394_ _21311_/A _21328_/Y _21390_/X _21465_/B _21327_/C vssd1 vssd1 vccd1 vccd1
+ _21399_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_135_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_952 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23133_ _23133_/A vssd1 vssd1 vccd1 vccd1 _23390_/D sky130_fd_sc_hd__clkbuf_1
X_20345_ _20343_/Y _20344_/X _20384_/B _20340_/Y _20341_/A vssd1 vssd1 vccd1 vccd1
+ _20345_/X sky130_fd_sc_hd__o2111a_1
XFILLER_135_868 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23026__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16161__C1 _19811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12317__A2 _11749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23064_ _23110_/S vssd1 vssd1 vccd1 vccd1 _23073_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_68_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20276_ _20274_/A _20274_/B _20274_/C _20400_/A vssd1 vssd1 vccd1 vccd1 _20328_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_108_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22015_ _22130_/A _22136_/A _13470_/A _13410_/X vssd1 vssd1 vccd1 vccd1 _22015_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_68_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13278__B1 _13469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22001__A2 _21892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11980_ _11980_/A _11980_/B _18469_/B _18998_/C vssd1 vssd1 vccd1 vccd1 _11980_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_99_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_716 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22917_ _22917_/A vssd1 vssd1 vccd1 vccd1 _23294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15731__A _15731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13650_ _13650_/A vssd1 vssd1 vccd1 vccd1 _22226_/C sky130_fd_sc_hd__clkbuf_2
X_22848_ _22859_/A _22828_/Y _22858_/A vssd1 vssd1 vccd1 vccd1 _22848_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_72_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12601_/A _12601_/B _12601_/C vssd1 vssd1 vccd1 vccd1 _13052_/C sky130_fd_sc_hd__nand3_4
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _22278_/B vssd1 vssd1 vccd1 vccd1 _22553_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17136__A2_N _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22779_ _22828_/B vssd1 vssd1 vccd1 vccd1 _22780_/B sky130_fd_sc_hd__inv_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12532_ _12532_/A _12532_/B vssd1 vssd1 vccd1 vccd1 _12532_/Y sky130_fd_sc_hd__nor2_1
X_15320_ _15366_/A _15366_/C _15241_/Y _15422_/A vssd1 vssd1 vccd1 vccd1 _15321_/B
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_0_0_bq_clk_i clkbuf_4_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _23510_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_169_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22564__A _22564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12463_ _19017_/A _18600_/C _18756_/B _19017_/D vssd1 vssd1 vccd1 vccd1 _12463_/Y
+ sky130_fd_sc_hd__nand4_4
X_15251_ _15251_/A vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18480__C _19846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14202_ _14911_/A _14886_/A _14202_/C _15116_/B vssd1 vssd1 vccd1 vccd1 _14800_/B
+ sky130_fd_sc_hd__nand4_1
X_15182_ _14212_/X _15166_/Y _15250_/A _15187_/C _15181_/X vssd1 vssd1 vccd1 vccd1
+ _15185_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_153_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ _12251_/X _12393_/Y _12300_/C vssd1 vssd1 vccd1 vccd1 _12394_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16281__B _16281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ _14133_/A _14133_/B vssd1 vssd1 vccd1 vccd1 _14137_/A sky130_fd_sc_hd__nand2_1
XANTENNA__23017__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19990_ _19974_/Y _19977_/Y _19982_/Y _19986_/B vssd1 vssd1 vccd1 vccd1 _19991_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_153_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13505__A1 _13498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18941_ _19709_/C _18941_/B _19709_/B vssd1 vssd1 vccd1 vccd1 _18942_/B sky130_fd_sc_hd__and3_1
XFILLER_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14064_ _14056_/C _14064_/B _14064_/C vssd1 vssd1 vccd1 vccd1 _14285_/C sky130_fd_sc_hd__nand3b_2
XFILLER_193_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12314__B _16529_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ _12748_/X _20479_/A _13014_/Y vssd1 vssd1 vccd1 vccd1 _20620_/B sky130_fd_sc_hd__o21ai_1
X_18872_ _18872_/A _18872_/B vssd1 vssd1 vccd1 vccd1 _18872_/Y sky130_fd_sc_hd__nand2_2
XFILLER_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17823_ _17535_/A _17536_/A _17949_/A _17949_/B vssd1 vssd1 vccd1 vccd1 _17823_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_181_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17754_ _17644_/A _17613_/A _17605_/Y vssd1 vssd1 vccd1 vccd1 _17754_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__11819__A1 _12297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14966_ _14966_/A _14966_/B vssd1 vssd1 vccd1 vccd1 _15036_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16705_ _16707_/A _16707_/B _16706_/A _16706_/B vssd1 vssd1 vccd1 vccd1 _16709_/B
+ sky130_fd_sc_hd__nand4_1
X_13917_ _23355_/Q vssd1 vssd1 vccd1 vccd1 _14027_/A sky130_fd_sc_hd__inv_2
X_17685_ _17535_/A _17536_/A _17538_/X _17934_/B vssd1 vssd1 vccd1 vccd1 _17945_/A
+ sky130_fd_sc_hd__o22ai_2
X_14897_ _14899_/A _14899_/B _14908_/C _14898_/A vssd1 vssd1 vccd1 vccd1 _14900_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19424_ _19424_/A vssd1 vssd1 vccd1 vccd1 _19616_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_62_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19113__A _19381_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16636_ _15861_/X _16370_/A _16153_/B _16617_/X _16614_/Y vssd1 vssd1 vccd1 vccd1
+ _16637_/C sky130_fd_sc_hd__o221ai_1
XFILLER_23_708 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13848_ _13848_/A _13848_/B vssd1 vssd1 vccd1 vccd1 _13848_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19355_ _19391_/A _19392_/A vssd1 vssd1 vccd1 vccd1 _19355_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12244__A1 _11815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12244__B2 _12243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16567_ _16567_/A _16567_/B _16567_/C vssd1 vssd1 vccd1 vccd1 _16759_/C sky130_fd_sc_hd__nand3_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13779_ _13772_/X _13776_/Y _13778_/Y vssd1 vssd1 vccd1 vccd1 _13842_/B sky130_fd_sc_hd__o21bai_4
XANTENNA__18952__A _19530_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21503__B2 _20786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18306_ _18267_/A _18251_/B _18305_/X vssd1 vssd1 vccd1 vccd1 _18306_/Y sky130_fd_sc_hd__a21oi_1
X_15518_ _15483_/X _15493_/A _15516_/A _15517_/Y vssd1 vssd1 vccd1 vccd1 _15518_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_188_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19286_ _19457_/A _23544_/Q _19457_/C vssd1 vssd1 vccd1 vccd1 _19286_/Y sky130_fd_sc_hd__nand3_1
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16498_ _17248_/C vssd1 vssd1 vccd1 vccd1 _16526_/C sky130_fd_sc_hd__buf_2
XFILLER_31_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22474__A _22474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ _18185_/A _18185_/B _18185_/C _18187_/B _18187_/A vssd1 vssd1 vccd1 vccd1
+ _18239_/A sky130_fd_sc_hd__o32a_1
X_15449_ _15420_/D _15420_/Y _15447_/Y _15448_/X vssd1 vssd1 vccd1 vccd1 _15451_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18168_ _20151_/C _17753_/B _17753_/A _18169_/A _18218_/A vssd1 vssd1 vccd1 vccd1
+ _18170_/A sky130_fd_sc_hd__a32o_1
XFILLER_175_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_684 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_790 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17119_ _17117_/Y _17118_/X _17125_/A _17298_/A vssd1 vssd1 vccd1 vccd1 _17120_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_116_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23008__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18099_ _18094_/X _18095_/X _18098_/X vssd1 vssd1 vccd1 vccd1 _18104_/B sky130_fd_sc_hd__o21ai_1
X_20130_ _20151_/A _20212_/A _18335_/B _20369_/A _20067_/B vssd1 vssd1 vccd1 vccd1
+ _20182_/A sky130_fd_sc_hd__a41oi_4
XFILLER_171_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20061_ _20061_/A vssd1 vssd1 vccd1 vccd1 _20151_/A sky130_fd_sc_hd__buf_2
XANTENNA__15816__A _19165_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12180__B1 _11935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17789__A3 _18211_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18199__B1 _23532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20963_ _21545_/A _12722_/X _20962_/Y vssd1 vssd1 vccd1 vccd1 _20963_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__21742__A1 _22014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17946__B1 _23527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22368__B _22564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22702_ _22701_/C _22800_/B _22701_/A _22701_/B vssd1 vssd1 vccd1 vccd1 _22702_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17410__A2 _16683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20894_ _20894_/A _20894_/B vssd1 vssd1 vccd1 vccd1 _21046_/B sky130_fd_sc_hd__nand2_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22633_ _22633_/A _22633_/B vssd1 vssd1 vccd1 vccd1 _22633_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22564_ _22564_/A _22564_/B _22564_/C vssd1 vssd1 vccd1 vccd1 _22564_/X sky130_fd_sc_hd__and3_1
XFILLER_179_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1024 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17174__A1 _16934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21515_ _21513_/Y _21633_/A _21386_/A _21456_/Y vssd1 vssd1 vccd1 vccd1 _21517_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_22_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16382__A _16382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22495_ _22496_/A _22496_/B _22545_/B _22544_/A vssd1 vssd1 vccd1 vccd1 _22501_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21446_ _21448_/B _21371_/B _21371_/C _21448_/A _21561_/B vssd1 vssd1 vccd1 vccd1
+ _21510_/B sky130_fd_sc_hd__a32o_1
XFILLER_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18674__A1 _15882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19871__B1 _19525_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18674__B2 _16604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21377_ _21377_/A _21377_/B _21377_/C vssd1 vssd1 vccd1 vccd1 _21378_/C sky130_fd_sc_hd__nand3_1
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23116_ _23116_/A vssd1 vssd1 vccd1 vccd1 _23382_/D sky130_fd_sc_hd__clkbuf_1
X_20328_ _20328_/A _20328_/B _20328_/C vssd1 vssd1 vccd1 vccd1 _20329_/A sky130_fd_sc_hd__or3_1
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15726__A _16593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23047_ _13977_/B input29/X _23051_/S vssd1 vssd1 vccd1 vccd1 _23048_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20259_ _20311_/B _20312_/A vssd1 vssd1 vccd1 vccd1 _20261_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18977__A2 _11865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12710__A2 _12648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_796 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _14821_/A _14821_/B _14821_/C vssd1 vssd1 vccd1 vccd1 _14822_/A sky130_fd_sc_hd__a21o_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12150__A _19193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18756__B _18756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A wb_dat_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14751_ _14752_/A _14751_/B _14752_/C vssd1 vssd1 vccd1 vccd1 _14887_/A sky130_fd_sc_hd__nand3_2
XFILLER_28_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ _12189_/A vssd1 vssd1 vccd1 vccd1 _16860_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _13485_/A _13485_/B _13701_/Y _13415_/X vssd1 vssd1 vccd1 vccd1 _13705_/C
+ sky130_fd_sc_hd__a211o_1
X_17470_ _17562_/A _17562_/B _17473_/C _17473_/D vssd1 vssd1 vccd1 vccd1 _17471_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__21182__B _21279_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _23339_/Q _14668_/X _14673_/X _23307_/Q _14678_/X vssd1 vssd1 vccd1 vccd1
+ _14682_/X sky130_fd_sc_hd__a221o_1
X_11894_ _19165_/C vssd1 vssd1 vccd1 vccd1 _17149_/A sky130_fd_sc_hd__buf_4
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16421_ _16421_/A vssd1 vssd1 vccd1 vccd1 _16421_/Y sky130_fd_sc_hd__inv_2
X_13633_ _13553_/A _13470_/A _13630_/Y _13632_/X vssd1 vssd1 vccd1 vccd1 _13633_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19868__A _19868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15963__A2 _15862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19140_ _19140_/A _19140_/B _19140_/C vssd1 vssd1 vccd1 vccd1 _19410_/C sky130_fd_sc_hd__nand3_2
XFILLER_13_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19154__A2 _16055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16352_ _16340_/B _16296_/Y _16338_/Y vssd1 vssd1 vccd1 vccd1 _16575_/B sky130_fd_sc_hd__o21ai_2
XFILLER_34_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13564_ _13650_/A _21778_/D _21778_/C _13709_/A _13563_/X vssd1 vssd1 vccd1 vccd1
+ _13720_/B sky130_fd_sc_hd__a41o_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22294__A _22476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15303_ _15303_/A _15363_/D _15350_/C _15303_/D vssd1 vssd1 vccd1 vccd1 _15303_/X
+ sky130_fd_sc_hd__and4_1
X_19071_ _19071_/A vssd1 vssd1 vccd1 vccd1 _19071_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17388__A _17388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12515_ _17594_/A vssd1 vssd1 vccd1 vccd1 _18756_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_121_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16283_ _16275_/X _16278_/Y _16983_/B vssd1 vssd1 vccd1 vccd1 _16283_/Y sky130_fd_sc_hd__o21ai_1
X_13495_ _13495_/A vssd1 vssd1 vccd1 vccd1 _13495_/X sky130_fd_sc_hd__buf_2
XFILLER_185_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18022_ _18022_/A _18022_/B _18022_/C _18022_/D vssd1 vssd1 vccd1 vccd1 _18028_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12446_ _12246_/Y _12247_/Y _19180_/D vssd1 vssd1 vccd1 vccd1 _12446_/Y sky130_fd_sc_hd__o21ai_1
X_15234_ _15001_/X _14978_/A _15233_/Y vssd1 vssd1 vccd1 vccd1 _15234_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_173_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22997__A0 _21902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ _11931_/A _11931_/B _11792_/A _11792_/B vssd1 vssd1 vccd1 vccd1 _12377_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ _15163_/Y _15164_/Y _15188_/A vssd1 vssd1 vccd1 vccd1 _15185_/A sky130_fd_sc_hd__o21ai_1
XFILLER_176_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12325__A _16921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14116_ _14116_/A vssd1 vssd1 vccd1 vccd1 _14116_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_output83_A _14591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19973_ _17966_/A _17966_/B _19668_/A vssd1 vssd1 vccd1 vccd1 _19973_/X sky130_fd_sc_hd__a21o_1
X_15096_ _15096_/A _15096_/B _15238_/C vssd1 vssd1 vccd1 vccd1 _15096_/Y sky130_fd_sc_hd__nand3_2
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18924_ _18925_/A _18925_/B _23542_/Q vssd1 vssd1 vccd1 vccd1 _18926_/A sky130_fd_sc_hd__a21oi_1
X_14047_ _14026_/X _14121_/A _14183_/A _14039_/Y _14858_/A vssd1 vssd1 vccd1 vccd1
+ _14056_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_141_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21357__B _21358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12701__A2 _13184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18855_ _18958_/B _18856_/A _18854_/X vssd1 vssd1 vccd1 vccd1 _18858_/B sky130_fd_sc_hd__a21o_1
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17806_ _17806_/A _17806_/B vssd1 vssd1 vccd1 vccd1 _17806_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15100__B1 _14632_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18786_ _18868_/A _18868_/B _18868_/C _18785_/Y vssd1 vssd1 vccd1 vccd1 _18786_/Y
+ sky130_fd_sc_hd__a31oi_4
X_15998_ _15998_/A _15998_/B vssd1 vssd1 vccd1 vccd1 _15999_/B sky130_fd_sc_hd__xor2_1
XFILLER_36_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15651__A1 _16921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17737_ _17737_/A vssd1 vssd1 vccd1 vccd1 _17840_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12465__A1 _11931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ _14855_/Y _14856_/X _14825_/B vssd1 vssd1 vccd1 vccd1 _14949_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12465__B2 _11961_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22921__A0 _20481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17668_ _17493_/A _17493_/C _17493_/B vssd1 vssd1 vccd1 vccd1 _17668_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_51_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19407_ _19140_/C _19140_/A _19140_/B _19146_/A vssd1 vssd1 vccd1 vccd1 _19420_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__16600__B1 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16619_ _16619_/A _16815_/D vssd1 vssd1 vccd1 vccd1 _17249_/A sky130_fd_sc_hd__nand2_4
XFILLER_196_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17599_ _17589_/Y _17597_/Y _17598_/Y vssd1 vssd1 vccd1 vccd1 _17770_/A sky130_fd_sc_hd__o21ai_2
X_19338_ _19966_/A _19201_/C _19951_/D _19196_/Y vssd1 vssd1 vccd1 vccd1 _19339_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11976__B1 _11912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19269_ _19297_/A _19297_/B _19266_/X _19265_/X vssd1 vssd1 vccd1 vccd1 _19298_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_21300_ _21438_/A _21430_/C _21435_/C _21455_/A vssd1 vssd1 vccd1 vccd1 _21300_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_117_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22280_ _22562_/A _22280_/B _22562_/C vssd1 vssd1 vccd1 vccd1 _22283_/A sky130_fd_sc_hd__nand3_1
XANTENNA__22988__A0 _13802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21231_ _21236_/A _21236_/C vssd1 vssd1 vccd1 vccd1 _21231_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18656__A1 _12004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12235__A _16066_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16930__A _16935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21162_ _21082_/B _21083_/B _21161_/Y vssd1 vssd1 vccd1 vccd1 _21162_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16131__A2 _16153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20113_ _20113_/A _20113_/B _20185_/B vssd1 vssd1 vccd1 vccd1 _20116_/A sky130_fd_sc_hd__nand3_1
XFILLER_120_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21093_ _21088_/Y _21091_/Y _21092_/Y vssd1 vssd1 vccd1 vccd1 _21159_/A sky130_fd_sc_hd__o21bai_4
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20044_ _19973_/X _19980_/C _20058_/A vssd1 vssd1 vccd1 vccd1 _20054_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__22755__A3 _22392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A wb_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17761__A _17761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _21943_/X _21944_/X _21936_/Y vssd1 vssd1 vccd1 vccd1 _21995_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__22912__A0 _12712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16377__A _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ _20943_/A _20943_/B _20940_/X _20941_/Y _21057_/B vssd1 vssd1 vccd1 vccd1
+ _20950_/A sky130_fd_sc_hd__o221ai_1
XFILLER_121_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1018 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_808 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20877_ _20877_/A _21017_/B _21017_/C _21018_/A vssd1 vssd1 vccd1 vccd1 _20878_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22616_ _22629_/A _22629_/B vssd1 vssd1 vccd1 vccd1 _22616_/Y sky130_fd_sc_hd__nand2_1
X_23596_ _23598_/CLK _23596_/D vssd1 vssd1 vccd1 vccd1 _23596_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17147__A1 _16908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22547_ _22677_/A _22548_/C _22090_/A _22126_/X vssd1 vssd1 vccd1 vccd1 _22549_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_167_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12300_ _12300_/A _12300_/B _12300_/C vssd1 vssd1 vccd1 vccd1 _12547_/A sky130_fd_sc_hd__nand3_2
XFILLER_10_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ _13766_/A vssd1 vssd1 vccd1 vccd1 _13634_/A sky130_fd_sc_hd__clkbuf_1
X_22478_ _13547_/X _22461_/A _22362_/B _22476_/X _22477_/Y vssd1 vssd1 vccd1 vccd1
+ _22478_/X sky130_fd_sc_hd__o311a_1
XFILLER_120_1130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22979__A0 _13264_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ _12231_/A _12231_/B vssd1 vssd1 vccd1 vccd1 _12231_/Y sky130_fd_sc_hd__nor2_1
X_21429_ _21428_/X _21386_/A _21386_/B _21386_/C _21389_/A vssd1 vssd1 vccd1 vccd1
+ _21468_/A sky130_fd_sc_hd__a41oi_4
XFILLER_120_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16840__A _16840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12162_ _12143_/Y _12152_/X _12139_/Y vssd1 vssd1 vccd1 vccd1 _12162_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16970_ _16964_/A _16964_/B _16964_/C vssd1 vssd1 vccd1 vccd1 _16970_/Y sky130_fd_sc_hd__a21oi_1
X_12093_ _12093_/A vssd1 vssd1 vccd1 vccd1 _12093_/X sky130_fd_sc_hd__buf_2
XANTENNA__21177__B _21177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20081__B _20081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14684__A2 _14672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15921_ _15921_/A _15921_/B _15921_/C vssd1 vssd1 vccd1 vccd1 _15922_/A sky130_fd_sc_hd__nand3_1
XANTENNA__15175__B _15233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18640_ _18804_/B _18630_/X _18830_/B _18639_/Y vssd1 vssd1 vccd1 vccd1 _18669_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__23535__CLK _23558_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _15852_/A vssd1 vssd1 vccd1 vccd1 _15852_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16830__B1 _15972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21193__A _21493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14803_ _14934_/B _14934_/C vssd1 vssd1 vccd1 vccd1 _14803_/Y sky130_fd_sc_hd__nand2_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _18571_/A _18571_/B vssd1 vssd1 vccd1 vccd1 _18571_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12447__A1 _18511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _15783_/A vssd1 vssd1 vccd1 vccd1 _15785_/A sky130_fd_sc_hd__buf_2
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16287__A _17108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ _13133_/C _20886_/A _20584_/A _20585_/B vssd1 vssd1 vccd1 vccd1 _13085_/B
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__22903__A0 _12667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _17832_/A _17522_/B _17522_/C _17522_/D vssd1 vssd1 vccd1 vccd1 _17523_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13704__A _22388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12998__A2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14734_ _23256_/A vssd1 vssd1 vccd1 vccd1 _14734_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_189_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _16800_/A vssd1 vssd1 vccd1 vccd1 _11947_/C sky130_fd_sc_hd__inv_2
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17453_ _17453_/A _17453_/B _17453_/C vssd1 vssd1 vccd1 vccd1 _17469_/A sky130_fd_sc_hd__nand3_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _23367_/Q _14635_/X _14664_/X vssd1 vssd1 vccd1 vccd1 _14665_/X sky130_fd_sc_hd__o21a_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _16464_/A _11760_/A _11760_/B _12373_/A _19040_/A vssd1 vssd1 vccd1 vccd1
+ _11877_/X sky130_fd_sc_hd__o32a_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16404_ _16404_/A _16404_/B vssd1 vssd1 vccd1 vccd1 _16405_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13947__A1 _13977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13616_ _13616_/A _13616_/B vssd1 vssd1 vccd1 vccd1 _13616_/Y sky130_fd_sc_hd__nand2_1
X_17384_ _17384_/A _17384_/B vssd1 vssd1 vccd1 vccd1 _23585_/D sky130_fd_sc_hd__nor2_2
X_14596_ _13802_/B _14532_/X _14534_/X _14595_/X vssd1 vssd1 vccd1 vccd1 _14596_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19123_ _19703_/B _19123_/B _19123_/C _19548_/A vssd1 vssd1 vccd1 vccd1 _19123_/Y
+ sky130_fd_sc_hd__nand4_2
X_16335_ _16335_/A _16335_/B vssd1 vssd1 vccd1 vccd1 _16418_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13547_ _13547_/A vssd1 vssd1 vccd1 vccd1 _13547_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12981__C _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19054_ _19046_/Y _19048_/Y _19037_/A _19036_/B _19036_/A vssd1 vssd1 vccd1 vccd1
+ _19055_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16266_ _16266_/A _16266_/B _16266_/C vssd1 vssd1 vccd1 vccd1 _16281_/C sky130_fd_sc_hd__nand3_2
XFILLER_127_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13478_ _13538_/A _13538_/B _13598_/A _13477_/X vssd1 vssd1 vccd1 vccd1 _13540_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_195_1028 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18005_ _17610_/X _16742_/A _17860_/Y _17859_/Y vssd1 vssd1 vccd1 vccd1 _18005_/X
+ sky130_fd_sc_hd__o22a_1
X_15217_ _15286_/A _15286_/C vssd1 vssd1 vccd1 vccd1 _15218_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17846__A _17975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12429_ _11982_/Y _12428_/Y _12125_/Y vssd1 vssd1 vccd1 vccd1 _12429_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_173_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16197_ _15604_/X _16658_/C _16191_/A _16657_/B vssd1 vssd1 vccd1 vccd1 _17148_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__18638__B2 _18484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18102__A3 _17766_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15148_ _15148_/A _15220_/C vssd1 vssd1 vccd1 vccd1 _23274_/D sky130_fd_sc_hd__xor2_1
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15366__A _15366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11894__A _19165_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19956_ _20043_/A _20043_/B _19955_/X vssd1 vssd1 vccd1 vccd1 _19960_/A sky130_fd_sc_hd__a21boi_1
XFILLER_142_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15079_ _15077_/X _15076_/Y _15054_/A _14068_/X _14069_/X vssd1 vssd1 vccd1 vccd1
+ _15079_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_68_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18907_ _18907_/A vssd1 vssd1 vccd1 vccd1 _19091_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12686__A1 _12674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19887_ _19723_/C _19831_/X _19723_/B _19827_/A _19876_/B vssd1 vssd1 vccd1 vccd1
+ _19888_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_95_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_744 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17581__A _17581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18838_ _12105_/Y _19656_/A _19029_/A _19543_/A _19180_/D vssd1 vssd1 vccd1 vccd1
+ _18841_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_28_619 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14427__A2 _14876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18769_ _11815_/X _17846_/X _18617_/X _18768_/X vssd1 vssd1 vccd1 vccd1 _18966_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20800_ _21047_/A _20800_/B vssd1 vssd1 vccd1 vccd1 _21036_/B sky130_fd_sc_hd__nand2_1
X_21780_ _13805_/Y _21778_/Y _21779_/X _13810_/Y vssd1 vssd1 vccd1 vccd1 _21780_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_36_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21364__A_N _21285_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20731_ _20699_/A _20699_/B _20699_/C _20718_/B vssd1 vssd1 vccd1 vccd1 _20731_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19118__A2 _12247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23450_ _23462_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 _23450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20662_ _20662_/A _20662_/B vssd1 vssd1 vccd1 vccd1 _21277_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13052__C _13052_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19669__A3 _18461_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22401_ _22398_/Y _22401_/B _22401_/C vssd1 vssd1 vccd1 vccd1 _22402_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__22365__C _22365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23381_ _23381_/CLK _23381_/D vssd1 vssd1 vccd1 vccd1 _23381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20593_ _21008_/C _21008_/A _20593_/C vssd1 vssd1 vccd1 vccd1 _20597_/B sky130_fd_sc_hd__nand3b_1
XFILLER_177_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17459__C _17605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22332_ _22332_/A _22332_/B _22332_/C vssd1 vssd1 vccd1 vccd1 _22333_/C sky130_fd_sc_hd__nand3_1
XANTENNA__11788__B _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22263_ _22434_/A _22263_/B _22510_/B vssd1 vssd1 vccd1 vccd1 _22263_/X sky130_fd_sc_hd__and3_1
XFILLER_145_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14902__A3 _14061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21214_ _21218_/C _21217_/A _21218_/B vssd1 vssd1 vccd1 vccd1 _21215_/C sky130_fd_sc_hd__a21o_1
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21278__A _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22194_ _22184_/Y _22193_/Y _22290_/A _22158_/A vssd1 vssd1 vccd1 vccd1 _22214_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_183_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21145_ _21345_/A _21141_/X _23564_/Q _21142_/Y vssd1 vssd1 vccd1 vccd1 _21146_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__15312__B1 _15366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23558__CLK _23558_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19054__A1 _19046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21076_ _20906_/X _20907_/X _21079_/A _20908_/X vssd1 vssd1 vccd1 vccd1 _21194_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20027_ _19785_/X _20205_/A _20032_/A _20032_/B _20196_/C vssd1 vssd1 vccd1 vccd1
+ _20042_/B sky130_fd_sc_hd__o221ai_4
XFILLER_74_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19357__A2 _17741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13524__A _13732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _12071_/A _12105_/C _11798_/A vssd1 vssd1 vccd1 vccd1 _11896_/B sky130_fd_sc_hd__a21boi_4
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15442__C _15442_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _13011_/D vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ _13875_/B _21864_/Y _21861_/Y vssd1 vssd1 vccd1 vccd1 _21979_/B sky130_fd_sc_hd__a21bo_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11739_/B vssd1 vssd1 vccd1 vccd1 _11741_/A sky130_fd_sc_hd__clkinv_4
XFILLER_187_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ _20934_/A _20929_/B vssd1 vssd1 vccd1 vccd1 _20929_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16040__A1 _15920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16040__B2 _12020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14450_ _15116_/B vssd1 vssd1 vccd1 vccd1 _14975_/C sky130_fd_sc_hd__buf_2
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11684_/A _18653_/C _11665_/A vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20357__A _23554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14051__B1 _14031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13401_ _13486_/A _22420_/B _22420_/C _13400_/Y vssd1 vssd1 vccd1 vccd1 _13443_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_128_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11593_ _12510_/A _16807_/A _11593_/C vssd1 vssd1 vccd1 vccd1 _11972_/A sky130_fd_sc_hd__nand3_1
X_14381_ _14381_/A _14381_/B vssd1 vssd1 vccd1 vccd1 _14381_/Y sky130_fd_sc_hd__nor2_1
XFILLER_195_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23579_ _23584_/CLK _23579_/D vssd1 vssd1 vccd1 vccd1 _23579_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16120_ _15971_/X _15964_/Y _15998_/A vssd1 vssd1 vccd1 vccd1 _16120_/Y sky130_fd_sc_hd__a21oi_2
X_13332_ _13701_/A vssd1 vssd1 vccd1 vccd1 _21987_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16051_ _16377_/A _15800_/Y _17226_/D _16372_/A _16046_/Y vssd1 vssd1 vccd1 vccd1
+ _16094_/B sky130_fd_sc_hd__o2111a_1
XFILLER_6_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13263_ _23322_/Q vssd1 vssd1 vccd1 vccd1 _13264_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15002_ _15459_/B _15001_/X _15459_/A _14991_/A vssd1 vssd1 vccd1 vccd1 _15002_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12214_ _12324_/A vssd1 vssd1 vccd1 vccd1 _12214_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13194_ _13171_/B _13171_/A _13149_/Y _13148_/X vssd1 vssd1 vccd1 vccd1 _13194_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_194_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14106__A1 _14029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19810_ _19819_/B _19819_/A _19820_/A vssd1 vssd1 vccd1 vccd1 _19810_/Y sky130_fd_sc_hd__a21boi_1
X_12145_ _12145_/A _12145_/B vssd1 vssd1 vccd1 vccd1 _12324_/A sky130_fd_sc_hd__nand2_4
XFILLER_123_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15854__B2 _15975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19741_ _19740_/A _19740_/B _19730_/A _19730_/B vssd1 vssd1 vccd1 vccd1 _19742_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_12076_ _19703_/C vssd1 vssd1 vccd1 vccd1 _19811_/A sky130_fd_sc_hd__clkbuf_4
X_16953_ _16953_/A _16953_/B _16953_/C vssd1 vssd1 vccd1 vccd1 _17173_/B sky130_fd_sc_hd__nand3_1
X_15904_ _15904_/A vssd1 vssd1 vccd1 vccd1 _16054_/A sky130_fd_sc_hd__buf_2
X_19672_ _19682_/A _19682_/B _19672_/C vssd1 vssd1 vccd1 vccd1 _19672_/Y sky130_fd_sc_hd__nand3_1
XFILLER_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16884_ _16879_/X _16882_/Y _16894_/D vssd1 vssd1 vccd1 vccd1 _16884_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__21635__B _21635_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18623_ _18778_/C _18778_/A _18778_/B _18931_/A _18615_/Y vssd1 vssd1 vccd1 vccd1
+ _18623_/X sky130_fd_sc_hd__a32o_1
XFILLER_2_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _15830_/X _16027_/D _17057_/A _16028_/A _16029_/B vssd1 vssd1 vccd1 vccd1
+ _15836_/C sky130_fd_sc_hd__a32oi_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18554_ _18554_/A _18554_/B _18554_/C vssd1 vssd1 vccd1 vccd1 _18555_/C sky130_fd_sc_hd__nand3_1
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15766_ _15766_/A vssd1 vssd1 vccd1 vccd1 _15766_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12978_ _13106_/B vssd1 vssd1 vccd1 vccd1 _12978_/Y sky130_fd_sc_hd__inv_2
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17505_ _17513_/A _17513_/B _17513_/C vssd1 vssd1 vccd1 vccd1 _17677_/C sky130_fd_sc_hd__and3_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14717_ _23412_/Q _14640_/A _14534_/X _23444_/Q _14716_/X vssd1 vssd1 vccd1 vccd1
+ _14717_/X sky130_fd_sc_hd__a221o_4
XANTENNA__16167__D _20062_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18485_ _18476_/X _18484_/X _12149_/X _15704_/A _19846_/A vssd1 vssd1 vccd1 vccd1
+ _18486_/A sky130_fd_sc_hd__o2111ai_4
X_11929_ _11618_/C _11606_/X _18999_/C _11672_/Y vssd1 vssd1 vccd1 vccd1 _11931_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_75_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15697_ _15630_/Y _15713_/B _14569_/X vssd1 vssd1 vccd1 vccd1 _15698_/B sky130_fd_sc_hd__a21oi_4
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16031__A1 _16464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22466__B _22566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17436_ _17434_/X _17435_/X _15682_/D _15974_/C _18947_/A vssd1 vssd1 vccd1 vccd1
+ _17571_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_127_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14648_ _23429_/Q vssd1 vssd1 vccd1 vccd1 _15735_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18308__B1 _18154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19181__A1_N _19168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14593__A1 _23579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _17196_/Y _17200_/Y _17369_/C _17024_/A vssd1 vssd1 vccd1 vccd1 _17522_/C
+ sky130_fd_sc_hd__a22o_2
X_14579_ _15674_/C _14575_/X _14576_/X _14578_/X vssd1 vssd1 vccd1 vccd1 _14579_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14593__B2 _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19106_ _19106_/A _19106_/B vssd1 vssd1 vccd1 vccd1 _19294_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16318_ _16318_/A _17845_/C _16318_/C vssd1 vssd1 vccd1 vccd1 _16321_/A sky130_fd_sc_hd__nand3_1
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17298_ _17298_/A _17298_/B vssd1 vssd1 vccd1 vccd1 _17299_/C sky130_fd_sc_hd__nand2_1
XANTENNA__17531__A1 _17943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16334__A2 _16408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20130__A3 _18335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_192 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19037_ _19037_/A _19052_/B vssd1 vssd1 vccd1 vccd1 _19037_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17576__A _19694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16249_ _16268_/B _16249_/B vssd1 vssd1 vccd1 vccd1 _16249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13002__D1 _20781_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16480__A _16480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18087__A2 _17960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_13_0_bq_clk_i clkbuf_3_6_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _23575_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_126_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12108__B1 _12104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13305__C1 _13304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19939_ _19939_/A vssd1 vssd1 vccd1 vccd1 _19939_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22950_ _22950_/A vssd1 vssd1 vccd1 vccd1 _23309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23463__D _23475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21901_ _13602_/C _21901_/B _22141_/B _21901_/D vssd1 vssd1 vccd1 vccd1 _22028_/A
+ sky130_fd_sc_hd__nand4b_4
XFILLER_56_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22881_ _23285_/Q _22881_/B _22887_/B vssd1 vssd1 vccd1 vccd1 _22881_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21832_ _21832_/A _22667_/D vssd1 vssd1 vccd1 vccd1 _21832_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14281__B1 _14245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23252__S _23254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18011__A2 _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21763_ _13825_/Y _21922_/A _21762_/Y _13410_/A vssd1 vssd1 vccd1 vccd1 _21783_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_93_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20714_ _20714_/A _20714_/B vssd1 vssd1 vccd1 vccd1 _20716_/B sky130_fd_sc_hd__nand2_1
X_23502_ _23510_/CLK _23502_/D vssd1 vssd1 vccd1 vccd1 _23502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21694_ _21694_/A _21704_/C _21694_/C vssd1 vssd1 vccd1 vccd1 _21698_/C sky130_fd_sc_hd__nand3_1
XFILLER_12_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19388__D _19569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19966__A _19966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14584__A1 _13379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23433_ _23433_/CLK _23433_/D vssd1 vssd1 vccd1 vccd1 _23433_/Q sky130_fd_sc_hd__dfxtp_1
X_20645_ _20921_/A _20921_/B _20645_/C vssd1 vssd1 vccd1 vccd1 _20645_/Y sky130_fd_sc_hd__nand3_2
XFILLER_177_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23364_ _23402_/CLK _23364_/D vssd1 vssd1 vccd1 vccd1 _23364_/Q sky130_fd_sc_hd__dfxtp_4
X_20576_ _20595_/C _20595_/B _13075_/Y _13072_/Y vssd1 vssd1 vccd1 vccd1 _20576_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__22392__A _22392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20905__A _21072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22315_ _22291_/Y _22313_/X _22323_/C vssd1 vssd1 vccd1 vccd1 _22315_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_106_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23295_ _23295_/CLK _23295_/D vssd1 vssd1 vccd1 vccd1 _23295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_760 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22246_ _22246_/A _22246_/B vssd1 vssd1 vccd1 vccd1 _22246_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17286__B1 _17260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22177_ _22290_/B _22166_/Y _22290_/A vssd1 vssd1 vccd1 vccd1 _22177_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__20062__D _20133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19027__A1 _19548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21128_ _21132_/A vssd1 vssd1 vccd1 vccd1 _21128_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17038__B1 _15968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1040 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21455__B _21455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13950_ _13948_/X _14029_/A _14188_/C vssd1 vssd1 vccd1 vccd1 _13951_/B sky130_fd_sc_hd__o21ai_1
X_21059_ _21084_/A _21212_/A _21202_/B _21056_/B vssd1 vssd1 vccd1 vccd1 _21097_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__17589__A1 _17974_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21385__A2 _21490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22582__A1 _21997_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_86 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16549__B _16549_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ _12901_/A _12901_/B _12901_/C _12901_/D vssd1 vssd1 vccd1 vccd1 _12902_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_100_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13881_ _14459_/D vssd1 vssd1 vccd1 vccd1 _14377_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21174__C _21174_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15620_ _23422_/Q _15665_/B vssd1 vssd1 vccd1 vccd1 _15634_/C sky130_fd_sc_hd__nand2_4
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _20532_/B vssd1 vssd1 vccd1 vccd1 _13115_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15528_/C _15528_/B _15339_/A vssd1 vssd1 vccd1 vccd1 _15552_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12763_/A vssd1 vssd1 vccd1 vccd1 _12792_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14502_/A vssd1 vssd1 vccd1 vccd1 _23270_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _18226_/A _18223_/X _18225_/B vssd1 vssd1 vccd1 vccd1 _18285_/A sky130_fd_sc_hd__o21a_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _16677_/A vssd1 vssd1 vccd1 vccd1 _16027_/B sky130_fd_sc_hd__clkbuf_2
X_15482_ _15420_/D _15420_/Y _15447_/Y _15448_/X vssd1 vssd1 vccd1 vccd1 _15483_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_43_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12694_/A vssd1 vssd1 vccd1 vccd1 _12695_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17221_ _17221_/A _17221_/B _17221_/C vssd1 vssd1 vccd1 vccd1 _17221_/X sky130_fd_sc_hd__and3_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14433_ _14806_/A _14448_/A _14867_/C _14433_/D vssd1 vssd1 vccd1 vccd1 _14465_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__22098__B1 _22099_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11645_ _15956_/A vssd1 vssd1 vccd1 vccd1 _16802_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15772__B1 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17152_ _17152_/A _17152_/B vssd1 vssd1 vccd1 vccd1 _17161_/A sky130_fd_sc_hd__nand2_1
Xinput15 wb_dat_i[17] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
X_14364_ _14414_/A _14416_/B _14414_/B vssd1 vssd1 vccd1 vccd1 _14365_/C sky130_fd_sc_hd__a21boi_1
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11576_ _23590_/Q vssd1 vssd1 vccd1 vccd1 _16815_/B sky130_fd_sc_hd__clkbuf_2
Xinput26 wb_dat_i[27] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_2
XANTENNA__16316__A2 _16451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 wb_dat_i[8] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_4
X_16103_ _16425_/B _16425_/C _16425_/A vssd1 vssd1 vccd1 vccd1 _16104_/A sky130_fd_sc_hd__a21oi_1
Xinput48 x[5] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_4
X_13315_ _21925_/B vssd1 vssd1 vccd1 vccd1 _21764_/C sky130_fd_sc_hd__clkbuf_2
X_17083_ _12518_/X _16311_/X _17069_/A _17070_/A _17077_/B vssd1 vssd1 vccd1 vccd1
+ _17083_/X sky130_fd_sc_hd__o311a_1
XFILLER_122_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16867__A3 _17605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14295_ _14256_/A _14324_/B _14255_/A vssd1 vssd1 vccd1 vccd1 _14298_/A sky130_fd_sc_hd__o21ai_1
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12036__C _16796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16034_ _12036_/A _12036_/B _18434_/B _15749_/B _15749_/A vssd1 vssd1 vccd1 vccd1
+ _16308_/D sky130_fd_sc_hd__a32oi_4
XANTENNA__19266__A1 _12353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13246_ _13769_/A vssd1 vssd1 vccd1 vccd1 _22365_/C sky130_fd_sc_hd__buf_2
XANTENNA__19266__B2 _19082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17546__D _19862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21073__B2 _12979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13177_ _13177_/A _13177_/B _13177_/C vssd1 vssd1 vccd1 vccd1 _13177_/X sky130_fd_sc_hd__and3_1
XFILLER_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12128_ _12010_/B _12125_/Y _12051_/A _18645_/A _12119_/Y vssd1 vssd1 vccd1 vccd1
+ _12399_/C sky130_fd_sc_hd__o221ai_4
X_17985_ _20133_/D vssd1 vssd1 vccd1 vccd1 _18100_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19724_ _19483_/Y _19692_/Y _19521_/B _19521_/C vssd1 vssd1 vccd1 vccd1 _19725_/C
+ sky130_fd_sc_hd__a22oi_4
XANTENNA__19116__A _19116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ _12059_/A _12200_/B _12205_/A _12059_/D vssd1 vssd1 vccd1 vccd1 _12064_/B
+ sky130_fd_sc_hd__nand4_2
X_16936_ _17166_/A _16936_/B _16936_/C vssd1 vssd1 vccd1 vccd1 _16936_/Y sky130_fd_sc_hd__nand3_2
XFILLER_81_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_736 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19655_ _16437_/X _20080_/A _19649_/A vssd1 vssd1 vccd1 vccd1 _19655_/X sky130_fd_sc_hd__o21a_1
X_16867_ _18859_/D _17605_/A _17605_/B _17107_/A _16860_/Y vssd1 vssd1 vccd1 vccd1
+ _16870_/A sky130_fd_sc_hd__a32o_1
XFILLER_65_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18606_ _11815_/X _18604_/X _18605_/Y vssd1 vssd1 vccd1 vccd1 _18606_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15818_ _15813_/A _15813_/B _15817_/Y vssd1 vssd1 vccd1 vccd1 _16020_/A sky130_fd_sc_hd__o21ai_2
X_19586_ _19376_/A _19572_/X _19573_/C vssd1 vssd1 vccd1 vccd1 _19587_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__13066__A1 _13131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15082__C _15356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16798_ _17043_/A _16798_/B _18947_/C vssd1 vssd1 vccd1 vccd1 _16812_/B sky130_fd_sc_hd__nand3_2
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14802__A2 _14911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18537_ _12378_/A _12378_/B _17593_/A _17591_/A _19364_/C vssd1 vssd1 vccd1 vccd1
+ _18537_/Y sky130_fd_sc_hd__o221ai_4
X_15749_ _15749_/A _15749_/B vssd1 vssd1 vccd1 vccd1 _15968_/A sky130_fd_sc_hd__nand2_4
XFILLER_34_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18468_ _18468_/A _23391_/Q _18810_/A vssd1 vssd1 vccd1 vccd1 _18469_/C sky130_fd_sc_hd__nor3_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17419_ _17265_/Y _17414_/X _17260_/Y vssd1 vssd1 vccd1 vccd1 _17426_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__14566__A1 _13253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18399_ _18400_/A _18414_/C _18400_/C vssd1 vssd1 vccd1 vccd1 _18399_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12508__A _12508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20430_ _20430_/A _20430_/B vssd1 vssd1 vccd1 vccd1 _20431_/C sky130_fd_sc_hd__xor2_4
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20361_ _20120_/X _20205_/X _20344_/X _20343_/Y _20339_/A vssd1 vssd1 vccd1 vccd1
+ _20361_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_146_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15819__A _17066_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14723__A _23594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12329__B1 _19512_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22100_ _21964_/A _21964_/C _21964_/B vssd1 vssd1 vccd1 vccd1 _22102_/C sky130_fd_sc_hd__a21boi_4
XFILLER_173_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23080_ _23367_/Q input15/X _23084_/S vssd1 vssd1 vccd1 vccd1 _23081_/A sky130_fd_sc_hd__mux2_1
X_20292_ _20295_/A _20295_/B vssd1 vssd1 vccd1 vccd1 _20337_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22031_ _22031_/A vssd1 vssd1 vccd1 vccd1 _22562_/C sky130_fd_sc_hd__buf_2
XANTENNA__21064__A1 _21545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18849__B _19364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17753__B _17753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22933_ _22933_/A vssd1 vssd1 vccd1 vccd1 _23301_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__21772__C1 _22264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22864_ _22836_/A _22839_/A _22862_/Y vssd1 vssd1 vccd1 vccd1 _22865_/B sky130_fd_sc_hd__o21a_1
XFILLER_73_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17991__A1 _12088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21815_ _22236_/A _21815_/B _21815_/C vssd1 vssd1 vccd1 vccd1 _21820_/A sky130_fd_sc_hd__nor3_2
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16385__A _17845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22795_ _22700_/C _22637_/A _22637_/B _22830_/A _22830_/C vssd1 vssd1 vccd1 vccd1
+ _22797_/B sky130_fd_sc_hd__a311o_1
XANTENNA__18535__A3 _17587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20619__B _21054_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21746_ _22057_/A _22020_/B _22024_/C _22033_/A vssd1 vssd1 vccd1 vccd1 _21906_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_52_783 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17743__A1 _17741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12280__A2 _11611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19696__A _19698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14557__A1 _13977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14557__B2 _12667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21677_ _21704_/C vssd1 vssd1 vccd1 vccd1 _21698_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23416_ _23416_/CLK _23416_/D vssd1 vssd1 vccd1 vccd1 _23416_/Q sky130_fd_sc_hd__dfxtp_2
X_20628_ _20628_/A _20628_/B _20628_/C vssd1 vssd1 vccd1 vccd1 _20783_/A sky130_fd_sc_hd__nand3_2
XFILLER_125_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11776__D1 _11749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22553__C _22553_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20559_ _20578_/A _20578_/B _20578_/C vssd1 vssd1 vccd1 vccd1 _20570_/A sky130_fd_sc_hd__nand3_1
X_23347_ _23347_/CLK _23347_/D vssd1 vssd1 vccd1 vccd1 _23347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13100_ _13205_/C _13205_/A _13205_/B vssd1 vssd1 vccd1 vccd1 _13100_/X sky130_fd_sc_hd__and3_1
XFILLER_192_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14080_ _14752_/A vssd1 vssd1 vccd1 vccd1 _14178_/B sky130_fd_sc_hd__buf_2
X_23278_ _23510_/CLK _23278_/D vssd1 vssd1 vccd1 vccd1 _23278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13031_ _21061_/A _12632_/A _13001_/A _13005_/Y vssd1 vssd1 vccd1 vccd1 _13031_/Y
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__21055__B2 _20471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22229_ _22086_/Y _22119_/X _22093_/D vssd1 vssd1 vccd1 vccd1 _22234_/A sky130_fd_sc_hd__o21ai_1
XFILLER_161_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15809__B2 _15800_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A x[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21170__A1_N _21276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16482__A1 _16478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17770_ _17770_/A _17770_/B vssd1 vssd1 vccd1 vccd1 _17770_/Y sky130_fd_sc_hd__nand2_1
X_14982_ _14976_/Y _14979_/X _14981_/X vssd1 vssd1 vccd1 vccd1 _15124_/A sky130_fd_sc_hd__o21ai_1
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22555__B2 _13465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23276__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16721_ _16715_/Y _16718_/Y _16720_/Y vssd1 vssd1 vccd1 vccd1 _16721_/Y sky130_fd_sc_hd__a21oi_2
X_13933_ _13933_/A _13933_/B vssd1 vssd1 vccd1 vccd1 _13933_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19440_ _19427_/X _19433_/Y _19439_/Y vssd1 vssd1 vccd1 vccd1 _19440_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19971__A2 _19670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16652_ _16139_/Y _16169_/Y _16645_/Y _16651_/Y vssd1 vssd1 vccd1 vccd1 _16722_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__21913__B _21913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13864_ _13864_/A vssd1 vssd1 vccd1 vccd1 _13864_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_823 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15603_ _15615_/A _15634_/A _15642_/A vssd1 vssd1 vccd1 vccd1 _16658_/B sky130_fd_sc_hd__nand3_2
X_19371_ _19371_/A _19371_/B vssd1 vssd1 vccd1 vccd1 _19374_/A sky130_fd_sc_hd__nand2_1
X_12815_ _13151_/A _12815_/B _12815_/C vssd1 vssd1 vccd1 vccd1 _12816_/A sky130_fd_sc_hd__or3_1
X_16583_ _16283_/Y _17026_/C _16774_/B vssd1 vssd1 vccd1 vccd1 _16584_/A sky130_fd_sc_hd__nand3b_1
X_13795_ _13615_/A _13791_/A _13793_/Y vssd1 vssd1 vccd1 vccd1 _13797_/A sky130_fd_sc_hd__o21ai_1
XFILLER_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18322_ _18322_/A _18349_/B vssd1 vssd1 vccd1 vccd1 _18388_/A sky130_fd_sc_hd__nand2_1
XFILLER_163_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15534_ _15225_/B _15446_/A _15488_/X vssd1 vssd1 vccd1 vccd1 _15538_/A sky130_fd_sc_hd__a21bo_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12746_ _20473_/A vssd1 vssd1 vccd1 vccd1 _20962_/A sky130_fd_sc_hd__buf_2
XANTENNA__16537__A2 _17445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _18253_/A _18253_/B vssd1 vssd1 vccd1 vccd1 _18254_/C sky130_fd_sc_hd__nor2_1
XFILLER_124_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14548__A1 _13945_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16445__D _17445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15465_ _15467_/B _15467_/C _15467_/A vssd1 vssd1 vccd1 vccd1 _15466_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__14548__B2 _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12328__A _19180_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12677_ _12677_/A vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_187_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17204_ _17035_/X _16923_/A _17200_/C _17200_/A _16917_/X vssd1 vssd1 vccd1 vccd1
+ _17204_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14416_ _14416_/A _14416_/B vssd1 vssd1 vccd1 vccd1 _14418_/B sky130_fd_sc_hd__nand2_1
X_18184_ _18110_/B _18110_/A _18108_/A vssd1 vssd1 vccd1 vccd1 _18185_/A sky130_fd_sc_hd__o21a_1
XANTENNA__19487__A1 _18656_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11628_ _12174_/A _12173_/A _12175_/A vssd1 vssd1 vccd1 vccd1 _12207_/A sky130_fd_sc_hd__o21ai_4
XFILLER_168_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15396_ _15391_/A _15391_/B _15435_/A _15435_/B vssd1 vssd1 vccd1 vccd1 _15396_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17135_ _17156_/B vssd1 vssd1 vccd1 vccd1 _17359_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14347_ _14361_/C _14361_/A _14347_/C vssd1 vssd1 vccd1 vccd1 _14347_/X sky130_fd_sc_hd__and3_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17066_ _19700_/C _19700_/D _17066_/C vssd1 vssd1 vccd1 vccd1 _17077_/B sky130_fd_sc_hd__and3_1
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14278_ _13914_/A _14263_/Y _14340_/B _14260_/Y vssd1 vssd1 vccd1 vccd1 _14279_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16017_ _16017_/A _16017_/B _16017_/C vssd1 vssd1 vccd1 vccd1 _16018_/A sky130_fd_sc_hd__nand3_1
X_13229_ _13226_/X _13224_/B _13394_/B _13228_/X vssd1 vssd1 vccd1 vccd1 _13659_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22794__A1 _22237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21376__A _21376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17968_ _18080_/A vssd1 vssd1 vccd1 vccd1 _20146_/A sky130_fd_sc_hd__buf_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19947__C1 _18434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19707_ _19831_/A _19831_/B _19831_/C vssd1 vssd1 vccd1 vccd1 _19723_/A sky130_fd_sc_hd__nand3_1
X_16919_ _15932_/A _16665_/A _17029_/A _16918_/Y vssd1 vssd1 vccd1 vccd1 _17133_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11837__A2 _16921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17899_ _17899_/A _17899_/B _18017_/D vssd1 vssd1 vccd1 vccd1 _17899_/X sky130_fd_sc_hd__and3_1
XFILLER_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19638_ _19638_/A _19638_/B _19638_/C vssd1 vssd1 vccd1 vccd1 _19638_/Y sky130_fd_sc_hd__nand3_1
XFILLER_93_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12247__C1 _12245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19569_ _19569_/A vssd1 vssd1 vccd1 vccd1 _19572_/A sky130_fd_sc_hd__inv_2
XFILLER_168_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15984__B1 _19017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21600_ _21602_/A _21602_/B _21599_/X vssd1 vssd1 vccd1 vccd1 _21645_/B sky130_fd_sc_hd__a21oi_1
XFILLER_178_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22580_ _22579_/Y _22573_/A _22574_/Y vssd1 vssd1 vccd1 vccd1 _22580_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_178_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21531_ _21529_/X _21576_/A _21614_/D vssd1 vssd1 vccd1 vccd1 _21541_/A sky130_fd_sc_hd__a21o_1
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12238__A _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21462_ _21463_/A _21463_/B _21461_/Y vssd1 vssd1 vccd1 vccd1 _21464_/A sky130_fd_sc_hd__a21bo_1
XFILLER_193_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20413_ _20452_/B _20415_/A _20415_/B _20362_/Y vssd1 vssd1 vccd1 vccd1 _20414_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_135_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23201_ _23201_/A vssd1 vssd1 vccd1 vccd1 _23420_/D sky130_fd_sc_hd__clkbuf_1
X_21393_ _21390_/X _21465_/B _21392_/X vssd1 vssd1 vccd1 vccd1 _21424_/A sky130_fd_sc_hd__a21oi_1
XFILLER_162_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20344_ _20295_/A _20295_/B _20336_/A _20336_/B vssd1 vssd1 vccd1 vccd1 _20344_/X
+ sky130_fd_sc_hd__a211o_1
X_23132_ _12121_/B input37/X _23134_/S vssd1 vssd1 vccd1 vccd1 _23133_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_964 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12317__A3 _16549_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23063_ _23063_/A vssd1 vssd1 vccd1 vccd1 _23359_/D sky130_fd_sc_hd__clkbuf_1
X_20275_ _20400_/B vssd1 vssd1 vccd1 vccd1 _20328_/A sky130_fd_sc_hd__inv_2
XFILLER_103_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_880 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22014_ _22014_/A _22364_/B _22380_/C _22381_/C vssd1 vssd1 vccd1 vccd1 _22136_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20902__B _20902_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19650__A1 _12323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22916_ _12756_/B input37/X _22918_/S vssd1 vssd1 vccd1 vccd1 _22917_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15731__B _15731_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22847_ _22847_/A vssd1 vssd1 vccd1 vccd1 _22847_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_1019 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12600_ _20782_/C vssd1 vssd1 vccd1 vccd1 _21036_/C sky130_fd_sc_hd__buf_2
XANTENNA__17004__A _23521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13580_ _13712_/D vssd1 vssd1 vccd1 vccd1 _13582_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_169_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22778_ _22630_/X _22813_/B _22858_/A vssd1 vssd1 vccd1 vccd1 _22780_/A sky130_fd_sc_hd__o21ai_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12531_/A _12531_/B _12531_/C vssd1 vssd1 vccd1 vccd1 _12531_/X sky130_fd_sc_hd__and3_1
X_21729_ _21722_/B _21728_/A _21728_/Y vssd1 vssd1 vccd1 vccd1 _21729_/X sky130_fd_sc_hd__o21a_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22564__B _22564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _15250_/A _15250_/B _15250_/C _15250_/D vssd1 vssd1 vccd1 vccd1 _15326_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_71_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12462_ _12474_/A vssd1 vssd1 vccd1 vccd1 _19017_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__12005__A2 _16619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ _14312_/D vssd1 vssd1 vccd1 vccd1 _15116_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_166_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18480__D _19180_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15181_ _15310_/B _14990_/A _14990_/B _15301_/A _15010_/A vssd1 vssd1 vccd1 vccd1
+ _15181_/X sky130_fd_sc_hd__a32o_1
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12393_ _12393_/A _12393_/B vssd1 vssd1 vccd1 vccd1 _12393_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _14172_/A _14172_/B _14276_/A vssd1 vssd1 vccd1 vccd1 _14133_/B sky130_fd_sc_hd__and3_1
XFILLER_180_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13505__A2 _13498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18940_ _18944_/C _19141_/A _19141_/B vssd1 vssd1 vccd1 vccd1 _19410_/A sky130_fd_sc_hd__nand3b_2
X_14063_ _14063_/A _14063_/B vssd1 vssd1 vccd1 vccd1 _14064_/C sky130_fd_sc_hd__nand2_1
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12713__B1 _12712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13014_ _13014_/A _20494_/D vssd1 vssd1 vccd1 vccd1 _13014_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18871_ _18808_/B _18808_/C _18808_/A vssd1 vssd1 vccd1 vccd1 _18871_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17822_ _17686_/X _17541_/Y _17680_/C _17832_/D vssd1 vssd1 vccd1 vccd1 _17949_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_842 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17753_ _17753_/A _17753_/B _20055_/C _20055_/D vssd1 vssd1 vccd1 vccd1 _17760_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_130_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14965_ _23270_/D _14965_/B _14849_/Y vssd1 vssd1 vccd1 vccd1 _15220_/A sky130_fd_sc_hd__or3b_1
XFILLER_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16207__A1 _15920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16704_ _16704_/A _16704_/B vssd1 vssd1 vccd1 vccd1 _16707_/B sky130_fd_sc_hd__nand2_1
XANTENNA__21200__B2 _12862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13916_ _13949_/A vssd1 vssd1 vccd1 vccd1 _14189_/A sky130_fd_sc_hd__clkbuf_2
X_17684_ _18207_/A _18208_/A _17538_/X _17527_/C _17935_/D vssd1 vssd1 vccd1 vccd1
+ _17684_/X sky130_fd_sc_hd__o221a_1
XANTENNA__15232__A1_N _15225_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14896_ _14896_/A _14896_/B _14896_/C vssd1 vssd1 vccd1 vccd1 _14898_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19533__A1_N _19534_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23561__D _23561_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21751__A2 _21906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19423_ _19423_/A _19423_/B _19423_/C vssd1 vssd1 vccd1 vccd1 _19424_/A sky130_fd_sc_hd__nand3_1
X_16635_ _16635_/A _16635_/B vssd1 vssd1 vccd1 vccd1 _16637_/B sky130_fd_sc_hd__nand2_1
XANTENNA__19113__B _19694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13847_ _13674_/A _13680_/D _13846_/Y vssd1 vssd1 vccd1 vccd1 _13848_/B sky130_fd_sc_hd__a21oi_2
XFILLER_16_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19354_ _19354_/A _19354_/B vssd1 vssd1 vccd1 vccd1 _19392_/A sky130_fd_sc_hd__nand2_1
X_16566_ _16566_/A _16566_/B _16566_/C vssd1 vssd1 vccd1 vccd1 _16567_/C sky130_fd_sc_hd__nand3_1
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12244__A2 _16523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13778_ _13776_/B _13777_/Y _13776_/A vssd1 vssd1 vccd1 vccd1 _13778_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18952__B _19703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18305_ _18305_/A _18305_/B vssd1 vssd1 vccd1 vccd1 _18305_/X sky130_fd_sc_hd__or2_1
XFILLER_149_917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15517_ _15517_/A _15540_/A vssd1 vssd1 vccd1 vccd1 _15517_/Y sky130_fd_sc_hd__nand2_1
X_19285_ _20031_/A _19294_/B _19278_/C _19281_/X vssd1 vssd1 vccd1 vccd1 _19457_/C
+ sky130_fd_sc_hd__o211ai_1
X_12729_ _12709_/A _12722_/X _12723_/X _12725_/X _12728_/Y vssd1 vssd1 vccd1 vccd1
+ _12734_/B sky130_fd_sc_hd__o221ai_2
X_16497_ _16497_/A vssd1 vssd1 vccd1 vccd1 _16526_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_175_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18236_ _18236_/A _18236_/B _18236_/C vssd1 vssd1 vccd1 vccd1 _18239_/C sky130_fd_sc_hd__nor3_1
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15448_ _15536_/A _14999_/Y _15446_/X _15445_/X vssd1 vssd1 vccd1 vccd1 _15448_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_176_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18167_ _18172_/C vssd1 vssd1 vccd1 vccd1 _18218_/A sky130_fd_sc_hd__clkbuf_2
X_15379_ _15379_/A _15379_/B _15377_/X vssd1 vssd1 vccd1 vccd1 _15382_/B sky130_fd_sc_hd__or3b_1
XFILLER_157_994 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_696 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17118_ _17118_/A _17118_/B _17301_/B vssd1 vssd1 vccd1 vccd1 _17118_/X sky130_fd_sc_hd__and3_1
X_18098_ _16478_/X _17465_/X _20210_/A _18328_/A _17992_/C vssd1 vssd1 vccd1 vccd1
+ _18098_/X sky130_fd_sc_hd__o41a_1
XFILLER_143_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17049_ _17050_/A _16819_/X _17249_/A _17250_/A vssd1 vssd1 vccd1 vccd1 _17975_/A
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_132_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20060_ _20060_/A _20060_/B _20060_/C vssd1 vssd1 vccd1 vccd1 _20071_/C sky130_fd_sc_hd__nand3_1
XFILLER_131_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15816__B _16314_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12180__A1 _11926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23591__CLK _23598_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18199__A1 _18154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15832__A _16634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20962_ _20962_/A _20962_/B _20962_/C vssd1 vssd1 vccd1 vccd1 _20962_/Y sky130_fd_sc_hd__nand3_2
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21742__A2 _13804_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22701_ _22701_/A _22701_/B _22701_/C _22800_/B vssd1 vssd1 vccd1 vccd1 _22707_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_198_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14448__A _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20893_ _23300_/Q vssd1 vssd1 vccd1 vccd1 _20902_/C sky130_fd_sc_hd__inv_2
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_366 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22632_ _22537_/X _22540_/Y _22615_/B vssd1 vssd1 vccd1 vccd1 _22632_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13432__A1 _13732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14167__B _15019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22563_ _13547_/A _22059_/X _22635_/A vssd1 vssd1 vccd1 vccd1 _22563_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_55_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21514_ _21514_/A vssd1 vssd1 vccd1 vccd1 _21633_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22494_ _22501_/A _22501_/B _22500_/B _22500_/C vssd1 vssd1 vccd1 vccd1 _22499_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21978__B1_N _21861_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21445_ _21445_/A _21445_/B _21561_/A vssd1 vssd1 vccd1 vccd1 _21561_/B sky130_fd_sc_hd__nand3_2
XFILLER_163_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11600__A _18947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21376_ _21376_/A _21376_/B vssd1 vssd1 vccd1 vccd1 _21378_/B sky130_fd_sc_hd__nor2_1
XANTENNA__16134__B1 _15975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19871__A1 _16464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18674__A2 _19040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20913__A _21174_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16685__A1 _16683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20327_ _20327_/A _20329_/B vssd1 vssd1 vccd1 vccd1 _20330_/B sky130_fd_sc_hd__nor2_1
XFILLER_190_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23115_ _19261_/C input7/X _23123_/S vssd1 vssd1 vccd1 vccd1 _23116_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14911__A _14911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20258_ _20256_/X _20250_/Y _20257_/Y vssd1 vssd1 vccd1 vccd1 _20312_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__19623__A1 _19381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23046_ _23046_/A vssd1 vssd1 vccd1 vccd1 _23351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12171__A1 _11851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13527__A _22392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20189_ _20189_/A _20189_/B _20189_/C vssd1 vssd1 vccd1 vccd1 _20206_/A sky130_fd_sc_hd__nand3_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _14174_/Y _14177_/B _14121_/B _14756_/A vssd1 vssd1 vccd1 vccd1 _14766_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ _11916_/X _11958_/X _11961_/Y vssd1 vssd1 vccd1 vccd1 _12189_/A sky130_fd_sc_hd__o21ai_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _13701_/A _21778_/D _13701_/C vssd1 vssd1 vccd1 vccd1 _13701_/Y sky130_fd_sc_hd__nand3_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _23402_/Q _14672_/X _14677_/X _23434_/Q _14680_/X vssd1 vssd1 vccd1 vccd1
+ _14681_/X sky130_fd_sc_hd__a221o_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11893_ _15718_/A vssd1 vssd1 vccd1 vccd1 _19165_/C sky130_fd_sc_hd__buf_2
XFILLER_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16420_ _16472_/A _16472_/B vssd1 vssd1 vccd1 vccd1 _16420_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13632_ _13632_/A vssd1 vssd1 vccd1 vccd1 _13632_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18772__B _18966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_591 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16351_ _16771_/B _16771_/C vssd1 vssd1 vccd1 vccd1 _16351_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13563_ _13563_/A _22035_/C _13563_/C vssd1 vssd1 vccd1 vccd1 _13563_/X sky130_fd_sc_hd__and3_1
XFILLER_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22294__B _22476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ _15409_/A _15363_/A _15419_/A vssd1 vssd1 vccd1 vccd1 _15302_/X sky130_fd_sc_hd__and3_1
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19070_ _18882_/B _18931_/X _19071_/A _19069_/Y vssd1 vssd1 vccd1 vccd1 _19075_/B
+ sky130_fd_sc_hd__o211ai_4
X_12514_ _16795_/C _12514_/B vssd1 vssd1 vccd1 vccd1 _17594_/A sky130_fd_sc_hd__nand2_2
XFILLER_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16282_ _16282_/A _16282_/B _16282_/C vssd1 vssd1 vccd1 vccd1 _16983_/B sky130_fd_sc_hd__nand3_1
XANTENNA__17388__B _19675_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13494_ _13555_/A _13494_/B _13494_/C vssd1 vssd1 vccd1 vccd1 _13494_/Y sky130_fd_sc_hd__nand3b_2
XANTENNA__16373__B1 _18461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17570__C1 _20317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16292__B _17974_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18021_ _18017_/B _17896_/C _18014_/Y vssd1 vssd1 vccd1 vccd1 _18022_/D sky130_fd_sc_hd__a21o_1
XANTENNA__23464__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15233_ _15233_/A _15233_/B _15233_/C vssd1 vssd1 vccd1 vccd1 _15233_/Y sky130_fd_sc_hd__nand3_1
X_12445_ _12445_/A _18497_/A _12445_/C vssd1 vssd1 vccd1 vccd1 _12445_/Y sky130_fd_sc_hd__nand3_1
XFILLER_154_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22997__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16125__B1 _16124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15164_ _15164_/A _15164_/B vssd1 vssd1 vccd1 vccd1 _15164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12376_ _11844_/A _12355_/A _12355_/B _12375_/X _11682_/Y vssd1 vssd1 vccd1 vccd1
+ _12376_/X sky130_fd_sc_hd__a311o_1
XFILLER_5_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1054 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14115_ _14172_/A _14172_/B vssd1 vssd1 vccd1 vccd1 _14115_/Y sky130_fd_sc_hd__nand2_4
XFILLER_113_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19972_ _19972_/A vssd1 vssd1 vccd1 vccd1 _20058_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15095_ _15099_/B vssd1 vssd1 vccd1 vccd1 _15095_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18923_ _19107_/B _19107_/C _19108_/A vssd1 vssd1 vccd1 vccd1 _18925_/B sky130_fd_sc_hd__nand3b_1
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14046_ _14588_/A _14050_/A _14061_/A _14120_/B vssd1 vssd1 vccd1 vccd1 _14858_/A
+ sky130_fd_sc_hd__o31a_2
XANTENNA_output76_A _14561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_850 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18854_ _11774_/A _11774_/B _12464_/Y _11961_/Y vssd1 vssd1 vccd1 vccd1 _18854_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_39_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18947__B _18947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17805_ _17805_/A _17805_/B vssd1 vssd1 vccd1 vccd1 _17805_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18785_ _18785_/A _18880_/B vssd1 vssd1 vccd1 vccd1 _18785_/Y sky130_fd_sc_hd__nand2_1
X_15997_ _16000_/A _15990_/Y _15996_/Y vssd1 vssd1 vccd1 vccd1 _16248_/A sky130_fd_sc_hd__o21ai_4
XFILLER_95_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23174__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22469__B _22553_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17736_ _17736_/A vssd1 vssd1 vccd1 vccd1 _17840_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14948_ _14931_/Y _14932_/X _14945_/C vssd1 vssd1 vccd1 vccd1 _14948_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12465__A2 _11931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22921__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15371__B _15371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17667_ _17667_/A _17667_/B vssd1 vssd1 vccd1 vccd1 _17670_/C sky130_fd_sc_hd__nand2_1
X_14879_ _14879_/A _14879_/B _14879_/C vssd1 vssd1 vccd1 vccd1 _14889_/B sky130_fd_sc_hd__nand3_1
XFILLER_36_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19406_ _19406_/A _19422_/B vssd1 vssd1 vccd1 vccd1 _19408_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16600__B2 _16319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16618_ _16153_/B _16617_/X _16614_/Y _19703_/C _16027_/D vssd1 vssd1 vccd1 vccd1
+ _16837_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_23_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17598_ _17960_/A _18093_/A vssd1 vssd1 vccd1 vccd1 _17598_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19337_ _19709_/A vssd1 vssd1 vccd1 vccd1 _19966_/A sky130_fd_sc_hd__clkbuf_2
X_16549_ _16549_/A _16549_/B _16549_/C _16549_/D vssd1 vssd1 vccd1 vccd1 _16549_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_188_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11976__A1 _11902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13900__A _14188_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19268_ _19275_/A _19275_/B _19275_/C vssd1 vssd1 vccd1 vccd1 _19268_/X sky130_fd_sc_hd__and3_1
XFILLER_176_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_514 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18219_ _18272_/A _19425_/C _20212_/D _18219_/D vssd1 vssd1 vccd1 vccd1 _18279_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_163_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19199_ _19662_/C _19543_/A _20062_/B _19199_/D vssd1 vssd1 vccd1 vccd1 _19201_/A
+ sky130_fd_sc_hd__nand4_4
XANTENNA__19302__B1 _19172_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22988__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21230_ _21119_/A _21119_/B _21119_/C _21123_/C vssd1 vssd1 vccd1 vccd1 _21236_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18656__A2 _12006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21829__A _21829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16930__B _16930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21161_ _21268_/A _21271_/B vssd1 vssd1 vccd1 vccd1 _21161_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21548__B _21548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20112_ _20112_/A _20112_/B vssd1 vssd1 vccd1 vccd1 _20185_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23466__D _23478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21092_ _20979_/A _20984_/B _20984_/C vssd1 vssd1 vccd1 vccd1 _21092_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__22204__A3 _22208_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20043_ _20043_/A _20043_/B vssd1 vssd1 vccd1 vccd1 _20043_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17761__B _17761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23165__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_683 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21994_ _21994_/A _21994_/B vssd1 vssd1 vccd1 vccd1 _21994_/Y sky130_fd_sc_hd__nand2_2
XFILLER_2_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22912__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19969__A _19969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ _20945_/A _20945_/B _20945_/C vssd1 vssd1 vccd1 vccd1 _20984_/B sky130_fd_sc_hd__nand3_4
XFILLER_198_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_388 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _20751_/Y _20754_/X _20756_/Y vssd1 vssd1 vccd1 vccd1 _20877_/A sky130_fd_sc_hd__a21o_1
XFILLER_183_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22615_ _22615_/A _22615_/B vssd1 vssd1 vccd1 vccd1 _22619_/B sky130_fd_sc_hd__nand2_1
XFILLER_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23595_ _23598_/CLK _23595_/D vssd1 vssd1 vccd1 vccd1 _23595_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_179_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13810__A _22014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22545__D _22663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22546_ _22545_/B _22545_/C _22754_/A _22484_/X vssd1 vssd1 vccd1 vccd1 _22548_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_10_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22477_ _21997_/X _22059_/X _22368_/Y vssd1 vssd1 vccd1 vccd1 _22477_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__12426__A _15718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22979__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ _12540_/B _12532_/B _12203_/Y _12220_/Y vssd1 vssd1 vccd1 vccd1 _12230_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_120_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21428_ _21455_/B vssd1 vssd1 vccd1 vccd1 _21428_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19844__A1 _20209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16840__B _18755_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12161_ _12491_/A _12491_/B _12217_/B _12217_/C vssd1 vssd1 vccd1 vccd1 _12161_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_135_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21359_ _21359_/A _21359_/B vssd1 vssd1 vccd1 vccd1 _21359_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_956 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12092_ _18503_/D _19000_/B _18503_/C vssd1 vssd1 vccd1 vccd1 _12093_/A sky130_fd_sc_hd__nand3_1
XFILLER_1_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23029_ _23029_/A vssd1 vssd1 vccd1 vccd1 _23344_/D sky130_fd_sc_hd__clkbuf_1
X_15920_ _15920_/A _15920_/B _16667_/B _15920_/D vssd1 vssd1 vccd1 vccd1 _15921_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19072__A2 _18931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15175__C _15175_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17083__A1 _12518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15851_ _15941_/A _15943_/A _15943_/B vssd1 vssd1 vccd1 vccd1 _15879_/A sky130_fd_sc_hd__nand3_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23156__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16830__A1 _12222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ _14975_/C _14911_/A _15301_/A _14448_/A vssd1 vssd1 vccd1 vccd1 _14802_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_36_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18570_ _18912_/B _19090_/C vssd1 vssd1 vccd1 vccd1 _18570_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__21193__B _21493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15782_ _15721_/X _15781_/Y _15719_/B vssd1 vssd1 vccd1 vccd1 _15782_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12994_ _20775_/D vssd1 vssd1 vccd1 vccd1 _20886_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22903__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17521_ _16994_/C _16994_/D _16994_/A vssd1 vssd1 vccd1 vccd1 _17524_/A sky130_fd_sc_hd__a21oi_1
X_14733_ _23260_/A vssd1 vssd1 vccd1 vccd1 _23256_/A sky130_fd_sc_hd__clkbuf_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ _23591_/Q vssd1 vssd1 vccd1 vccd1 _16800_/A sky130_fd_sc_hd__buf_2
XFILLER_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17433_/X _17437_/X _17445_/A _20062_/C _17440_/A vssd1 vssd1 vccd1 vccd1
+ _17453_/C sky130_fd_sc_hd__o2111ai_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _23335_/Q _14636_/X _14642_/X _23303_/Q _14657_/X vssd1 vssd1 vccd1 vccd1
+ _14664_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11876_ _18675_/B vssd1 vssd1 vccd1 vccd1 _19040_/A sky130_fd_sc_hd__buf_2
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16403_ _16403_/A _16403_/B _16403_/C vssd1 vssd1 vccd1 vccd1 _16405_/A sky130_fd_sc_hd__nand3_2
X_13615_ _13615_/A vssd1 vssd1 vccd1 vccd1 _13616_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17383_ _17382_/B _17533_/A _17382_/D _17382_/A vssd1 vssd1 vccd1 vccd1 _17384_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14595_ _14070_/X _14545_/A _14539_/X _12121_/B vssd1 vssd1 vccd1 vccd1 _14595_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19122_ _19118_/Y _19119_/Y _19530_/A _19121_/X _19705_/A vssd1 vssd1 vccd1 vccd1
+ _19125_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_125_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16334_ _16066_/A _16408_/A _15852_/X _16071_/Y vssd1 vssd1 vccd1 vccd1 _16335_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13546_ _13540_/Y _13543_/Y _13544_/Y _13545_/Y vssd1 vssd1 vccd1 vccd1 _13697_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_185_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19053_ _18828_/Y _18840_/Y _18846_/A _18875_/B vssd1 vssd1 vccd1 vccd1 _19055_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_9_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16897__A1 _16054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16265_ _16347_/A _16265_/B vssd1 vssd1 vccd1 vccd1 _16266_/C sky130_fd_sc_hd__nand2_2
XFILLER_187_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13477_ _13477_/A vssd1 vssd1 vccd1 vccd1 _13477_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18004_ _17958_/A _17752_/X _18211_/B _17611_/X vssd1 vssd1 vccd1 vccd1 _18004_/X
+ sky130_fd_sc_hd__o22a_1
X_15216_ _15144_/B _15144_/A _15063_/A _15066_/Y vssd1 vssd1 vccd1 vccd1 _15286_/C
+ sky130_fd_sc_hd__o22ai_4
XFILLER_127_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12428_ _19019_/C _18445_/B vssd1 vssd1 vccd1 vccd1 _12428_/Y sky130_fd_sc_hd__nand2_1
X_16196_ _16661_/A vssd1 vssd1 vccd1 vccd1 _17631_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_142_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15147_ _15066_/Y _15145_/X _15146_/Y vssd1 vssd1 vccd1 vccd1 _15220_/C sky130_fd_sc_hd__o21a_1
X_12359_ _14735_/A _19534_/C _12355_/Y _12358_/X vssd1 vssd1 vccd1 vccd1 _12363_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19955_ _19847_/X _19848_/Y _20079_/A _19659_/Y vssd1 vssd1 vccd1 vccd1 _19955_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_15078_ _15195_/B _14068_/X _14069_/X _15077_/X vssd1 vssd1 vccd1 vccd1 _15078_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18958__A _19900_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12135__A1 _12130_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17862__A _20142_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18906_ _18900_/X _18901_/X _18903_/Y _18905_/X vssd1 vssd1 vccd1 vccd1 _18907_/A
+ sky130_fd_sc_hd__o211ai_1
X_14029_ _14029_/A _14086_/A _14029_/C vssd1 vssd1 vccd1 vccd1 _14029_/X sky130_fd_sc_hd__and3_2
X_19886_ _19827_/A _19830_/A _19882_/X vssd1 vssd1 vccd1 vccd1 _19888_/A sky130_fd_sc_hd__a21o_1
XFILLER_171_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18837_ _19703_/D vssd1 vssd1 vccd1 vccd1 _19543_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16478__A _17285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18768_ _12308_/A _17443_/A _17444_/A _19113_/C _12066_/A vssd1 vssd1 vccd1 vccd1
+ _18768_/X sky130_fd_sc_hd__a32o_1
XFILLER_64_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17719_ _12088_/A _17644_/X _17467_/X _17760_/A vssd1 vssd1 vccd1 vccd1 _17719_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17377__A2 _18059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18699_ _18751_/A _18751_/B _18751_/C vssd1 vssd1 vccd1 vccd1 _18706_/A sky130_fd_sc_hd__nand3_1
X_20730_ _20728_/Y _20729_/Y _20716_/C _20716_/A vssd1 vssd1 vccd1 vccd1 _20730_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_91_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20661_ _21046_/A _20894_/B vssd1 vssd1 vccd1 vccd1 _20662_/B sky130_fd_sc_hd__nand2_1
XFILLER_91_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14726__A _23596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22400_ _22400_/A _22400_/B _22412_/A _22400_/D vssd1 vssd1 vccd1 vccd1 _22401_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20592_ _21008_/B vssd1 vssd1 vccd1 vccd1 _20593_/C sky130_fd_sc_hd__clkbuf_2
X_23380_ _23381_/CLK _23380_/D vssd1 vssd1 vccd1 vccd1 _23380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_823 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22331_ _22330_/Y _22210_/Y _22225_/A _22232_/X vssd1 vssd1 vccd1 vccd1 _22333_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__12136__A1_N _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__C _18755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22262_ _21829_/A _13431_/X _22261_/Y vssd1 vssd1 vccd1 vccd1 _22434_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__18629__A2 _18490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22381__C _22381_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21213_ _21217_/A _21218_/B _21218_/C vssd1 vssd1 vccd1 vccd1 _21319_/B sky130_fd_sc_hd__nand3_2
XFILLER_118_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19029__A _19029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22193_ _22160_/Y _22192_/Y _22182_/X vssd1 vssd1 vccd1 vccd1 _22193_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21144_ _23564_/Q _21144_/B vssd1 vssd1 vccd1 vccd1 _21144_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18868__A _18868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21075_ _21063_/Y _21066_/Y _20969_/A _12722_/X vssd1 vssd1 vccd1 vccd1 _21163_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__19054__A2 _19048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20026_ _20207_/D vssd1 vssd1 vccd1 vccd1 _20196_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21977_ _21975_/Y _21977_/B vssd1 vssd1 vccd1 vccd1 _21979_/A sky130_fd_sc_hd__and2b_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15442__D _15442_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11720_/A _11724_/A _11694_/X _11860_/C _11960_/B vssd1 vssd1 vccd1 vccd1
+ _16364_/A sky130_fd_sc_hd__o311ai_4
XANTENNA__20372__A1 _20371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ _21281_/A _21282_/A vssd1 vssd1 vccd1 vccd1 _21592_/A sky130_fd_sc_hd__nand2_2
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20638__A _23296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _23388_/Q vssd1 vssd1 vccd1 vccd1 _11665_/A sky130_fd_sc_hd__clkbuf_4
X_20859_ _20858_/Y _20724_/A _20736_/A _20867_/A _20867_/B vssd1 vssd1 vccd1 vccd1
+ _20859_/Y sky130_fd_sc_hd__a32oi_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13400_ _21883_/A _13600_/C _21883_/C vssd1 vssd1 vccd1 vccd1 _13400_/Y sky130_fd_sc_hd__nand3_4
XFILLER_179_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16328__B1 _16325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14380_ _14492_/C _14380_/B vssd1 vssd1 vccd1 vccd1 _14380_/Y sky130_fd_sc_hd__nor2_1
X_23578_ _23578_/CLK _23578_/D vssd1 vssd1 vccd1 vccd1 _23578_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21321__B1 _21215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11592_ _11634_/B vssd1 vssd1 vccd1 vccd1 _16807_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__18261__B1_N _23532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13331_ _13660_/A vssd1 vssd1 vccd1 vccd1 _13701_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_823 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22529_ _22529_/A _22629_/A _22629_/B vssd1 vssd1 vccd1 vccd1 _22530_/A sky130_fd_sc_hd__or3b_1
XFILLER_155_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_931 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16050_ _16372_/A _17226_/D _16046_/Y _16757_/A vssd1 vssd1 vccd1 vccd1 _16094_/A
+ sky130_fd_sc_hd__a22oi_4
X_13262_ _13483_/B _21739_/A _23322_/Q vssd1 vssd1 vccd1 vccd1 _13766_/A sky130_fd_sc_hd__a21o_2
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15001_ _15001_/A vssd1 vssd1 vccd1 vccd1 _15001_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11995__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ _12093_/X _12151_/Y _12107_/X _19648_/A _18952_/D vssd1 vssd1 vccd1 vccd1
+ _12216_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_68_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ _13171_/Y _13174_/B _13174_/A vssd1 vssd1 vccd1 vccd1 _13193_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ _12144_/A vssd1 vssd1 vccd1 vccd1 _16437_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_97_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14106__A2 _14015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18778__A _18778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12603__B _21036_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19740_ _19740_/A _19740_/B _19880_/B _19893_/B vssd1 vssd1 vccd1 vccd1 _19742_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__15854__A2 _16370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12075_ _15860_/D vssd1 vssd1 vccd1 vccd1 _19703_/C sky130_fd_sc_hd__buf_2
X_16952_ _16944_/X _16949_/Y _17184_/A vssd1 vssd1 vccd1 vccd1 _16952_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__21916__B _22045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15903_ _15899_/X _16209_/A _15902_/Y vssd1 vssd1 vccd1 vccd1 _15907_/A sky130_fd_sc_hd__o21ai_1
X_19671_ _17643_/X _19668_/X _19669_/X _19670_/X vssd1 vssd1 vccd1 vccd1 _19672_/C
+ sky130_fd_sc_hd__o31a_1
X_16883_ _16864_/A _16890_/B _16880_/X _16871_/X vssd1 vssd1 vccd1 vccd1 _16894_/D
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18622_ _18518_/B _18520_/B _18518_/A vssd1 vssd1 vccd1 vccd1 _18622_/X sky130_fd_sc_hd__a21bo_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _15834_/A vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _18902_/B _18553_/B vssd1 vssd1 vccd1 vccd1 _18554_/C sky130_fd_sc_hd__nor2_1
XFILLER_46_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15765_ _15765_/A vssd1 vssd1 vccd1 vccd1 _16447_/A sky130_fd_sc_hd__buf_4
X_12977_ _12977_/A _12977_/B _12977_/C vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__nand3_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _17513_/A _17513_/B _17513_/C vssd1 vssd1 vccd1 vccd1 _17504_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18944__C _18944_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11928_ _12474_/A vssd1 vssd1 vccd1 vccd1 _18859_/D sky130_fd_sc_hd__buf_2
X_14716_ _23380_/Q _14635_/A _14715_/X vssd1 vssd1 vccd1 vccd1 _14716_/X sky130_fd_sc_hd__o21a_1
X_18484_ _18484_/A vssd1 vssd1 vccd1 vccd1 _18484_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15696_ _15686_/A _15686_/B _15678_/Y vssd1 vssd1 vccd1 vccd1 _15698_/A sky130_fd_sc_hd__a21oi_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16031__A2 _16058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17435_ _17435_/A vssd1 vssd1 vccd1 vccd1 _17435_/X sky130_fd_sc_hd__buf_2
X_14647_ _14647_/A vssd1 vssd1 vccd1 vccd1 _14647_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11859_ _11720_/A _11644_/C _11694_/X _11733_/Y _16796_/A vssd1 vssd1 vccd1 vccd1
+ _12017_/A sky130_fd_sc_hd__o311a_1
XFILLER_198_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17366_ _17200_/B _17195_/Y _17203_/Y vssd1 vssd1 vccd1 vccd1 _17369_/C sky130_fd_sc_hd__o21ai_2
XFILLER_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14578_ _13304_/X _14550_/X _14539_/X _12245_/X _14577_/X vssd1 vssd1 vccd1 vccd1
+ _14578_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19105_ _19105_/A _19105_/B vssd1 vssd1 vccd1 vccd1 _23523_/D sky130_fd_sc_hd__nor2_1
XFILLER_9_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16317_ _16384_/A _16355_/A _16316_/Y vssd1 vssd1 vccd1 vccd1 _16318_/A sky130_fd_sc_hd__o21ai_1
X_13529_ _21919_/C vssd1 vssd1 vccd1 vccd1 _22380_/C sky130_fd_sc_hd__clkbuf_2
X_17297_ _17477_/A _17477_/B _17297_/C _17297_/D vssd1 vssd1 vccd1 vccd1 _17299_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20130__A4 _20369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23065__A0 _14883_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19036_ _19036_/A _19036_/B vssd1 vssd1 vccd1 vccd1 _19052_/B sky130_fd_sc_hd__nand2_2
XFILLER_146_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16248_ _16248_/A _16248_/B _16248_/C _16248_/D vssd1 vssd1 vccd1 vccd1 _16268_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19494__D _19494_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12356__A1 _14735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16179_ _16010_/X _16179_/B _16179_/C vssd1 vssd1 vccd1 vccd1 _16254_/B sky130_fd_sc_hd__nand3b_4
XFILLER_115_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18087__A3 _18016_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15808__C _17860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17295__A1 _17104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19938_ _19889_/A _19889_/B _19889_/C _19897_/C vssd1 vssd1 vccd1 vccd1 _19938_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_99_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19869_ _20142_/B vssd1 vssd1 vccd1 vccd1 _20269_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_29_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21545__C _21592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21900_ _23328_/Q _23329_/Q vssd1 vssd1 vccd1 vccd1 _22141_/B sky130_fd_sc_hd__nor2_1
XFILLER_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22880_ _22881_/B _22887_/B _23285_/Q vssd1 vssd1 vccd1 vccd1 _22891_/A sky130_fd_sc_hd__a21bo_1
XFILLER_56_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13344__B _13377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21831_ _22510_/B vssd1 vssd1 vccd1 vccd1 _22667_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__21842__A _21842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22879__B1 _22878_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18011__A3 _17391_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12292__B1 _12238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21762_ _21923_/A _22064_/C _21919_/C _21924_/A vssd1 vssd1 vccd1 vccd1 _21762_/Y
+ sky130_fd_sc_hd__nand4_2
XANTENNA__20458__A _23560_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_926 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23501_ _23510_/CLK _23501_/D vssd1 vssd1 vccd1 vccd1 _23501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20713_ _20728_/A _20713_/B vssd1 vssd1 vccd1 vccd1 _20714_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21693_ _21665_/A _21631_/B _21631_/C _21631_/A _21542_/X vssd1 vssd1 vccd1 vccd1
+ _21698_/A sky130_fd_sc_hd__a41o_1
XANTENNA__14033__A1 _14015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14456__A _14819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23432_ _23432_/CLK _23432_/D vssd1 vssd1 vccd1 vccd1 _23432_/Q sky130_fd_sc_hd__dfxtp_1
X_20644_ _20917_/A vssd1 vssd1 vccd1 vccd1 _20921_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__19966__B _20062_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23363_ _23363_/CLK _23363_/D vssd1 vssd1 vccd1 vccd1 _23363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20575_ _20589_/A _20736_/A _20589_/C vssd1 vssd1 vccd1 vccd1 _20575_/Y sky130_fd_sc_hd__nand3_1
XFILLER_20_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22392__B _22392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23056__A0 _14031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22314_ _22314_/A _22314_/B vssd1 vssd1 vccd1 vccd1 _22323_/C sky130_fd_sc_hd__nor2_1
XFILLER_191_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23294_ _23295_/CLK _23294_/D vssd1 vssd1 vccd1 vccd1 _23294_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_164_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22245_ _21981_/A _21981_/B _21981_/C _22118_/Y vssd1 vssd1 vccd1 vccd1 _22246_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_164_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22176_ _22176_/A vssd1 vssd1 vccd1 vccd1 _22290_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21127_ _20995_/A _20995_/B _20995_/C _21130_/A vssd1 vssd1 vccd1 vccd1 _21127_/Y
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__19027__A2 _19485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21058_ _21084_/A _21212_/A _21084_/C _21057_/Y _20947_/A vssd1 vssd1 vccd1 vccd1
+ _21089_/A sky130_fd_sc_hd__a32oi_4
XFILLER_115_1052 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18786__A1 _18868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1003 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12900_ _12900_/A _13034_/A _13044_/A _13044_/B vssd1 vssd1 vccd1 vccd1 _12901_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20009_ _19937_/Y _19896_/B _19897_/B vssd1 vssd1 vccd1 vccd1 _20012_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__16549__C _16549_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13880_ _14430_/D vssd1 vssd1 vccd1 vccd1 _14459_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_143_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _13177_/B _13177_/C _12827_/A vssd1 vssd1 vccd1 vccd1 _12833_/B sky130_fd_sc_hd__a21oi_2
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15750__A _16593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15550_ _15522_/A _15547_/Y _15558_/C vssd1 vssd1 vccd1 vccd1 _15552_/A sky130_fd_sc_hd__o21bai_4
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _23452_/Q vssd1 vssd1 vccd1 vccd1 _12763_/A sky130_fd_sc_hd__inv_2
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_634 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20368__A _20368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_656 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14853_/A _14501_/B vssd1 vssd1 vccd1 vccd1 _14502_/A sky130_fd_sc_hd__and2_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11713_/A _11713_/B vssd1 vssd1 vccd1 vccd1 _16677_/A sky130_fd_sc_hd__nand2_1
X_15481_ _15460_/A _15460_/B _15458_/B vssd1 vssd1 vccd1 vccd1 _15499_/A sky130_fd_sc_hd__o21a_1
XFILLER_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12689_/X _12850_/B _12692_/Y vssd1 vssd1 vccd1 vccd1 _12694_/A sky130_fd_sc_hd__a21oi_2
XFILLER_70_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17220_ _17220_/A _17220_/B _17220_/C vssd1 vssd1 vccd1 vccd1 _17220_/X sky130_fd_sc_hd__and3_1
X_14432_ _14436_/A _14436_/C _14436_/B vssd1 vssd1 vccd1 vccd1 _14465_/A sky130_fd_sc_hd__a21o_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _23586_/Q _23584_/Q _11644_/C _11739_/B vssd1 vssd1 vccd1 vccd1 _15956_/A
+ sky130_fd_sc_hd__nor4_2
XFILLER_187_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17151_ _17151_/A _17151_/B _17151_/C vssd1 vssd1 vccd1 vccd1 _17152_/B sky130_fd_sc_hd__nand3_2
XFILLER_196_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14363_ _14353_/X _14357_/X _14358_/Y _14362_/Y vssd1 vssd1 vccd1 vccd1 _14414_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__20648__A2 _12722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11575_ _11739_/A vssd1 vssd1 vccd1 vccd1 _12071_/A sky130_fd_sc_hd__clkbuf_2
Xinput16 wb_dat_i[18] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_2
Xinput27 wb_dat_i[28] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_2
XFILLER_195_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16102_ _16089_/X _16090_/X _16072_/Y _16097_/Y vssd1 vssd1 vccd1 vccd1 _16425_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16316__A3 _16451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23047__A0 _13977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput38 wb_dat_i[9] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_4
X_13314_ _23476_/Q vssd1 vssd1 vccd1 vccd1 _21925_/B sky130_fd_sc_hd__clkbuf_2
X_17082_ _12086_/A _16451_/B _16451_/C _17077_/A vssd1 vssd1 vccd1 vccd1 _17082_/X
+ sky130_fd_sc_hd__o31a_1
Xinput49 x[6] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_4
XFILLER_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14327__A2 _14203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14294_ _14294_/A _14294_/B vssd1 vssd1 vccd1 vccd1 _14310_/B sky130_fd_sc_hd__nand2_1
XFILLER_143_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16033_ _16033_/A vssd1 vssd1 vccd1 vccd1 _16033_/X sky130_fd_sc_hd__buf_4
X_13245_ _13523_/A _22476_/C _13680_/A _13247_/A vssd1 vssd1 vccd1 vccd1 _13249_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19266__A2 _20368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13176_ _13176_/A _21182_/D _13176_/C vssd1 vssd1 vccd1 vccd1 _13176_/X sky130_fd_sc_hd__and3_1
XFILLER_151_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ _18444_/A vssd1 vssd1 vccd1 vccd1 _18645_/A sky130_fd_sc_hd__buf_2
X_17984_ _17994_/A _17994_/B _17992_/A vssd1 vssd1 vccd1 vccd1 _17984_/Y sky130_fd_sc_hd__nand3_1
XFILLER_97_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23564__D _23564_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19723_ _19723_/A _19723_/B _19723_/C vssd1 vssd1 vccd1 vccd1 _19725_/B sky130_fd_sc_hd__nand3_1
X_12058_ _12204_/B vssd1 vssd1 vccd1 vccd1 _12059_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_16935_ _16935_/A vssd1 vssd1 vccd1 vccd1 _17166_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19654_ _19503_/X _19647_/Y _19650_/X _19653_/X vssd1 vssd1 vccd1 vccd1 _19654_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16866_ _16866_/A vssd1 vssd1 vccd1 vccd1 _17605_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__16788__B1 _16778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18605_ _18537_/Y _18932_/A _18599_/B _18599_/A vssd1 vssd1 vccd1 vccd1 _18605_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15817_ _15834_/A _16029_/B vssd1 vssd1 vccd1 vccd1 _15817_/Y sky130_fd_sc_hd__nand2_1
X_19585_ _19588_/B vssd1 vssd1 vccd1 vccd1 _19747_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16797_ _16808_/A _16808_/B _16796_/X vssd1 vssd1 vccd1 vccd1 _18947_/C sky130_fd_sc_hd__o21ai_4
XANTENNA__15082__D _15082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_995 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19132__A _19391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18536_ _11611_/A _11611_/B _12222_/X _12223_/X vssd1 vssd1 vccd1 vccd1 _18536_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15748_ _15729_/X _16187_/A _15662_/C vssd1 vssd1 vccd1 vccd1 _15749_/B sky130_fd_sc_hd__o21ai_4
XFILLER_93_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17201__A1 _16663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ _18649_/A _18469_/B _12410_/C _18998_/C _11754_/A vssd1 vssd1 vccd1 vccd1
+ _18483_/A sky130_fd_sc_hd__a41oi_4
XFILLER_34_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15679_ _16187_/A _15637_/D _15677_/Y _15678_/Y vssd1 vssd1 vccd1 vccd1 _15974_/C
+ sky130_fd_sc_hd__a31o_4
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17418_ _17429_/A vssd1 vssd1 vccd1 vccd1 _17485_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__12026__B1 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18398_ _18398_/A _18417_/A _18398_/C vssd1 vssd1 vccd1 vccd1 _18407_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12508__B _19543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17587__A _17587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17349_ _17187_/A _17192_/X _17187_/B vssd1 vssd1 vccd1 vccd1 _17351_/B sky130_fd_sc_hd__a21boi_1
XFILLER_14_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12227__C _12227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20360_ _20359_/C _20358_/Y _20359_/Y _20312_/B vssd1 vssd1 vccd1 vccd1 _20420_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_147_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12329__A1 _12346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19019_ _19327_/B _19019_/B _19019_/C vssd1 vssd1 vccd1 vccd1 _19019_/Y sky130_fd_sc_hd__nand3_1
X_20291_ _20295_/B _20295_/A vssd1 vssd1 vccd1 vccd1 _20291_/X sky130_fd_sc_hd__or2_1
XFILLER_161_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15538__C _15538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22030_ _22028_/Y _22141_/C _13486_/B vssd1 vssd1 vccd1 vccd1 _22030_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__21064__A2 _21061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22261__A1 _22139_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18849__C _18849_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18211__A _18211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17753__C _20055_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22013__A1 _13465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18768__A1 _12308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22932_ _20902_/B input13/X _22940_/S vssd1 vssd1 vccd1 vccd1 _22933_/A sky130_fd_sc_hd__mux2_1
XANTENNA__21772__B1 _22276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22863_ _22834_/A _22834_/B _22834_/C _22839_/A _22862_/Y vssd1 vssd1 vccd1 vccd1
+ _22865_/A sky130_fd_sc_hd__a311oi_1
XANTENNA__17991__A2 _18002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21814_ _21987_/B vssd1 vssd1 vccd1 vccd1 _22236_/A sky130_fd_sc_hd__clkinv_2
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22794_ _22237_/X _22754_/B _22791_/X _22792_/X vssd1 vssd1 vccd1 vccd1 _22797_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20619__C _21035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13802__B _13802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21745_ _21745_/A _21745_/B vssd1 vssd1 vccd1 vccd1 _22020_/B sky130_fd_sc_hd__nand2_2
XFILLER_52_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17743__A2 _17742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_795 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_946 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21676_ _21646_/A _21675_/Y _21673_/Y vssd1 vssd1 vccd1 vccd1 _21704_/C sky130_fd_sc_hd__o21ai_2
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23415_ _23416_/CLK _23415_/D vssd1 vssd1 vccd1 vccd1 _23415_/Q sky130_fd_sc_hd__dfxtp_1
X_20627_ _20502_/X _20504_/X _23448_/Q _20496_/X vssd1 vssd1 vccd1 vccd1 _20627_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_149_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11776__C1 _11747_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23346_ _23378_/CLK _23346_/D vssd1 vssd1 vccd1 vccd1 _23346_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16703__B1 _16662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20558_ _13079_/B _13049_/A _20556_/X _20557_/Y vssd1 vssd1 vccd1 vccd1 _20578_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_138_54 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23277_ _23510_/CLK _23277_/D vssd1 vssd1 vccd1 vccd1 _23277_/Q sky130_fd_sc_hd__dfxtp_1
X_20489_ _21493_/A _21493_/B _20784_/C vssd1 vssd1 vccd1 vccd1 _20490_/B sky130_fd_sc_hd__and3_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13030_ _12725_/A _12854_/Y _13002_/Y _13003_/Y vssd1 vssd1 vccd1 vccd1 _13030_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22228_ _22086_/Y _22119_/X _22093_/D _22225_/Y _22227_/Y vssd1 vssd1 vccd1 vccd1
+ _22228_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_191_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13532__A3 _13527_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15809__A2 _17409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22159_ _22267_/A _22268_/A _22159_/C vssd1 vssd1 vccd1 vccd1 _22271_/A sky130_fd_sc_hd__nand3_2
XFILLER_65_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16482__A2 _16458_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A wb_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14981_ _15353_/A _15353_/B _15010_/A vssd1 vssd1 vccd1 vccd1 _14981_/X sky130_fd_sc_hd__and3_1
XANTENNA__18759__A1 _12324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17416__D1 _17723_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13265__A _23474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16720_ _16010_/X _16176_/Y _16256_/Y _16719_/Y vssd1 vssd1 vccd1 vccd1 _16720_/Y
+ sky130_fd_sc_hd__o22ai_4
X_13932_ _15353_/A _15353_/B _14312_/D _14374_/D vssd1 vssd1 vccd1 vccd1 _13933_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_101_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16651_ _16646_/Y _16647_/X _16648_/Y _16650_/Y vssd1 vssd1 vccd1 vccd1 _16651_/Y
+ sky130_fd_sc_hd__o22ai_2
X_13863_ _21832_/A _22800_/A vssd1 vssd1 vccd1 vccd1 _13863_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_835 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12814_ _13151_/A _12785_/X _12815_/C _12816_/B _12816_/C vssd1 vssd1 vccd1 vccd1
+ _12817_/A sky130_fd_sc_hd__o32a_1
X_15602_ _23422_/Q vssd1 vssd1 vccd1 vccd1 _15642_/A sky130_fd_sc_hd__inv_2
X_19370_ _12246_/Y _12247_/Y _19709_/B _19709_/C vssd1 vssd1 vccd1 vccd1 _19371_/B
+ sky130_fd_sc_hd__o211a_1
X_13794_ _13453_/A _13410_/A _13615_/A _21916_/A _13793_/Y vssd1 vssd1 vccd1 vccd1
+ _13794_/Y sky130_fd_sc_hd__o221ai_4
X_16582_ _16582_/A _16582_/B _16582_/C vssd1 vssd1 vccd1 vccd1 _16774_/B sky130_fd_sc_hd__nand3_2
X_18321_ _18207_/X _18208_/X _18320_/Y vssd1 vssd1 vccd1 vccd1 _18395_/A sky130_fd_sc_hd__o21ai_1
XFILLER_16_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15533_ _15533_/A vssd1 vssd1 vccd1 vccd1 _15538_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _12997_/A vssd1 vssd1 vccd1 vccd1 _20473_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _18252_/A _18252_/B vssd1 vssd1 vccd1 vccd1 _18254_/B sky130_fd_sc_hd__nor2_1
XFILLER_148_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464_ _15429_/A _15429_/B _15463_/Y vssd1 vssd1 vccd1 vccd1 _15467_/A sky130_fd_sc_hd__o21ai_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15745__A1 _15742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12875_/C _12712_/A _12675_/X vssd1 vssd1 vccd1 vccd1 _12677_/A sky130_fd_sc_hd__a21o_1
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17203_ _17200_/B _17195_/Y _17202_/Y vssd1 vssd1 vccd1 vccd1 _17203_/Y sky130_fd_sc_hd__a21oi_2
X_14415_ _14418_/A _14415_/B _14415_/C vssd1 vssd1 vccd1 vccd1 _14495_/A sky130_fd_sc_hd__nand3b_1
XFILLER_128_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11627_ _12510_/A _16619_/A _16815_/A vssd1 vssd1 vccd1 vccd1 _12175_/A sky130_fd_sc_hd__a21o_1
XANTENNA__21818__A1 _22420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18183_ _18110_/B _18110_/A _18185_/C _18185_/B _18108_/A vssd1 vssd1 vccd1 vccd1
+ _18186_/A sky130_fd_sc_hd__o221a_1
XFILLER_156_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15395_ _15395_/A _15395_/B _15395_/C vssd1 vssd1 vccd1 vccd1 _15395_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__19487__A2 _19173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_951 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17134_ _17134_/A _17134_/B _17134_/C vssd1 vssd1 vccd1 vccd1 _17156_/B sky130_fd_sc_hd__and3_1
X_14346_ _14361_/C _14361_/A _14347_/C vssd1 vssd1 vccd1 vccd1 _14346_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21294__A2 _21061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22491__A1 _21891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17065_ _17068_/A _17069_/A _17070_/A vssd1 vssd1 vccd1 vccd1 _17077_/A sky130_fd_sc_hd__o21ai_2
XFILLER_13_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14277_ _14039_/A _14260_/A _15225_/C _14457_/A _14049_/Y vssd1 vssd1 vccd1 vccd1
+ _14279_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_195_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16016_ _15949_/X _16015_/Y _16002_/B _16006_/Y vssd1 vssd1 vccd1 vccd1 _16017_/C
+ sky130_fd_sc_hd__o211ai_1
X_13228_ _23320_/Q vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14720__A2 _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22794__A2 _22754_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21376__B _21376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _20563_/A _20563_/B _21177_/B _13158_/A _13156_/A vssd1 vssd1 vccd1 vccd1
+ _13159_/X sky130_fd_sc_hd__a32o_1
XFILLER_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _17967_/A vssd1 vssd1 vccd1 vccd1 _18080_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18966__A _18966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19706_ _19819_/A _19820_/A _19218_/X _18003_/A vssd1 vssd1 vccd1 vccd1 _19831_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16918_ _23428_/Q vssd1 vssd1 vccd1 vccd1 _16918_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17898_ _18079_/A _19957_/A _20164_/C _17898_/D vssd1 vssd1 vccd1 vccd1 _17898_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__13606__C _23471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19637_ _18919_/X _19443_/B _19442_/A _19442_/B vssd1 vssd1 vccd1 vccd1 _19637_/Y
+ sky130_fd_sc_hd__o211ai_1
X_16849_ _16848_/Y _16828_/Y _16841_/B vssd1 vssd1 vccd1 vccd1 _16849_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19568_ _19568_/A vssd1 vssd1 vccd1 vccd1 _19573_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19175__A1 _18993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18519_ _18523_/A _18529_/A _18516_/X _18518_/X vssd1 vssd1 vccd1 vccd1 _18519_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
X_19499_ _19499_/A vssd1 vssd1 vccd1 vccd1 _20209_/A sky130_fd_sc_hd__buf_2
XFILLER_178_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21530_ _21616_/A _21617_/A _21614_/D _21529_/X vssd1 vssd1 vccd1 vccd1 _21541_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_167_918 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23112__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21461_ _21463_/C _21463_/D vssd1 vssd1 vccd1 vccd1 _21461_/Y sky130_fd_sc_hd__nand2_1
X_23200_ _15664_/A input35/X _23206_/S vssd1 vssd1 vccd1 vccd1 _23201_/A sky130_fd_sc_hd__mux2_1
XANTENNA__23469__D _23481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20412_ _20431_/B _20412_/B vssd1 vssd1 vccd1 vccd1 _20414_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21392_ _21317_/Y _21318_/X _21319_/Y _21311_/A _21327_/C vssd1 vssd1 vccd1 vccd1
+ _21392_/X sky130_fd_sc_hd__a32o_1
XFILLER_88_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23131_ _23131_/A vssd1 vssd1 vccd1 vccd1 _23389_/D sky130_fd_sc_hd__clkbuf_1
X_20343_ _20343_/A vssd1 vssd1 vccd1 vccd1 _20343_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16161__A1 _15971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23062_ _14188_/A input38/X _23062_/S vssd1 vssd1 vccd1 vccd1 _23063_/A sky130_fd_sc_hd__mux2_1
X_20274_ _20274_/A _20274_/B _20274_/C _20400_/A vssd1 vssd1 vccd1 vccd1 _20400_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_162_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20471__A _21493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20245__B1 _20183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22013_ _13465_/A _22484_/A _22012_/Y vssd1 vssd1 vccd1 vccd1 _22130_/A sky130_fd_sc_hd__o21ai_2
XFILLER_102_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19650__A2 _20080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20796__A1 _20799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21993__B1 _22090_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_990 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17413__A1 _16408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22915_ _22915_/A vssd1 vssd1 vccd1 vccd1 _23293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22846_ _22859_/A _22828_/Y _22845_/Y _22858_/A vssd1 vssd1 vccd1 vccd1 _22847_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19166__A1 _12052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20349__C _23554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22777_ _22630_/X _22813_/B _22828_/B vssd1 vssd1 vccd1 vccd1 _22777_/Y sky130_fd_sc_hd__o21ai_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12530_ _12540_/C vssd1 vssd1 vccd1 vccd1 _18565_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21728_ _21728_/A _21728_/B _21728_/C vssd1 vssd1 vccd1 vccd1 _21728_/Y sky130_fd_sc_hd__nand3_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ _11847_/A _11936_/A _12460_/Y vssd1 vssd1 vccd1 vccd1 _12461_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_40_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21659_ _21659_/A _21659_/B vssd1 vssd1 vccd1 vccd1 _23552_/D sky130_fd_sc_hd__xnor2_1
X_14200_ _14883_/A _14094_/X _14878_/A _14089_/Y vssd1 vssd1 vccd1 vccd1 _14202_/C
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__18677__B1 _18503_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15180_ _15249_/B vssd1 vssd1 vccd1 vccd1 _15187_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12392_ _12393_/A _12393_/B _12392_/C vssd1 vssd1 vccd1 vccd1 _12392_/X sky130_fd_sc_hd__and3_1
XFILLER_166_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ _14131_/A vssd1 vssd1 vccd1 vccd1 _14217_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23329_ _23430_/CLK _23329_/D vssd1 vssd1 vccd1 vccd1 _23329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ _14588_/A _14050_/X _14061_/X _14901_/A _14760_/B vssd1 vssd1 vccd1 vccd1
+ _14063_/B sky130_fd_sc_hd__o311a_1
XFILLER_106_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13013_ _20494_/D _20498_/A vssd1 vssd1 vccd1 vccd1 _20628_/A sky130_fd_sc_hd__nand2_2
XFILLER_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18870_ _18869_/X _18665_/Y _18666_/X _18785_/A _18880_/B vssd1 vssd1 vccd1 vccd1
+ _18870_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_133_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17821_ _17821_/A _17821_/B vssd1 vssd1 vccd1 vccd1 _17949_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17752_ _17752_/A vssd1 vssd1 vccd1 vccd1 _17752_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12477__B1 _12478_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14964_ _14964_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _23272_/D sky130_fd_sc_hd__nor2_1
XFILLER_130_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16703_ _16225_/A _16928_/A _16662_/B _16662_/A vssd1 vssd1 vccd1 vccd1 _16704_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_130_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13915_ _23352_/Q _23350_/Q _23351_/Q vssd1 vssd1 vccd1 vccd1 _13949_/A sky130_fd_sc_hd__nor3_1
X_17683_ _17703_/A vssd1 vssd1 vccd1 vccd1 _17935_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_47_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14895_ _14174_/B _14887_/A _14754_/X _14757_/Y vssd1 vssd1 vccd1 vccd1 _14896_/C
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__14819__A _14819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19422_ _19422_/A _19422_/B vssd1 vssd1 vccd1 vccd1 _19423_/C sky130_fd_sc_hd__nand2_1
XFILLER_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16634_ _18755_/C _18755_/D _16634_/C vssd1 vssd1 vccd1 vccd1 _16635_/B sky130_fd_sc_hd__and3_1
XFILLER_90_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15966__A1 _16119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13846_ _13341_/X _13474_/A _13668_/A vssd1 vssd1 vccd1 vccd1 _13846_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19353_ _19353_/A _19353_/B _19353_/C vssd1 vssd1 vccd1 vccd1 _19398_/B sky130_fd_sc_hd__nand3_2
X_16565_ _16565_/A _16565_/B _16565_/C vssd1 vssd1 vccd1 vccd1 _16567_/B sky130_fd_sc_hd__nand3_1
XFILLER_16_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13777_ _13634_/X _13630_/Y _13768_/Y _13771_/Y _13636_/X vssd1 vssd1 vccd1 vccd1
+ _13777_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_188_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12244__A3 _16523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18304_ _18296_/X _18295_/X _18267_/Y _18301_/B vssd1 vssd1 vccd1 vccd1 _18304_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_149_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15516_ _15516_/A _15517_/A _15540_/A vssd1 vssd1 vccd1 vccd1 _15516_/X sky130_fd_sc_hd__and3_1
X_19284_ _19294_/C _19294_/D _19284_/C _19293_/A vssd1 vssd1 vccd1 vccd1 _19457_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_149_929 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12728_ _12728_/A _12728_/B vssd1 vssd1 vccd1 vccd1 _12728_/Y sky130_fd_sc_hd__nand2_1
X_16496_ _12149_/X _16167_/C _15704_/A _16529_/C _16549_/C vssd1 vssd1 vccd1 vccd1
+ _16496_/X sky130_fd_sc_hd__a32o_1
XANTENNA__16915__B1 _16662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18235_ _18236_/B _18236_/C _18236_/A vssd1 vssd1 vccd1 vccd1 _18322_/A sky130_fd_sc_hd__o21a_1
XFILLER_175_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15447_ _14995_/A _14995_/B _15445_/X _15536_/A _15446_/X vssd1 vssd1 vccd1 vccd1
+ _15447_/Y sky130_fd_sc_hd__a2111oi_4
X_12659_ _20675_/B vssd1 vssd1 vccd1 vccd1 _20966_/B sky130_fd_sc_hd__buf_2
XFILLER_129_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18166_ _19967_/C vssd1 vssd1 vccd1 vccd1 _20151_/C sky130_fd_sc_hd__buf_2
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15378_ _15379_/A _15379_/B _15377_/X vssd1 vssd1 vccd1 vccd1 _15382_/A sky130_fd_sc_hd__o21bai_1
XFILLER_184_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ _17302_/A _17301_/A _17301_/B vssd1 vssd1 vccd1 vccd1 _17117_/Y sky130_fd_sc_hd__a21oi_1
X_14329_ _14329_/A _14340_/A vssd1 vssd1 vccd1 vccd1 _14353_/A sky130_fd_sc_hd__nand2_1
X_18097_ _18097_/A vssd1 vssd1 vccd1 vccd1 _18328_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17048_ _15884_/A _16147_/A _16625_/X _17252_/A vssd1 vssd1 vccd1 vccd1 _17048_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20291__A _20295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15816__C _16314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ _18999_/A _23396_/Q _18999_/C vssd1 vssd1 vccd1 vccd1 _19308_/C sky130_fd_sc_hd__nand3_4
XFILLER_140_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20961_ _20961_/A vssd1 vssd1 vccd1 vccd1 _21545_/A sky130_fd_sc_hd__buf_2
XFILLER_94_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22011__A _22064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14729__A _14729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22700_ _22700_/A _22790_/A _22700_/C _22700_/D vssd1 vssd1 vccd1 vccd1 _22701_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_38_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20892_ _20843_/B _20842_/A _20842_/B vssd1 vssd1 vccd1 vccd1 _20980_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22631_ _22631_/A _22631_/B vssd1 vssd1 vccd1 vccd1 _22631_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13432__A2 _13431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19320__A _19320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22562_ _22562_/A _22562_/B _22562_/C vssd1 vssd1 vccd1 vccd1 _22635_/A sky130_fd_sc_hd__nand3_2
XANTENNA__16367__D1 _12149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21513_ _21513_/A vssd1 vssd1 vccd1 vccd1 _21513_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22493_ _22493_/A _22493_/B _22493_/C vssd1 vssd1 vccd1 vccd1 _22500_/C sky130_fd_sc_hd__nand3_1
XFILLER_186_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21444_ _21445_/B _21561_/A _21445_/A vssd1 vssd1 vccd1 vccd1 _21448_/A sky130_fd_sc_hd__a21o_1
XANTENNA__18659__B1 _18959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23266__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_34 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12943__A1 _12571_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21375_ _21184_/C _21285_/Y _21373_/Y vssd1 vssd1 vccd1 vccd1 _21376_/B sky130_fd_sc_hd__a21oi_2
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23114_ _23182_/S vssd1 vssd1 vccd1 vccd1 _23123_/S sky130_fd_sc_hd__clkbuf_2
X_20326_ _20328_/A _20328_/C _20328_/B _20329_/B _20327_/A vssd1 vssd1 vccd1 vccd1
+ _20330_/A sky130_fd_sc_hd__o311a_1
XANTENNA__16685__A2 _16684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22758__A2 _22566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23045_ _13945_/X input18/X _23051_/S vssd1 vssd1 vccd1 vccd1 _23046_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20257_ _20256_/X _20250_/Y _20255_/A vssd1 vssd1 vccd1 vccd1 _20257_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12171__A2 _11852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20188_ _20188_/A vssd1 vssd1 vccd1 vccd1 _20189_/C sky130_fd_sc_hd__inv_2
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21744__B _21744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13120__A1 _13121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _11961_/A _23256_/B vssd1 vssd1 vccd1 vccd1 _11961_/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18552__B1_N _12536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13700_ _13578_/Y _13590_/Y _13587_/Y vssd1 vssd1 vccd1 vccd1 _13730_/A sky130_fd_sc_hd__a21bo_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11682__A1 _11851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14680_ _23370_/Q _14667_/X _14679_/X vssd1 vssd1 vccd1 vccd1 _14680_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11892_ _12032_/B _11877_/X _11881_/Y _11891_/Y vssd1 vssd1 vccd1 vccd1 _11912_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_879 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21182__D _21182_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13631_ _13495_/A _13418_/A _13312_/A _13279_/A vssd1 vssd1 vccd1 vccd1 _13632_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22829_ _22829_/A _22829_/B vssd1 vssd1 vccd1 vccd1 _22840_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13562_ _21988_/A _21988_/B _21778_/C _21778_/D _13709_/A vssd1 vssd1 vccd1 vccd1
+ _13720_/A sky130_fd_sc_hd__a32o_1
X_16350_ _16350_/A _16581_/B vssd1 vssd1 vccd1 vccd1 _16771_/C sky130_fd_sc_hd__nand2_1
X_12513_ _12513_/A vssd1 vssd1 vccd1 vccd1 _17590_/A sky130_fd_sc_hd__clkbuf_4
X_15301_ _15301_/A vssd1 vssd1 vccd1 vccd1 _15363_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16281_ _16281_/A _16281_/B _16281_/C _16281_/D vssd1 vssd1 vccd1 vccd1 _16282_/C
+ sky130_fd_sc_hd__nand4_1
X_13493_ _13553_/A _13732_/A _13482_/A _13400_/Y _13440_/Y vssd1 vssd1 vccd1 vccd1
+ _13494_/C sky130_fd_sc_hd__o221ai_1
XANTENNA__17570__B1 _16056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17388__C _19512_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16373__B2 _15972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14374__A _15195_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18020_ _18114_/A _18014_/B _18075_/A _18075_/B vssd1 vssd1 vccd1 vccd1 _18022_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__16292__C _18172_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15232_ _15225_/C _15054_/A _15231_/C _15293_/A vssd1 vssd1 vccd1 vccd1 _15275_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12444_ _12444_/A vssd1 vssd1 vccd1 vccd1 _12445_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_932 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17858__D1 _17766_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15163_ _15163_/A _15188_/A vssd1 vssd1 vccd1 vccd1 _15163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ _19082_/A _16480_/A _12379_/A _19082_/B vssd1 vssd1 vccd1 vccd1 _12375_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_165_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_954 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14114_ _14135_/A vssd1 vssd1 vccd1 vccd1 _14114_/X sky130_fd_sc_hd__buf_2
XFILLER_153_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19971_ _12509_/X _19670_/B _19807_/A vssd1 vssd1 vccd1 vccd1 _19972_/A sky130_fd_sc_hd__o21ai_1
X_15094_ _15094_/A _15094_/B _15094_/C vssd1 vssd1 vccd1 vccd1 _15099_/B sky130_fd_sc_hd__nand3_1
XFILLER_158_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18922_ _18922_/A vssd1 vssd1 vccd1 vccd1 _19108_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14045_ _14189_/A _14086_/A _14029_/C _14044_/B vssd1 vssd1 vccd1 vccd1 _14061_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_140_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18853_ _18959_/A _18959_/B vssd1 vssd1 vccd1 vccd1 _18858_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18822__B1 _19029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17804_ _17802_/Y _17803_/X _17709_/Y vssd1 vssd1 vccd1 vccd1 _17805_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__18947__C _18947_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18784_ _18784_/A _18784_/B _18784_/C vssd1 vssd1 vccd1 vccd1 _18880_/B sky130_fd_sc_hd__nand3_2
X_15996_ _16000_/A _16000_/B _16000_/C _15867_/Y vssd1 vssd1 vccd1 vccd1 _15996_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23572__D _23572_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17735_ _17435_/X _17434_/X _17567_/X _17259_/A vssd1 vssd1 vccd1 vccd1 _17736_/A
+ sky130_fd_sc_hd__o211ai_2
X_14947_ _14947_/A _14947_/B vssd1 vssd1 vccd1 vccd1 _14947_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17389__B1 _17305_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18050__A1 _17535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13453__A _13453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17666_ _17666_/A _17666_/B vssd1 vssd1 vccd1 vccd1 _17667_/B sky130_fd_sc_hd__nand2_1
X_14878_ _14878_/A _14970_/B vssd1 vssd1 vccd1 vccd1 _14879_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12870__B1 _12875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16061__B1 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19405_ _19400_/Y _19401_/Y _19403_/X _19404_/Y vssd1 vssd1 vccd1 vccd1 _19422_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_63_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16617_ _16832_/A vssd1 vssd1 vccd1 vccd1 _16617_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13829_ _21786_/A _21786_/B _13799_/X _13813_/X vssd1 vssd1 vccd1 vccd1 _13829_/Y
+ sky130_fd_sc_hd__o211ai_2
X_17597_ _17597_/A _17760_/A vssd1 vssd1 vccd1 vccd1 _17597_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__12069__A _23592_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14072__C1 _14188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_326 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19535__D1 _19700_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19336_ _18993_/Y _19173_/X _19333_/Y _19335_/Y vssd1 vssd1 vccd1 vccd1 _19341_/A
+ sky130_fd_sc_hd__o211ai_1
X_16548_ _16549_/A _16549_/D _16549_/B _16549_/C vssd1 vssd1 vccd1 vccd1 _16548_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19267_ _19265_/X _19266_/X _19297_/B _19297_/A vssd1 vssd1 vccd1 vccd1 _19275_/C
+ sky130_fd_sc_hd__o211ai_2
X_16479_ _16479_/A vssd1 vssd1 vccd1 vccd1 _16479_/X sky130_fd_sc_hd__clkbuf_4
X_18218_ _18218_/A vssd1 vssd1 vccd1 vccd1 _19425_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_164_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19198_ _19703_/A vssd1 vssd1 vccd1 vccd1 _20062_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_102_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_526 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19302__A1 _19172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18149_ _18149_/A _18149_/B _18149_/C _18149_/D vssd1 vssd1 vccd1 vccd1 _18149_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17595__A _17595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17849__D1 _17605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21160_ _21228_/A _21228_/B vssd1 vssd1 vccd1 vccd1 _21232_/A sky130_fd_sc_hd__nand2_1
X_20111_ _20111_/A _20111_/B _20111_/C _20111_/D vssd1 vssd1 vccd1 vccd1 _20112_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_172_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21091_ _21083_/A _21083_/B _21089_/Y _21090_/X vssd1 vssd1 vccd1 vccd1 _21091_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20042_ _20042_/A _20042_/B vssd1 vssd1 vccd1 vccd1 _20201_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21993_ _22096_/B _22090_/A _22090_/D _22090_/C vssd1 vssd1 vccd1 vccd1 _22086_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20944_ _20940_/X _20941_/Y _21057_/B _21057_/A vssd1 vssd1 vccd1 vccd1 _20945_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_57_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20875_ _21017_/B _21017_/C _21542_/A _21017_/A vssd1 vssd1 vccd1 vccd1 _20878_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16674__A _16674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14602__A1 _13603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14602__B2 _12875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22614_ _22730_/B _22540_/B _22537_/X vssd1 vssd1 vccd1 vccd1 _22615_/A sky130_fd_sc_hd__a21boi_1
XFILLER_198_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23594_ _23598_/CLK _23594_/D vssd1 vssd1 vccd1 vccd1 _23594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19541__A1 _19547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13810__B _13810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22545_ _22670_/A _22545_/B _22545_/C _22663_/D vssd1 vssd1 vccd1 vccd1 _22677_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_50_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11611__A _11611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14905__A2 _15366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22476_ _22476_/A _22476_/B _22476_/C vssd1 vssd1 vccd1 vccd1 _22476_/X sky130_fd_sc_hd__and3_1
XFILLER_148_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12426__B _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21427_ _21425_/Y _21426_/X _21407_/A _21407_/B vssd1 vssd1 vccd1 vccd1 _21473_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19844__A2 _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16840__C _18755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _12015_/Y _12027_/Y _12046_/A _12046_/B vssd1 vssd1 vccd1 vccd1 _12160_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_136_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21358_ _21358_/A _21358_/B _21358_/C vssd1 vssd1 vccd1 vccd1 _21359_/B sky130_fd_sc_hd__nand3_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20309_ _20354_/B _20257_/Y _20311_/A _20308_/Y vssd1 vssd1 vccd1 vccd1 _20310_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_151_968 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12091_ _12227_/A _12059_/A _12088_/X _19082_/A vssd1 vssd1 vccd1 vccd1 _12231_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_21289_ _21380_/A _21380_/B vssd1 vssd1 vccd1 vccd1 _21317_/A sky130_fd_sc_hd__nand2_2
XFILLER_122_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17607__A1 _17243_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23028_ _23344_/Q input25/X _23034_/S vssd1 vssd1 vccd1 vccd1 _23029_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17607__B2 _17243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15079__D1 _14069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17083__A2 _16311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15850_ _18675_/A _16370_/A _15858_/A vssd1 vssd1 vccd1 vccd1 _15943_/B sky130_fd_sc_hd__o21ai_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input20_A wb_dat_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ _14934_/A _14934_/B _14934_/C _14934_/D vssd1 vssd1 vccd1 vccd1 _14805_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_188_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16830__A2 _12223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _16027_/A _16027_/B _17066_/C _17062_/B vssd1 vssd1 vccd1 vccd1 _15781_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _20584_/A _20585_/B _13133_/C _20775_/D vssd1 vssd1 vccd1 vccd1 _13085_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _17353_/Y _17357_/Y _17515_/X _17523_/B vssd1 vssd1 vccd1 vccd1 _17537_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _18435_/B _16795_/B _14725_/Y _23582_/D vssd1 vssd1 vccd1 vccd1 _23260_/A
+ sky130_fd_sc_hd__a31o_2
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11944_ _12071_/A vssd1 vssd1 vccd1 vccd1 _16140_/A sky130_fd_sc_hd__buf_2
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _17440_/A _17450_/Y _16479_/A _17733_/A vssd1 vssd1 vccd1 vccd1 _17453_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11875_ _11875_/A vssd1 vssd1 vccd1 vccd1 _18675_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__16594__A1 _16382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14663_ _23398_/Q _14640_/X _14647_/X _23430_/Q _14662_/X vssd1 vssd1 vccd1 vccd1
+ _14663_/X sky130_fd_sc_hd__a221o_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21921__C _21921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _16402_/A _16402_/B vssd1 vssd1 vccd1 vccd1 _16403_/C sky130_fd_sc_hd__nand2_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13614_ _22126_/A _13407_/Y _13434_/B _13433_/A vssd1 vssd1 vccd1 vccd1 _13619_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17382_ _17382_/A _17382_/B _17533_/A _17382_/D vssd1 vssd1 vccd1 vccd1 _17384_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__13947__A3 _13945_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14594_ input51/X _14518_/X _14593_/X vssd1 vssd1 vccd1 vccd1 _14594_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19121_ _19121_/A vssd1 vssd1 vccd1 vccd1 _19121_/X sky130_fd_sc_hd__clkbuf_2
X_16333_ _16421_/A vssd1 vssd1 vccd1 vccd1 _16475_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_197_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13545_ _13545_/A vssd1 vssd1 vccd1 vccd1 _13545_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_854 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23581__CLK _23582_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19052_ _19052_/A _19052_/B vssd1 vssd1 vccd1 vccd1 _19055_/A sky130_fd_sc_hd__nand2_1
XANTENNA__22419__A1 _22754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13476_ _13476_/A _13476_/B _13476_/C vssd1 vssd1 vccd1 vccd1 _13477_/A sky130_fd_sc_hd__nand3_1
XANTENNA__16897__A2 _16055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16264_ _16347_/B _16347_/C vssd1 vssd1 vccd1 vccd1 _16265_/B sky130_fd_sc_hd__nand2_1
XFILLER_185_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18003_ _18003_/A vssd1 vssd1 vccd1 vccd1 _18211_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_145_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12907__B2 _12906_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15215_ _15213_/Y _15286_/B vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__and2b_1
X_12427_ _18448_/A vssd1 vssd1 vccd1 vccd1 _12427_/X sky130_fd_sc_hd__clkbuf_2
X_16195_ _16195_/A _16667_/D vssd1 vssd1 vccd1 vccd1 _16661_/A sky130_fd_sc_hd__nand2_2
XFILLER_127_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14832__A _23505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14109__B1 _14015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ _12508_/A _16549_/B _16549_/D _18778_/C vssd1 vssd1 vccd1 vccd1 _12358_/X
+ sky130_fd_sc_hd__and4_1
X_15146_ _15063_/A _15066_/Y _15286_/A _15144_/X vssd1 vssd1 vccd1 vccd1 _15146_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_127_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15857__B1 _15855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19954_ _19951_/B _19951_/C _20081_/B _20366_/C vssd1 vssd1 vccd1 vccd1 _20043_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_15077_ _15077_/A _15077_/B _15077_/C vssd1 vssd1 vccd1 vccd1 _15077_/X sky130_fd_sc_hd__and3_1
X_12289_ _12289_/A _12289_/B vssd1 vssd1 vccd1 vccd1 _12547_/B sky130_fd_sc_hd__nor2_2
XFILLER_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18905_ _18897_/C _18897_/D _18904_/Y vssd1 vssd1 vccd1 vccd1 _18905_/X sky130_fd_sc_hd__a21o_1
X_14028_ _14193_/A vssd1 vssd1 vccd1 vccd1 _14029_/C sky130_fd_sc_hd__clkbuf_2
X_19885_ _19883_/Y _19884_/X _19877_/Y vssd1 vssd1 vccd1 vccd1 _19889_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__17862__B _17959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16806__C1 _15964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18836_ _18836_/A _18836_/B vssd1 vssd1 vccd1 vccd1 _19703_/D sky130_fd_sc_hd__nand2_2
XFILLER_110_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18767_ _18767_/A _18767_/B _18767_/C vssd1 vssd1 vccd1 vccd1 _18966_/A sky130_fd_sc_hd__nand3_4
X_15979_ _15982_/A _15979_/B vssd1 vssd1 vccd1 vccd1 _15979_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17718_ _17597_/Y _17711_/Y _17715_/Y _17717_/Y vssd1 vssd1 vccd1 vccd1 _17838_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19220__B1 _19013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18698_ _18696_/Y _18697_/X _18667_/Y _18672_/Y vssd1 vssd1 vccd1 vccd1 _18751_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16034__B1 _15749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17649_ _17792_/A _17788_/A _17649_/C vssd1 vssd1 vccd1 vccd1 _17657_/C sky130_fd_sc_hd__nand3_2
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20660_ _20660_/A vssd1 vssd1 vccd1 vccd1 _21046_/A sky130_fd_sc_hd__buf_2
XFILLER_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19319_ _19172_/A _19172_/B _19172_/C _19183_/C vssd1 vssd1 vccd1 vccd1 _19325_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__21866__C1 _21864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20591_ _20578_/X _20736_/B _20576_/Y _20568_/Y vssd1 vssd1 vccd1 vccd1 _21008_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22330_ _22201_/Y _22205_/Y _22207_/B vssd1 vssd1 vccd1 vccd1 _22330_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_191_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__D _18755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22261_ _22139_/B _22139_/C _22139_/A vssd1 vssd1 vccd1 vccd1 _22261_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__15560__A2 _15552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21212_ _21212_/A _21212_/B _21212_/C _21212_/D vssd1 vssd1 vccd1 vccd1 _21218_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_145_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22192_ _22700_/A _22554_/A _22192_/C _22192_/D vssd1 vssd1 vccd1 vccd1 _22192_/Y
+ sky130_fd_sc_hd__nand4_4
X_21143_ _21345_/A _21141_/X _21142_/Y vssd1 vssd1 vccd1 vccd1 _21144_/B sky130_fd_sc_hd__o21a_1
XANTENNA__19039__B1 _18840_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12262__A _12475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18868__B _18868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21074_ _21071_/Y _21073_/Y _20905_/Y vssd1 vssd1 vccd1 vccd1 _21078_/A sky130_fd_sc_hd__o21ai_1
XFILLER_86_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20025_ _20113_/B _20025_/B vssd1 vssd1 vccd1 vccd1 _20207_/D sky130_fd_sc_hd__nand2_1
XFILLER_59_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11885__B2 _11784_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16273__B1 _16275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13093__A _23456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19211__B1 _19013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ _21976_/A _23272_/Q _21976_/C vssd1 vssd1 vccd1 vccd1 _21977_/B sky130_fd_sc_hd__nand3_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_771 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20927_ _20783_/Y _20790_/B _20778_/X _20934_/A vssd1 vssd1 vccd1 vccd1 _20941_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20638__B _23297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _11980_/A _11823_/B _11983_/A vssd1 vssd1 vccd1 vccd1 _11684_/A sky130_fd_sc_hd__nand3_1
XFILLER_70_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20858_ _20589_/A _20589_/C _20722_/A _20853_/B vssd1 vssd1 vccd1 vccd1 _20858_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23577_ _23578_/CLK _23577_/D vssd1 vssd1 vccd1 vccd1 _23577_/Q sky130_fd_sc_hd__dfxtp_1
X_11591_ _11808_/A vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__buf_2
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20789_ _20789_/A _20789_/B _20789_/C vssd1 vssd1 vccd1 vccd1 _20819_/A sky130_fd_sc_hd__nand3_2
XFILLER_183_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13330_ _13701_/C vssd1 vssd1 vccd1 vccd1 _21987_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22528_ _22528_/A _22528_/B vssd1 vssd1 vccd1 vccd1 _22629_/B sky130_fd_sc_hd__nand2_1
XFILLER_168_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ _23333_/Q vssd1 vssd1 vccd1 vccd1 _21739_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22459_ _22414_/X _22415_/Y _22400_/B _22400_/A vssd1 vssd1 vccd1 vccd1 _22541_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__19817__A2 _17763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15551__A2 _15528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16997__A_N _23523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12212_ _12199_/A _12199_/B _12210_/Y _12211_/X vssd1 vssd1 vccd1 vccd1 _12531_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_15000_ _15000_/A _15000_/B vssd1 vssd1 vccd1 vccd1 _15000_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13562__A1 _21988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13192_ _13191_/A _13191_/B _13191_/C _13191_/D vssd1 vssd1 vccd1 vccd1 _13192_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12143_ _12107_/X _12110_/Y _12104_/X vssd1 vssd1 vccd1 vccd1 _12143_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__13268__A _13766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12172__A _16122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18778__B _18778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ _12222_/A _12223_/A vssd1 vssd1 vccd1 vccd1 _15860_/D sky130_fd_sc_hd__nand2_1
X_16951_ _16951_/A vssd1 vssd1 vccd1 vccd1 _17184_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20045__D1 _20320_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18789__C1 _18479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15902_ _15908_/B _15902_/B vssd1 vssd1 vccd1 vccd1 _15902_/Y sky130_fd_sc_hd__nand2_1
X_19670_ _19670_/A _19670_/B _19670_/C vssd1 vssd1 vccd1 vccd1 _19670_/X sky130_fd_sc_hd__or3_1
X_16882_ _16890_/B _16893_/C vssd1 vssd1 vccd1 vccd1 _16882_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18621_ _18615_/A _18615_/B _18615_/C _18617_/X vssd1 vssd1 vccd1 vccd1 _18931_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_37_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _16160_/A vssd1 vssd1 vccd1 vccd1 _17057_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22077__B1_N _22218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_72 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _12537_/B _12528_/A _12536_/B vssd1 vssd1 vccd1 vccd1 _18555_/B sky130_fd_sc_hd__a21bo_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _15761_/X _15762_/Y _15763_/Y vssd1 vssd1 vccd1 vccd1 _15883_/A sky130_fd_sc_hd__o21ai_2
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _12975_/A _12975_/B _12975_/C vssd1 vssd1 vccd1 vccd1 _12977_/C sky130_fd_sc_hd__a21o_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _17345_/A _17350_/D _17350_/C vssd1 vssd1 vccd1 vccd1 _17513_/C sky130_fd_sc_hd__a21bo_1
XFILLER_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _23348_/Q _14531_/A _14546_/A _23316_/Q _14657_/A vssd1 vssd1 vccd1 vccd1
+ _14715_/X sky130_fd_sc_hd__a221o_1
XFILLER_75_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _16593_/A vssd1 vssd1 vccd1 vccd1 _18859_/A sky130_fd_sc_hd__buf_2
XFILLER_75_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18483_ _18483_/A vssd1 vssd1 vccd1 vccd1 _18484_/A sky130_fd_sc_hd__buf_2
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15695_ _15648_/A _15693_/Y _15694_/Y vssd1 vssd1 vccd1 vccd1 _15983_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__17764__B1 _17465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _17434_/A vssd1 vssd1 vccd1 vccd1 _17434_/X sky130_fd_sc_hd__buf_2
XANTENNA__18508__A2_N _18504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14646_ _14646_/A vssd1 vssd1 vccd1 vccd1 _18434_/A sky130_fd_sc_hd__buf_4
X_11858_ _11912_/A _11912_/B vssd1 vssd1 vccd1 vccd1 _11903_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13450__B _21921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_487 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17365_ _17365_/A _17365_/B _17365_/C _17365_/D vssd1 vssd1 vccd1 vccd1 _17522_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA__12347__A _17546_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14577_ _23267_/Q _14551_/X _14547_/A _12608_/X vssd1 vssd1 vccd1 vccd1 _14577_/X
+ sky130_fd_sc_hd__a22o_1
X_11789_ _11789_/A _11789_/B vssd1 vssd1 vccd1 vccd1 _11847_/A sky130_fd_sc_hd__nand2_2
X_19104_ _19104_/A _19289_/B _19104_/C vssd1 vssd1 vccd1 vccd1 _19105_/B sky130_fd_sc_hd__and3_1
XFILLER_159_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ _18461_/A _16451_/B _16451_/C _15972_/X _16194_/A vssd1 vssd1 vccd1 vccd1
+ _16316_/Y sky130_fd_sc_hd__o32ai_4
XFILLER_186_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13528_ _13814_/B vssd1 vssd1 vccd1 vccd1 _21919_/C sky130_fd_sc_hd__buf_2
X_17296_ _17477_/A _17477_/B _17297_/C _17297_/D vssd1 vssd1 vccd1 vccd1 _17299_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_846 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19035_ _19138_/A _19139_/A _19035_/C vssd1 vssd1 vccd1 vccd1 _19036_/B sky130_fd_sc_hd__nand3_1
XFILLER_118_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23065__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16247_ _16254_/A _16254_/B _16247_/C _16247_/D vssd1 vssd1 vccd1 vccd1 _16248_/D
+ sky130_fd_sc_hd__nand4_2
X_13459_ _13517_/A _13513_/A _13463_/A vssd1 vssd1 vccd1 vccd1 _13461_/B sky130_fd_sc_hd__a21bo_1
XFILLER_63_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19808__A2 _18003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12356__A2 _11747_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16178_ _16175_/B _16175_/C _16175_/A vssd1 vssd1 vccd1 vccd1 _16179_/C sky130_fd_sc_hd__a21o_1
XFILLER_115_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18492__A1 _12323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15129_ _15129_/A _15129_/B vssd1 vssd1 vccd1 vccd1 _15132_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15096__C _15238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12108__A2 _12093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13305__A1 _23322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19937_ _19889_/B _19889_/C _19889_/A vssd1 vssd1 vccd1 vccd1 _19937_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_130_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19868_ _19868_/A vssd1 vssd1 vccd1 vccd1 _20142_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__21545__D _21635_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17452__C1 _20062_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18819_ _12004_/X _12006_/X _19505_/A _19504_/A _19157_/A vssd1 vssd1 vccd1 vccd1
+ _18835_/A sky130_fd_sc_hd__o221ai_4
XANTENNA__13069__B1 _13061_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19799_ _19966_/A _20062_/C _19799_/C _19967_/A vssd1 vssd1 vccd1 vccd1 _20013_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21830_ _23481_/Q vssd1 vssd1 vccd1 vccd1 _22510_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22879__A1 _22878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21761_ _21766_/A _21767_/A _21919_/C vssd1 vssd1 vccd1 vccd1 _21922_/A sky130_fd_sc_hd__nand3_2
XANTENNA__12292__B2 _12374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20712_ _20712_/A _20718_/B vssd1 vssd1 vccd1 vccd1 _20716_/A sky130_fd_sc_hd__nand2_1
X_23500_ _23510_/CLK _23500_/D vssd1 vssd1 vccd1 vccd1 _23500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21692_ _21688_/A _21688_/B _21688_/D _21691_/X vssd1 vssd1 vccd1 vccd1 _21717_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_196_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14033__A2 _14029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15230__A1 _14834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23431_ _23431_/CLK _23431_/D vssd1 vssd1 vccd1 vccd1 _23431_/Q sky130_fd_sc_hd__dfxtp_1
X_20643_ _20479_/X _20639_/Y _12601_/C _20894_/B vssd1 vssd1 vccd1 vccd1 _20917_/A
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12257__A _17133_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19966__C _20133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23362_ _23363_/CLK _23362_/D vssd1 vssd1 vccd1 vccd1 _23362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20574_ _20579_/B vssd1 vssd1 vccd1 vccd1 _20589_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22313_ _22310_/Y _22199_/A _22288_/Y _22289_/Y vssd1 vssd1 vccd1 vccd1 _22313_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__22392__C _22392_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23056__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20905__C _20905_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23293_ _23296_/CLK _23293_/D vssd1 vssd1 vccd1 vccd1 _23293_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_194_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14472__A _14933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22244_ _22439_/D _22439_/C _22439_/B vssd1 vssd1 vccd1 vccd1 _22246_/A sky130_fd_sc_hd__nand3_1
XFILLER_106_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17286__A2 _17285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22175_ _22167_/X _22170_/Y _22174_/Y vssd1 vssd1 vccd1 vccd1 _22176_/A sky130_fd_sc_hd__o21ai_2
XFILLER_79_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21126_ _21134_/A _21134_/B vssd1 vssd1 vccd1 vccd1 _21126_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13816__A _13816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21057_ _21057_/A _21057_/B vssd1 vssd1 vccd1 vccd1 _21057_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20008_ _19937_/Y _19938_/Y _20004_/Y _20007_/Y vssd1 vssd1 vccd1 vccd1 _20111_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_189_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18786__A2 _18868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16549__D _16549_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _20532_/A vssd1 vssd1 vccd1 vccd1 _13115_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_185_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12864_/A _12864_/B _12760_/Y vssd1 vssd1 vccd1 vccd1 _12770_/C sky130_fd_sc_hd__a21o_4
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20433__B1_N _20431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ _21820_/A _21817_/Y _21819_/B vssd1 vssd1 vccd1 vccd1 _21964_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__20368__B _20368_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14846_/A _14846_/B _14847_/A _14847_/B vssd1 vssd1 vccd1 vccd1 _14501_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _12036_/A _11721_/A _11708_/Y vssd1 vssd1 vccd1 vccd1 _11713_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15480_ _15476_/B _15476_/A _15475_/A vssd1 vssd1 vccd1 vccd1 _15503_/A sky130_fd_sc_hd__o21ai_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12577_/A _20639_/A _12580_/A _20639_/D _12683_/Y vssd1 vssd1 vccd1 vccd1
+ _12692_/Y sky130_fd_sc_hd__a41oi_4
XFILLER_43_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _23585_/Q vssd1 vssd1 vccd1 vccd1 _11739_/B sky130_fd_sc_hd__buf_2
X_14431_ _14427_/Y _14428_/X _14456_/B vssd1 vssd1 vccd1 vccd1 _14436_/B sky130_fd_sc_hd__o21ai_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12167__A _12167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17150_ _17150_/A _17150_/B vssd1 vssd1 vccd1 vccd1 _17151_/C sky130_fd_sc_hd__nand2_1
X_11574_ _23598_/Q vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14362_ _14358_/C _14358_/B _14359_/X _14361_/X vssd1 vssd1 vccd1 vccd1 _14362_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_10_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 wb_dat_i[19] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 wb_dat_i[29] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_2
X_16101_ _16093_/Y _16096_/Y _16091_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 _16425_/B
+ sky130_fd_sc_hd__o22ai_1
Xinput39 wb_stb_i vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_2
X_13313_ _13466_/A vssd1 vssd1 vccd1 vccd1 _13313_/X sky130_fd_sc_hd__buf_2
XFILLER_183_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17081_ _16823_/Y _16825_/Y _17073_/Y _16843_/Y vssd1 vssd1 vccd1 vccd1 _17126_/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA__23047__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14293_ _14367_/A _14367_/B _14367_/C vssd1 vssd1 vccd1 vccd1 _14294_/B sky130_fd_sc_hd__a21boi_1
XFILLER_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13244_ _13520_/A _13732_/B _13732_/C _13243_/Y vssd1 vssd1 vccd1 vccd1 _13247_/A
+ sky130_fd_sc_hd__o31ai_1
X_16032_ _16032_/A vssd1 vssd1 vccd1 vccd1 _16032_/X sky130_fd_sc_hd__buf_4
XFILLER_170_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19266__A3 _18928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18420__A_N _23537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13175_ _13148_/X _13149_/Y _13171_/Y _13174_/Y vssd1 vssd1 vccd1 vccd1 _13175_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_124_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12126_ _12426_/B _12426_/C vssd1 vssd1 vccd1 vccd1 _18444_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17983_ _17988_/A _17988_/D vssd1 vssd1 vccd1 vccd1 _17992_/A sky130_fd_sc_hd__nand2_1
XFILLER_151_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_990 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19722_ _19722_/A _19722_/B _19722_/C vssd1 vssd1 vccd1 vccd1 _19725_/A sky130_fd_sc_hd__nand3_1
X_12057_ _12057_/A _12057_/B _12057_/C vssd1 vssd1 vccd1 vccd1 _12204_/B sky130_fd_sc_hd__nand3_1
X_16934_ _16934_/A _16934_/B _16934_/C vssd1 vssd1 vccd1 vccd1 _16934_/X sky130_fd_sc_hd__and3_2
XFILLER_77_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19116__C _19116_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20033__A1 _20031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19653_ _19653_/A _19862_/B _19862_/C vssd1 vssd1 vccd1 vccd1 _19653_/X sky130_fd_sc_hd__and3_1
XFILLER_120_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16865_ _16865_/A vssd1 vssd1 vccd1 vccd1 _17605_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16788__A1 _16988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18604_ _18604_/A vssd1 vssd1 vccd1 vccd1 _18604_/X sky130_fd_sc_hd__buf_2
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15941__A _15941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15816_ _19165_/C _16314_/B _16314_/C vssd1 vssd1 vccd1 vccd1 _16029_/B sky130_fd_sc_hd__and3_1
X_19584_ _19475_/X _19527_/Y _19571_/Y _19574_/X _19583_/Y vssd1 vssd1 vccd1 vccd1
+ _19592_/B sky130_fd_sc_hd__o221ai_1
X_16796_ _16796_/A _23597_/Q vssd1 vssd1 vccd1 vccd1 _16796_/X sky130_fd_sc_hd__and2_2
XFILLER_93_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18535_ _12508_/D _17586_/A _17587_/A _18532_/Y _18534_/Y vssd1 vssd1 vccd1 vccd1
+ _18540_/A sky130_fd_sc_hd__a32o_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _15735_/C _15662_/B _15665_/B _15677_/Y vssd1 vssd1 vccd1 vccd1 _15749_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _21276_/A _13181_/B _12958_/Y _12949_/Y vssd1 vssd1 vccd1 vccd1 _12959_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18934__C1 _17595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18466_ _11758_/A _18810_/A _18997_/B vssd1 vssd1 vccd1 vccd1 _18475_/A sky130_fd_sc_hd__a21o_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15678_ _23418_/Q _15735_/B vssd1 vssd1 vccd1 vccd1 _15678_/Y sky130_fd_sc_hd__nand2_2
XFILLER_178_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17417_ _17557_/B _17417_/B _17557_/A vssd1 vssd1 vccd1 vccd1 _17429_/A sky130_fd_sc_hd__nand3_1
XFILLER_178_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14629_ _16191_/A _14575_/X _14626_/X _14628_/X vssd1 vssd1 vccd1 vccd1 _14629_/X
+ sky130_fd_sc_hd__a22o_1
X_18397_ _18400_/A _18414_/C _18400_/C vssd1 vssd1 vccd1 vccd1 _18398_/C sky130_fd_sc_hd__nand3_1
XANTENNA__12077__A _19811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12508__C _19811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17348_ _17220_/X _17179_/X _17346_/A vssd1 vssd1 vccd1 vccd1 _17351_/A sky130_fd_sc_hd__o21ai_1
XFILLER_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18162__B1 _20215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23038__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15388__A _15538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17279_ _17258_/Y _17268_/Y _17276_/Y _17278_/Y vssd1 vssd1 vccd1 vccd1 _17297_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19018_ _19018_/A vssd1 vssd1 vccd1 vccd1 _19018_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12329__A2 _18755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13526__B2 _21891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20290_ _20237_/Y _20290_/B vssd1 vssd1 vccd1 vccd1 _20295_/A sky130_fd_sc_hd__nand2b_1
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22261__A2 _22139_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18849__D _19017_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17753__D _20055_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22014__A _22014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18211__B _18211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17108__A _19662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22013__A2 _22484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19965__A1 _19218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18768__A2 _17443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21853__A _21853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19965__B2 _17565_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22931_ _22953_/A vssd1 vssd1 vccd1 vccd1 _22940_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__16779__A1 _16275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15851__A _15941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19323__A _19323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22862_ _22830_/X _22860_/X _22861_/X vssd1 vssd1 vccd1 vccd1 _22862_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23490__D _23502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21813_ _21811_/X _21812_/Y _21803_/Y _21806_/X vssd1 vssd1 vccd1 vccd1 _21813_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22793_ _22560_/A _22560_/B _22237_/X _22791_/X _22792_/X vssd1 vssd1 vccd1 vccd1
+ _22797_/C sky130_fd_sc_hd__a2111oi_4
XFILLER_97_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21744_ _21744_/A _21744_/B _21744_/C vssd1 vssd1 vccd1 vccd1 _22057_/A sky130_fd_sc_hd__nor3_2
XFILLER_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15739__C1 _16122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20619__D _21036_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21675_ _21666_/A _21630_/B _21649_/C vssd1 vssd1 vccd1 vccd1 _21675_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20626_ _20475_/A _20475_/B _20485_/Y vssd1 vssd1 vccd1 vccd1 _20626_/Y sky130_fd_sc_hd__a21oi_1
X_23414_ _23416_/CLK _23414_/D vssd1 vssd1 vccd1 vccd1 _23414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11776__B1 _11741_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23345_ _23345_/CLK _23345_/D vssd1 vssd1 vccd1 vccd1 _23345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20557_ _20557_/A _20557_/B vssd1 vssd1 vccd1 vccd1 _20557_/Y sky130_fd_sc_hd__nand2_1
XFILLER_153_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_451 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23276_ _23559_/CLK _23276_/D vssd1 vssd1 vccd1 vccd1 _23276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20488_ _13029_/A _13029_/B _13001_/X vssd1 vssd1 vccd1 vccd1 _20488_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22227_ _22225_/A _22231_/B _22223_/X _22226_/X vssd1 vssd1 vccd1 vccd1 _22227_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_65_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18402__A _23535_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22158_ _22158_/A vssd1 vssd1 vccd1 vccd1 _22290_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_65_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21109_ _21109_/A vssd1 vssd1 vccd1 vccd1 _21228_/A sky130_fd_sc_hd__clkbuf_2
X_14980_ _14980_/A vssd1 vssd1 vccd1 vccd1 _15010_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22089_ _22089_/A _22089_/B vssd1 vssd1 vccd1 vccd1 _22094_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13931_ _23495_/Q vssd1 vssd1 vccd1 vccd1 _14374_/D sky130_fd_sc_hd__buf_2
XANTENNA__17960__B _17960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_524 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16650_ _16650_/A _16650_/B vssd1 vssd1 vccd1 vccd1 _16650_/Y sky130_fd_sc_hd__nor2_1
X_13862_ _22713_/C vssd1 vssd1 vccd1 vccd1 _22800_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15601_ _23423_/Q vssd1 vssd1 vccd1 vccd1 _15634_/A sky130_fd_sc_hd__inv_2
X_12813_ _12810_/A _12810_/B _12812_/Y vssd1 vssd1 vccd1 vccd1 _12816_/C sky130_fd_sc_hd__a21oi_1
XFILLER_74_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16581_ _16581_/A _16581_/B _16581_/C vssd1 vssd1 vccd1 vccd1 _16582_/B sky130_fd_sc_hd__nand3_1
X_13793_ _13793_/A _13793_/B vssd1 vssd1 vccd1 vccd1 _13793_/Y sky130_fd_sc_hd__nand2_2
XFILLER_62_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18320_ _18304_/Y _18306_/Y _18307_/Y vssd1 vssd1 vccd1 vccd1 _18320_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13281__A _13766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15532_ _15516_/A _15517_/Y _15518_/X vssd1 vssd1 vccd1 vccd1 _15545_/B sky130_fd_sc_hd__o21a_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12744_ _12874_/B _12756_/A vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__nand2_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18251_ _18251_/A _18251_/B vssd1 vssd1 vccd1 vccd1 _18302_/B sky130_fd_sc_hd__nand2_1
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12008__A1 _11822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17688__A _23527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15463_ _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15463_/Y sky130_fd_sc_hd__nand2_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15745__A2 _16447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _23293_/Q vssd1 vssd1 vccd1 vccd1 _12675_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_187_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17202_ _17202_/A _17202_/B vssd1 vssd1 vccd1 vccd1 _17202_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ _14414_/A _14414_/B _14416_/B vssd1 vssd1 vccd1 vccd1 _14415_/C sky130_fd_sc_hd__nand3_1
X_18182_ _18182_/A _18182_/B vssd1 vssd1 vccd1 vccd1 _18185_/B sky130_fd_sc_hd__and2_1
XFILLER_175_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11626_ _11634_/B vssd1 vssd1 vccd1 vccd1 _16619_/A sky130_fd_sc_hd__buf_4
X_15394_ _15214_/A _15214_/B _15392_/Y _15393_/Y _15286_/Y vssd1 vssd1 vccd1 vccd1
+ _15395_/C sky130_fd_sc_hd__o221ai_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17133_ _17133_/A _17133_/B _17133_/C vssd1 vssd1 vccd1 vccd1 _17134_/A sky130_fd_sc_hd__and3_1
XFILLER_184_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18695__A1 _18673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14345_ _14356_/A _14356_/B _14356_/C _14403_/C _14403_/D vssd1 vssd1 vccd1 vccd1
+ _14350_/B sky130_fd_sc_hd__a32o_1
XFILLER_183_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22491__A2 _22558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12625__A _23449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13508__A1 _13732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17064_ _17064_/A _17260_/A vssd1 vssd1 vccd1 vccd1 _17070_/A sky130_fd_sc_hd__nand2_1
XFILLER_170_101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14276_ _14276_/A vssd1 vssd1 vccd1 vccd1 _14457_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16015_ _15725_/Y _15898_/X _15944_/Y vssd1 vssd1 vccd1 vccd1 _16015_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_143_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13227_ _21745_/A vssd1 vssd1 vccd1 vccd1 _13394_/B sky130_fd_sc_hd__buf_2
XANTENNA__23575__D _23575_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13158_ _13158_/A _21182_/D vssd1 vssd1 vccd1 vccd1 _13158_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _18445_/A vssd1 vssd1 vccd1 vccd1 _19010_/A sky130_fd_sc_hd__buf_2
X_17966_ _17966_/A _17966_/B vssd1 vssd1 vccd1 vccd1 _17967_/A sky130_fd_sc_hd__nand2_1
X_13089_ _13072_/Y _13089_/B _13089_/C vssd1 vssd1 vccd1 vccd1 _20595_/A sky130_fd_sc_hd__nand3b_1
XFILLER_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17407__C1 _17233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19947__A1 _19156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21203__B1 _12862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19705_ _19705_/A _19819_/A _19820_/A _19966_/A vssd1 vssd1 vccd1 vccd1 _19831_/B
+ sky130_fd_sc_hd__nand4_1
X_16917_ _16923_/B vssd1 vssd1 vccd1 vccd1 _16917_/X sky130_fd_sc_hd__buf_2
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17897_ _17899_/A _17886_/X _18030_/A _17896_/Y vssd1 vssd1 vccd1 vccd1 _17901_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_120_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19636_ _19636_/A _19636_/B vssd1 vssd1 vccd1 vccd1 _19636_/Y sky130_fd_sc_hd__nor2_1
X_16848_ _17057_/A _18607_/C _18607_/A _19703_/B _16027_/D vssd1 vssd1 vccd1 vccd1
+ _16848_/Y sky130_fd_sc_hd__a32oi_2
XFILLER_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19567_ _19567_/A _19567_/B _19567_/C vssd1 vssd1 vccd1 vccd1 _19588_/B sky130_fd_sc_hd__nand3_2
X_16779_ _16275_/X _16278_/Y _16989_/B _16989_/A vssd1 vssd1 vccd1 vccd1 _16998_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_92_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15984__A2 _16123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19175__A2 _19173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18518_ _18518_/A _18518_/B _18520_/B vssd1 vssd1 vccd1 vccd1 _18518_/X sky130_fd_sc_hd__and3_1
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19498_ _19522_/A _19521_/B _19577_/C vssd1 vssd1 vccd1 vccd1 _19575_/B sky130_fd_sc_hd__nand3_2
XFILLER_22_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18449_ _18452_/A _18453_/A _18456_/A vssd1 vssd1 vccd1 vccd1 _18462_/A sky130_fd_sc_hd__o21ai_1
X_21460_ _21513_/A _21460_/B _21460_/C vssd1 vssd1 vccd1 vccd1 _21463_/D sky130_fd_sc_hd__nand3b_1
XFILLER_147_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22009__A _22218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20411_ _20411_/A _20411_/B _20411_/C vssd1 vssd1 vccd1 vccd1 _20412_/B sky130_fd_sc_hd__nand3_1
XANTENNA__18686__A1 _12214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21391_ _21391_/A _21465_/A _21391_/C vssd1 vssd1 vccd1 vccd1 _21465_/B sky130_fd_sc_hd__nand3_2
XFILLER_105_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23130_ _12113_/X input36/X _23134_/S vssd1 vssd1 vccd1 vccd1 _23131_/A sky130_fd_sc_hd__mux2_1
X_20342_ _20337_/Y _20384_/B _20340_/Y _20341_/X vssd1 vssd1 vccd1 vccd1 _20342_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_146_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21848__A _21852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12707__C1 _13184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23061_ _23061_/A vssd1 vssd1 vccd1 vccd1 _23358_/D sky130_fd_sc_hd__clkbuf_1
X_20273_ _20271_/C _20271_/Y _20269_/X _20270_/X vssd1 vssd1 vccd1 vccd1 _20400_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_1_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20471__B _21493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22012_ _22564_/A _22564_/B _22172_/C vssd1 vssd1 vccd1 vccd1 _22012_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__23485__D _23497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21993__A1 _22096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11930__B1 _11677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23195__A0 _14569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16677__A _16677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17413__A2 _16741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22914_ _12675_/X input36/X _22918_/S vssd1 vssd1 vccd1 vccd1 _22915_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20953__C1 _21358_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22845_ _22849_/A _22849_/B vssd1 vssd1 vccd1 vccd1 _22845_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_71_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19166__A2 _19838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22170__A1 _13642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22776_ _22810_/B _22774_/X _22775_/Y vssd1 vssd1 vccd1 vccd1 _22828_/B sky130_fd_sc_hd__o21a_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11997__B1 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21727_ _21717_/A _21717_/B _21723_/Y vssd1 vssd1 vccd1 vccd1 _21728_/A sky130_fd_sc_hd__o21bai_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21658_ _21624_/B _21656_/X _21657_/X vssd1 vssd1 vccd1 vccd1 _21659_/B sky130_fd_sc_hd__o21ai_1
X_12460_ _12184_/A _12185_/A _12474_/A vssd1 vssd1 vccd1 vccd1 _12460_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_149_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_120 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20609_ _20608_/B _20608_/C _20608_/A vssd1 vssd1 vccd1 vccd1 _20765_/A sky130_fd_sc_hd__a21oi_1
X_12391_ _12391_/A _12391_/B _12391_/C vssd1 vssd1 vccd1 vccd1 _12396_/B sky130_fd_sc_hd__nand3_2
XFILLER_71_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21589_ _21524_/C _21524_/B _21524_/A _21588_/X vssd1 vssd1 vccd1 vccd1 _21589_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_149_87 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14130_ _14130_/A _14130_/B _14130_/C vssd1 vssd1 vccd1 vccd1 _14131_/A sky130_fd_sc_hd__nand3_1
XFILLER_152_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23328_ _23430_/CLK _23328_/D vssd1 vssd1 vccd1 vccd1 _23328_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_153_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14061_ _14061_/A vssd1 vssd1 vccd1 vccd1 _14061_/X sky130_fd_sc_hd__clkbuf_2
X_23259_ _23259_/A vssd1 vssd1 vccd1 vccd1 _23580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input50_A x[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13012_ _12748_/X _20479_/A _13014_/A vssd1 vssd1 vccd1 vccd1 _20498_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__12713__A2 _12601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17820_ _18253_/B _18256_/A _18253_/A vssd1 vssd1 vccd1 vccd1 _17820_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13276__A _23476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17971__A _19534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23538__CLK _23538_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17751_ _17751_/A _17751_/B _17751_/C vssd1 vssd1 vccd1 vccd1 _17773_/B sky130_fd_sc_hd__nand3_2
XFILLER_130_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21493__A _21493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_14963_ _15289_/C _14962_/A _14960_/A _14960_/B vssd1 vssd1 vccd1 vccd1 _14964_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_102_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16702_ _16662_/Y _16663_/X _16457_/D _17388_/A vssd1 vssd1 vccd1 vccd1 _16707_/A
+ sky130_fd_sc_hd__o211ai_1
X_13914_ _13914_/A vssd1 vssd1 vccd1 vccd1 _13933_/A sky130_fd_sc_hd__buf_2
X_17682_ _17682_/A _17682_/B vssd1 vssd1 vccd1 vccd1 _17703_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14894_ _14756_/B _15000_/A _14890_/A _14457_/A _15004_/A vssd1 vssd1 vccd1 vccd1
+ _14896_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19421_ _19399_/A _19399_/B _19399_/C _19420_/Y vssd1 vssd1 vccd1 vccd1 _19422_/A
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__14819__B _23504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16633_ _17431_/A _16632_/X _16628_/Y vssd1 vssd1 vccd1 vccd1 _16637_/A sky130_fd_sc_hd__o21ai_1
XFILLER_74_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_398 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13845_ _22420_/A _21815_/B _21815_/C vssd1 vssd1 vccd1 vccd1 _13848_/A sky130_fd_sc_hd__or3_1
XANTENNA__15966__A2 _16153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15820__D1 _16462_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19352_ _19735_/A _19325_/Y _19345_/X _19346_/Y vssd1 vssd1 vccd1 vccd1 _19353_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_16564_ _16564_/A _16564_/B vssd1 vssd1 vccd1 vccd1 _16565_/C sky130_fd_sc_hd__nand2_1
XFILLER_62_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17168__A1 _16934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13776_ _13776_/A _13776_/B vssd1 vssd1 vccd1 vccd1 _13776_/Y sky130_fd_sc_hd__nand2_2
X_18303_ _18267_/Y _18297_/X _18417_/D _18314_/C _18302_/Y vssd1 vssd1 vccd1 vccd1
+ _18362_/A sky130_fd_sc_hd__o2111ai_1
X_15515_ _15517_/A _15540_/A _15516_/A vssd1 vssd1 vccd1 vccd1 _15515_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19283_ _19281_/X _19294_/C _19294_/D _19282_/Y _23544_/Q vssd1 vssd1 vccd1 vccd1
+ _19283_/X sky130_fd_sc_hd__a41o_1
XANTENNA__18952__D _18952_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12727_ _12712_/X _12704_/A _12726_/Y vssd1 vssd1 vccd1 vccd1 _12728_/B sky130_fd_sc_hd__o21ai_4
X_16495_ _16482_/X _16495_/B _16495_/C vssd1 vssd1 vccd1 vccd1 _16566_/C sky130_fd_sc_hd__nand3b_1
X_18234_ _18233_/Y _18227_/B _18179_/D _18185_/B vssd1 vssd1 vccd1 vccd1 _18236_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_176_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15446_ _15446_/A _15446_/B _15446_/C _15446_/D vssd1 vssd1 vccd1 vccd1 _15446_/X
+ sky130_fd_sc_hd__and4_1
X_12658_ _12577_/A _20639_/A _12580_/A _12640_/A vssd1 vssd1 vccd1 vccd1 _20675_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18165_ _18165_/A _18165_/B vssd1 vssd1 vccd1 vccd1 _18176_/A sky130_fd_sc_hd__nor2_1
XFILLER_129_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ _11828_/B vssd1 vssd1 vccd1 vccd1 _19156_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_156_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15377_ _15377_/A _15377_/B vssd1 vssd1 vccd1 vccd1 _15377_/X sky130_fd_sc_hd__xor2_1
XFILLER_8_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12589_ _20532_/A _20532_/B vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__nand2_4
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ _19494_/D _17243_/B _17107_/A _17112_/A vssd1 vssd1 vccd1 vccd1 _17301_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14328_ _13914_/A _14263_/Y _14260_/Y vssd1 vssd1 vccd1 vccd1 _14340_/A sky130_fd_sc_hd__o21ai_1
X_18096_ _18096_/A vssd1 vssd1 vccd1 vccd1 _18097_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17047_ _17047_/A _17047_/B _17047_/C vssd1 vssd1 vccd1 vccd1 _17089_/A sky130_fd_sc_hd__nand3_2
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14259_ _13965_/X _13966_/X _14261_/A _13972_/A vssd1 vssd1 vccd1 vccd1 _14330_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_143_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17628__C1 _19840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21975__A1 _21976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15103__B1 _15175_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12090__A _12090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18998_ _11841_/A _18998_/B _18998_/C _18998_/D vssd1 vssd1 vccd1 vccd1 _18999_/A
+ sky130_fd_sc_hd__nand4b_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12468__A1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17949_ _17949_/A _17949_/B vssd1 vssd1 vccd1 vccd1 _18139_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12468__B2 _18675_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16497__A _16497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20960_ _20962_/A _21079_/A _20962_/C vssd1 vssd1 vccd1 vccd1 _20960_/Y sky130_fd_sc_hd__nand3_4
XFILLER_26_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19619_ _19764_/A vssd1 vssd1 vccd1 vccd1 _19932_/A sky130_fd_sc_hd__clkbuf_2
X_20891_ _20890_/B _21124_/A _20890_/A vssd1 vssd1 vccd1 vccd1 _20989_/B sky130_fd_sc_hd__a21oi_1
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15811__D1 _15974_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22630_ _22813_/A vssd1 vssd1 vccd1 vccd1 _22630_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14090__B1 _14089_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22561_ _22637_/C _22636_/C _22641_/B _22800_/B vssd1 vssd1 vccd1 vccd1 _22650_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__16367__C1 _15964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16906__A1 _16360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21512_ _21544_/A _21512_/B vssd1 vssd1 vccd1 vccd1 _21517_/A sky130_fd_sc_hd__xnor2_1
XFILLER_139_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22492_ _22545_/B _22544_/A _22493_/C vssd1 vssd1 vccd1 vccd1 _22500_/B sky130_fd_sc_hd__a21o_1
XFILLER_166_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19305__C1 _19652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21443_ _21292_/Y _21433_/A _21453_/C vssd1 vssd1 vccd1 vccd1 _21445_/A sky130_fd_sc_hd__o21ai_1
XFILLER_194_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12265__A _18952_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12943__A2 _13177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21374_ _13177_/A _21176_/C _21635_/B _21373_/Y _21285_/Y vssd1 vssd1 vccd1 vccd1
+ _21376_/A sky130_fd_sc_hd__o311a_1
XANTENNA__16134__A2 _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19871__A3 _19304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20325_ _20325_/A _20376_/A vssd1 vssd1 vccd1 vccd1 _20329_/B sky130_fd_sc_hd__or2_2
XFILLER_162_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23113_ _23169_/A vssd1 vssd1 vccd1 vccd1 _23182_/S sky130_fd_sc_hd__buf_2
XFILLER_162_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23044_ _23044_/A vssd1 vssd1 vccd1 vccd1 _23350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20256_ _20207_/A _20117_/X _20207_/C _20196_/C _20031_/X vssd1 vssd1 vccd1 vccd1
+ _20256_/X sky130_fd_sc_hd__a41o_1
XFILLER_135_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22758__A3 _22566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13096__A _21455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_67 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20187_ _20113_/A _20112_/B _20112_/A vssd1 vssd1 vccd1 vccd1 _20188_/A sky130_fd_sc_hd__a21boi_2
XFILLER_103_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12459__A1 _12104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13120__A2 _13121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _16808_/A _11960_/B vssd1 vssd1 vccd1 vccd1 _11961_/A sky130_fd_sc_hd__nand2_2
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11682__A2 _11852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _11891_/A _11891_/B vssd1 vssd1 vccd1 vccd1 _11891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ _13630_/A _13630_/B vssd1 vssd1 vccd1 vccd1 _13630_/Y sky130_fd_sc_hd__nor2_2
XFILLER_60_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22828_ _22828_/A _22828_/B vssd1 vssd1 vccd1 vccd1 _22828_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__22143__A1 _22028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13561_ _13561_/A vssd1 vssd1 vccd1 vccd1 _13709_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22759_ _22759_/A _22759_/B vssd1 vssd1 vccd1 vccd1 _22762_/B sky130_fd_sc_hd__nand2_1
XFILLER_198_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14655__A _14655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15300_ _15300_/A _15388_/B vssd1 vssd1 vccd1 vccd1 _15330_/A sky130_fd_sc_hd__xnor2_2
XFILLER_197_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12512_ _16807_/A _23260_/B vssd1 vssd1 vccd1 vccd1 _12513_/A sky130_fd_sc_hd__nand2_2
XFILLER_185_524 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16280_ _16276_/A _16106_/Y _16581_/A vssd1 vssd1 vccd1 vccd1 _16282_/B sky130_fd_sc_hd__o21ai_1
X_13492_ _13492_/A vssd1 vssd1 vccd1 vccd1 _13553_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16373__A2 _15698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14374__B _15195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17388__D _17898_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15231_ _15231_/A _15293_/A _15231_/C _15054_/A vssd1 vssd1 vccd1 vccd1 _15293_/B
+ sky130_fd_sc_hd__nor4b_2
XFILLER_185_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16292__D _17326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12443_ _12443_/A _12443_/B _12443_/C vssd1 vssd1 vccd1 vccd1 _12444_/A sky130_fd_sc_hd__nand3_1
XFILLER_166_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19311__A2 _19304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15162_ _15162_/A _15228_/B vssd1 vssd1 vccd1 vccd1 _15191_/B sky130_fd_sc_hd__and2_1
XFILLER_176_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12374_ _12374_/A vssd1 vssd1 vccd1 vccd1 _19082_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_966 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14136__A1 _14181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14113_ _15001_/A _14026_/X _15231_/A _14110_/X _14112_/Y vssd1 vssd1 vccd1 vccd1
+ _14130_/A sky130_fd_sc_hd__o32ai_1
XFILLER_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19970_ _20142_/A _20268_/C _20146_/B _20142_/D vssd1 vssd1 vccd1 vccd1 _19980_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_153_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15093_ _15093_/A _15093_/B vssd1 vssd1 vccd1 vccd1 _15129_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__14687__A2 _14672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18921_ _18921_/A _19443_/A vssd1 vssd1 vccd1 vccd1 _19107_/C sky130_fd_sc_hd__nand2_1
X_14044_ _14193_/D _14044_/B vssd1 vssd1 vccd1 vccd1 _14050_/A sky130_fd_sc_hd__nor2_1
XFILLER_140_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18852_ _18959_/A _18959_/B _18852_/C _18959_/C vssd1 vssd1 vccd1 vccd1 _18862_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_122_874 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13437__C _13804_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17803_ _17798_/X _17799_/Y _17779_/Y _17786_/Y vssd1 vssd1 vccd1 vccd1 _17803_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18783_ _18784_/A _18784_/B _18784_/C vssd1 vssd1 vccd1 vccd1 _18785_/A sky130_fd_sc_hd__a21o_1
XFILLER_95_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23208__A _23254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15995_ _15995_/A _16181_/A _16181_/B vssd1 vssd1 vccd1 vccd1 _16000_/C sky130_fd_sc_hd__nand3_1
XANTENNA__22112__A _22112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17734_ _17250_/X _17249_/X _20317_/B _17845_/D vssd1 vssd1 vccd1 vccd1 _17734_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_94_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14946_ _14855_/Y _14856_/X _14825_/B _14941_/Y _14945_/Y vssd1 vssd1 vccd1 vccd1
+ _14953_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__17389__A1 _12323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16110__A _16549_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17665_ _17806_/B _17556_/X _17559_/Y _17666_/A _17666_/B vssd1 vssd1 vccd1 vccd1
+ _17670_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14877_ _14883_/C _14883_/A _15114_/B _15112_/D vssd1 vssd1 vccd1 vccd1 _14889_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19404_ _19242_/Y _19226_/A _19240_/Y _19239_/X vssd1 vssd1 vccd1 vccd1 _19404_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_16616_ _12509_/A _16370_/A _16635_/A vssd1 vssd1 vccd1 vccd1 _16837_/A sky130_fd_sc_hd__o21ai_1
X_13828_ _13818_/A _13818_/B _13826_/X vssd1 vssd1 vccd1 vccd1 _21786_/B sky130_fd_sc_hd__a21oi_2
XFILLER_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17596_ _17591_/X _17593_/X _17605_/A _17595_/X _17605_/B vssd1 vssd1 vccd1 vccd1
+ _17760_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19535__C1 _19700_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19335_ _19335_/A _19335_/B vssd1 vssd1 vccd1 vccd1 _19335_/Y sky130_fd_sc_hd__nand2_1
X_16547_ _16528_/A _16544_/A _16546_/X _16066_/A _16458_/X vssd1 vssd1 vccd1 vccd1
+ _16554_/A sky130_fd_sc_hd__a2111o_1
XFILLER_16_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13759_ _13759_/A _13759_/B vssd1 vssd1 vccd1 vccd1 _13763_/B sky130_fd_sc_hd__nand2_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19266_ _12353_/X _20368_/A _18928_/X _18373_/A _19082_/A vssd1 vssd1 vccd1 vccd1
+ _19266_/X sky130_fd_sc_hd__o32a_1
XANTENNA__11976__A3 _11902_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16478_ _17285_/A vssd1 vssd1 vccd1 vccd1 _16478_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_148_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18217_ _18217_/A vssd1 vssd1 vccd1 vccd1 _20317_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15429_ _15429_/A _15429_/B vssd1 vssd1 vccd1 vccd1 _15430_/B sky130_fd_sc_hd__xor2_1
XANTENNA__14375__A1 _15195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19197_ _12053_/X _11926_/X _19194_/X _19196_/Y vssd1 vssd1 vccd1 vccd1 _19197_/Y
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__12085__A _12509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16780__A _18434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19302__A2 _19172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18148_ _18148_/A _18148_/B vssd1 vssd1 vccd1 vccd1 _18149_/C sky130_fd_sc_hd__nand2_1
XANTENNA__17849__C1 _17581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18079_ _18079_/A vssd1 vssd1 vccd1 vccd1 _18272_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20110_ _20110_/A _20110_/B vssd1 vssd1 vccd1 vccd1 _20112_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21090_ _21095_/A _21212_/B _21097_/A vssd1 vssd1 vccd1 vccd1 _21090_/X sky130_fd_sc_hd__a21o_1
X_20041_ _20041_/A vssd1 vssd1 vccd1 vccd1 _23529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15627__A1 _15618_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_546 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21992_ _21992_/A _22508_/C _22226_/C vssd1 vssd1 vccd1 vccd1 _22090_/C sky130_fd_sc_hd__and3_1
XFILLER_96_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14459__B _14469_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20943_ _20943_/A _20943_/B vssd1 vssd1 vccd1 vccd1 _21057_/A sky130_fd_sc_hd__nor2_2
XFILLER_96_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _20751_/Y _20754_/X _20756_/Y vssd1 vssd1 vccd1 vccd1 _21017_/A sky130_fd_sc_hd__a21oi_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22125__A1 _22644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16674__B _19011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22613_ _22537_/X _22540_/Y _22615_/B vssd1 vssd1 vccd1 vccd1 _22619_/A sky130_fd_sc_hd__a21o_1
X_23593_ _23598_/CLK _23593_/D vssd1 vssd1 vccd1 vccd1 _23593_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22544_ _22544_/A _22544_/B vssd1 vssd1 vccd1 vccd1 _22545_/C sky130_fd_sc_hd__nand2_1
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11611__B _11611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22475_ _22475_/A _22475_/B _22475_/C _22475_/D vssd1 vssd1 vccd1 vccd1 _22501_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_154_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12377__B1 _11792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21426_ _21397_/A _21424_/X _21397_/B _21476_/A vssd1 vssd1 vccd1 vccd1 _21426_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__22833__C1 _22861_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18501__B1 _16604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21357_ _21358_/A _21358_/B _21430_/C vssd1 vssd1 vccd1 vccd1 _21433_/A sky130_fd_sc_hd__nand3_2
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_55 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20308_ _23551_/Q _20199_/B _20199_/C _20311_/B vssd1 vssd1 vccd1 vccd1 _20308_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_151_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12090_ _12090_/A vssd1 vssd1 vccd1 vccd1 _19082_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21288_ _21290_/C _21290_/B vssd1 vssd1 vccd1 vccd1 _21380_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20239_ _20236_/X _20237_/Y _20151_/D _20158_/C vssd1 vssd1 vccd1 vccd1 _20242_/B
+ sky130_fd_sc_hd__o211ai_4
X_23027_ _23027_/A vssd1 vssd1 vccd1 vccd1 _23343_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13341__A2 _13456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15079__C1 _14068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14800_ _14800_/A _14800_/B vssd1 vssd1 vccd1 vccd1 _14934_/D sky130_fd_sc_hd__nand2_1
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _15983_/A vssd1 vssd1 vccd1 vccd1 _17062_/B sky130_fd_sc_hd__buf_2
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _23457_/Q vssd1 vssd1 vccd1 vccd1 _20775_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _14731_/A vssd1 vssd1 vccd1 vccd1 _23582_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input13_A wb_dat_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _11766_/A _15882_/A _11942_/Y vssd1 vssd1 vccd1 vccd1 _11966_/A sky130_fd_sc_hd__o21ai_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12852__A1 _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _19534_/B _17450_/B _17450_/C _20317_/C vssd1 vssd1 vccd1 vccd1 _17450_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21490__B _21490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _23366_/Q _14635_/X _14661_/X vssd1 vssd1 vccd1 vccd1 _14662_/X sky130_fd_sc_hd__o21a_1
XFILLER_189_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _18503_/C _18503_/D vssd1 vssd1 vccd1 vccd1 _11875_/A sky130_fd_sc_hd__nand2_4
XANTENNA__16594__A2 _18675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _16360_/X _15884_/X _16322_/B _16389_/X _16323_/A vssd1 vssd1 vccd1 vccd1
+ _16403_/B sky130_fd_sc_hd__o221ai_1
X_13613_ _13613_/A vssd1 vssd1 vccd1 vccd1 _22126_/A sky130_fd_sc_hd__clkbuf_2
X_17381_ _17381_/A _17381_/B _17381_/C vssd1 vssd1 vccd1 vccd1 _17382_/D sky130_fd_sc_hd__nand3_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12604__A1 _12571_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14593_ _23579_/Q _14551_/X _14526_/X _12756_/B vssd1 vssd1 vccd1 vccd1 _14593_/X
+ sky130_fd_sc_hd__a22o_1
X_19120_ _19203_/A _12509_/A _18934_/Y vssd1 vssd1 vccd1 vccd1 _19121_/A sky130_fd_sc_hd__o21ai_1
XFILLER_41_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16332_ _16061_/Y _16089_/X _16330_/Y _16331_/Y vssd1 vssd1 vccd1 vccd1 _16421_/A
+ sky130_fd_sc_hd__o211ai_2
X_13544_ _13544_/A _13544_/B vssd1 vssd1 vccd1 vccd1 _13544_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19051_ _19037_/Y _19038_/Y _19066_/A _19066_/B vssd1 vssd1 vccd1 vccd1 _19058_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16263_ _16260_/Y _16261_/Y _16262_/X vssd1 vssd1 vccd1 vccd1 _16266_/B sky130_fd_sc_hd__o21ai_2
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22419__A2 _13599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13475_ _13460_/A _13460_/D _13474_/Y vssd1 vssd1 vccd1 vccd1 _13476_/C sky130_fd_sc_hd__a21o_1
XFILLER_173_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18002_ _18002_/A vssd1 vssd1 vccd1 vccd1 _18330_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15214_ _15214_/A _15214_/B vssd1 vssd1 vccd1 vccd1 _15286_/B sky130_fd_sc_hd__nand2_1
XFILLER_145_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12426_ _15718_/A _12426_/B _12426_/C vssd1 vssd1 vccd1 vccd1 _18448_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19296__A1 _19261_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16194_ _16194_/A _16194_/B _16194_/C vssd1 vssd1 vccd1 vccd1 _16194_/Y sky130_fd_sc_hd__nor3_2
XFILLER_154_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15145_ _15067_/A _15064_/X _15286_/A _15144_/X vssd1 vssd1 vccd1 vccd1 _15145_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12357_ _16500_/D vssd1 vssd1 vccd1 vccd1 _16549_/D sky130_fd_sc_hd__buf_2
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output81_A _14579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15857__B2 _15856_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19953_ _19953_/A vssd1 vssd1 vccd1 vccd1 _20366_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_141_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15076_ _15077_/A _15077_/B _15077_/C vssd1 vssd1 vccd1 vccd1 _15076_/Y sky130_fd_sc_hd__a21oi_1
X_12288_ _12288_/A _12288_/B _12288_/C vssd1 vssd1 vccd1 vccd1 _12364_/B sky130_fd_sc_hd__nand3_1
X_18904_ _18904_/A _18904_/B vssd1 vssd1 vccd1 vccd1 _18904_/Y sky130_fd_sc_hd__nand2_1
X_14027_ _14027_/A vssd1 vssd1 vccd1 vccd1 _14086_/A sky130_fd_sc_hd__clkbuf_2
X_19884_ _19835_/Y _19836_/Y _19882_/X _19827_/A vssd1 vssd1 vccd1 vccd1 _19884_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17862__C _17959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1042 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23583__D _23583_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18835_ _18835_/A vssd1 vssd1 vccd1 vccd1 _19656_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18766_ _18932_/A _18932_/B _12353_/A _18604_/X _18759_/Y vssd1 vssd1 vccd1 vccd1
+ _18767_/C sky130_fd_sc_hd__o221ai_4
X_15978_ _19017_/D _16314_/B _16314_/C vssd1 vssd1 vccd1 vccd1 _15979_/B sky130_fd_sc_hd__and3_1
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17717_ _16408_/X _17506_/A _17724_/A vssd1 vssd1 vccd1 vccd1 _17717_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__19220__A1 _19012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14929_ _14789_/A _14857_/B _14789_/C vssd1 vssd1 vccd1 vccd1 _14929_/Y sky130_fd_sc_hd__a21oi_1
X_18697_ _18880_/A _18773_/A _18753_/B vssd1 vssd1 vccd1 vccd1 _18697_/X sky130_fd_sc_hd__and3_1
XFILLER_91_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16034__B2 _15749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17648_ _17792_/A _17788_/A _17649_/C vssd1 vssd1 vccd1 vccd1 _17657_/B sky130_fd_sc_hd__a21o_1
XFILLER_1_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14596__A1 _13802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17579_ _16479_/X _17565_/X _17433_/X _17437_/X vssd1 vssd1 vccd1 vccd1 _17580_/B
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__12808__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19318_ _19302_/Y _19303_/Y _19316_/Y _19317_/X vssd1 vssd1 vccd1 vccd1 _19350_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_17_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21866__B1 _21861_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20590_ _20588_/Y _20589_/X _20576_/Y vssd1 vssd1 vccd1 vccd1 _21008_/A sky130_fd_sc_hd__o21bai_2
XFILLER_176_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19249_ _18880_/Y _18773_/C _18773_/D _18882_/Y vssd1 vssd1 vccd1 vccd1 _19249_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22260_ _22208_/X _22209_/X _22210_/Y _22216_/X vssd1 vssd1 vccd1 vccd1 _22260_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21211_ _21211_/A _21211_/B vssd1 vssd1 vccd1 vccd1 _21212_/D sky130_fd_sc_hd__nand2_1
X_22191_ _22191_/A _22191_/B vssd1 vssd1 vccd1 vccd1 _22554_/A sky130_fd_sc_hd__nand2_2
XFILLER_172_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21142_ _21542_/A _21345_/A _21344_/A _21344_/B vssd1 vssd1 vccd1 vccd1 _21142_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_133_958 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12262__B _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21073_ _21172_/A _21299_/A _21500_/A _12979_/A vssd1 vssd1 vccd1 vccd1 _21073_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23493__D _23505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20024_ _20021_/A _20023_/Y _20184_/B _20184_/A vssd1 vssd1 vccd1 vccd1 _20025_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_141_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16669__B _16669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input5_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19211__A1 _19012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21975_ _21976_/C _21976_/A _23272_/Q vssd1 vssd1 vccd1 vccd1 _21975_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ _20934_/A _20934_/B _20940_/B vssd1 vssd1 vccd1 vccd1 _20926_/Y sky130_fd_sc_hd__o21ai_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_783 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ _20860_/A vssd1 vssd1 vccd1 vccd1 _20857_/Y sky130_fd_sc_hd__inv_2
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23576_ _23578_/CLK _23576_/D vssd1 vssd1 vccd1 vccd1 _23576_/Q sky130_fd_sc_hd__dfxtp_1
X_11590_ _23598_/Q vssd1 vssd1 vccd1 vccd1 _11808_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_167_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17525__B2 _18059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20788_ _12633_/A _20786_/Y _20790_/A vssd1 vssd1 vccd1 vccd1 _20789_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__14339__A1 _14108_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22527_ _22436_/A _22436_/B _22443_/B _22729_/B vssd1 vssd1 vccd1 vccd1 _22528_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_194_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14933__A _14933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13260_ _13377_/A _13377_/D _13260_/C vssd1 vssd1 vccd1 vccd1 _13483_/B sky130_fd_sc_hd__nand3_4
X_22458_ _22417_/A _22417_/B _22417_/C _22428_/B _22428_/A vssd1 vssd1 vccd1 vccd1
+ _22516_/B sky130_fd_sc_hd__a32o_1
XFILLER_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_955 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12211_ _12211_/A _18559_/A _12211_/C vssd1 vssd1 vccd1 vccd1 _12211_/X sky130_fd_sc_hd__and3_1
XFILLER_108_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21409_ _21240_/Y _21246_/X _21340_/Y _21576_/A _21528_/C vssd1 vssd1 vccd1 vccd1
+ _21409_/X sky130_fd_sc_hd__o311a_1
XANTENNA__13562__A2 _21988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ _13191_/A _13191_/B _13191_/C _13191_/D vssd1 vssd1 vccd1 vccd1 _13191_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22389_ _22463_/B _22463_/C vssd1 vssd1 vccd1 vccd1 _22389_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _12015_/Y _12027_/Y _12141_/Y vssd1 vssd1 vccd1 vccd1 _12157_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__17963__B _18434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13268__B _13766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12172__B _16122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18778__C _18778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ _11916_/X _11947_/C _23258_/B _11961_/A vssd1 vssd1 vccd1 vccd1 _12223_/A
+ sky130_fd_sc_hd__o211ai_1
X_16950_ _16950_/A _16950_/B vssd1 vssd1 vccd1 vccd1 _16951_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20045__C1 _17414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18789__B1 _18476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15901_ _16032_/A _16033_/A _16856_/C _16856_/D vssd1 vssd1 vccd1 vccd1 _15902_/B
+ sky130_fd_sc_hd__o211ai_4
X_16881_ _16128_/X _16592_/B _16880_/X vssd1 vssd1 vccd1 vccd1 _16893_/C sky130_fd_sc_hd__a21oi_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18620_ _18620_/A vssd1 vssd1 vccd1 vccd1 _18620_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15832_ _16634_/C vssd1 vssd1 vccd1 vccd1 _16027_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22337__A1 _22756_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19202__A1 _19013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _18549_/Y _18550_/X _18547_/C vssd1 vssd1 vccd1 vccd1 _18555_/A sky130_fd_sc_hd__o21ai_1
X_15763_ _15931_/A _15761_/A _15637_/D vssd1 vssd1 vccd1 vccd1 _15763_/Y sky130_fd_sc_hd__o21ai_2
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12975_/A _12975_/B _12975_/C vssd1 vssd1 vccd1 vccd1 _12977_/B sky130_fd_sc_hd__nand3_1
XFILLER_79_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17213__B1 _23524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _17502_/A _17502_/B _17502_/C vssd1 vssd1 vccd1 vccd1 _17513_/B sky130_fd_sc_hd__nand3_1
X_14714_ _23411_/Q _14640_/A _14698_/X _23443_/Q _14713_/X vssd1 vssd1 vccd1 vccd1
+ _14714_/X sky130_fd_sc_hd__a221o_2
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _11926_/A vssd1 vssd1 vccd1 vccd1 _11926_/X sky130_fd_sc_hd__clkbuf_4
X_18482_ _18473_/X _18480_/Y _18481_/X vssd1 vssd1 vccd1 vccd1 _18482_/Y sky130_fd_sc_hd__a21boi_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ _15674_/C _15645_/A _15656_/X vssd1 vssd1 vccd1 vccd1 _15694_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17764__A1 _17644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17764__B2 _17763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_636 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17433_ _17433_/A vssd1 vssd1 vccd1 vccd1 _17433_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _23396_/Q _14640_/X _14575_/X _23428_/Q _14644_/X vssd1 vssd1 vccd1 vccd1
+ _14645_/X sky130_fd_sc_hd__a221o_1
XANTENNA__14578__A1 _13304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11857_ _11844_/A _11844_/B _19218_/A _11850_/Y _11856_/X vssd1 vssd1 vccd1 vccd1
+ _11912_/B sky130_fd_sc_hd__o311ai_4
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14578__B2 _12245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17364_ _16582_/C _16351_/Y _16761_/Y vssd1 vssd1 vccd1 vccd1 _17365_/A sky130_fd_sc_hd__o21ai_1
XFILLER_186_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14576_ input48/X _14518_/X _14545_/X _14863_/A vssd1 vssd1 vccd1 vccd1 _14576_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11788_ _11788_/A _12262_/B _18755_/A _18755_/B vssd1 vssd1 vccd1 vccd1 _11788_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12347__B _19903_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19103_ _19104_/A _19289_/B _19104_/C vssd1 vssd1 vccd1 vccd1 _19105_/A sky130_fd_sc_hd__a21oi_1
X_16315_ _16315_/A vssd1 vssd1 vccd1 vccd1 _16355_/A sky130_fd_sc_hd__clkbuf_2
X_13527_ _22392_/C vssd1 vssd1 vccd1 vccd1 _13527_/X sky130_fd_sc_hd__clkbuf_2
X_17295_ _17104_/B _17243_/X _17096_/X _17397_/A _17239_/X vssd1 vssd1 vccd1 vccd1
+ _17477_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_186_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19034_ _12243_/X _17408_/X _19031_/X _18958_/C vssd1 vssd1 vccd1 vccd1 _19035_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16246_ _16251_/B _16246_/B _16246_/C _16725_/A vssd1 vssd1 vccd1 vccd1 _16247_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_174_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13458_ _13458_/A _13458_/B _13458_/C vssd1 vssd1 vccd1 vccd1 _13463_/A sky130_fd_sc_hd__nand3_1
XANTENNA__13002__A1 _12712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19269__B2 _19265_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12356__A3 _11749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22273__B1 _22192_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ _12409_/A vssd1 vssd1 vccd1 vccd1 _18461_/B sky130_fd_sc_hd__clkbuf_2
X_16177_ _16000_/A _15990_/Y _16176_/Y vssd1 vssd1 vccd1 vccd1 _16254_/A sky130_fd_sc_hd__o21ai_2
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13389_ _22145_/C vssd1 vssd1 vccd1 vccd1 _21778_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_142_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15128_ _15130_/B _15130_/C vssd1 vssd1 vccd1 vccd1 _15129_/B sky130_fd_sc_hd__nand2_1
XFILLER_142_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18492__A2 _18474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12108__A3 _12103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19936_ _19931_/Y _19928_/C _19933_/Y _19928_/B _19935_/Y vssd1 vssd1 vccd1 vccd1
+ _20184_/B sky130_fd_sc_hd__a41oi_4
X_15059_ _15538_/C _14933_/A _14944_/B _14939_/B _15064_/A vssd1 vssd1 vccd1 vccd1
+ _15067_/C sky130_fd_sc_hd__a311o_1
XFILLER_141_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_820 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19867_ _19867_/A _19867_/B vssd1 vssd1 vccd1 vccd1 _20003_/A sky130_fd_sc_hd__nand2_2
XANTENNA__17452__B1 _17445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__A _23588_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18818_ _18818_/A vssd1 vssd1 vccd1 vccd1 _19157_/A sky130_fd_sc_hd__buf_2
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19798_ _19203_/X _17976_/A _17733_/A _19218_/X vssd1 vssd1 vccd1 vccd1 _20013_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18749_ _18749_/A vssd1 vssd1 vccd1 vccd1 _20031_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21760_ _21760_/A vssd1 vssd1 vccd1 vccd1 _21760_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_411 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20711_ _20711_/A _20718_/A vssd1 vssd1 vccd1 vccd1 _20712_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21691_ _21691_/A _21691_/B _21691_/C vssd1 vssd1 vccd1 vccd1 _21691_/X sky130_fd_sc_hd__and3_1
X_23430_ _23430_/CLK _23430_/D vssd1 vssd1 vccd1 vccd1 _23430_/Q sky130_fd_sc_hd__dfxtp_1
X_20642_ _20916_/A vssd1 vssd1 vccd1 vccd1 _20921_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20573_ _20571_/X _20572_/Y _20566_/X vssd1 vssd1 vccd1 vccd1 _20579_/B sky130_fd_sc_hd__a21oi_1
X_23361_ _23363_/CLK _23361_/D vssd1 vssd1 vccd1 vccd1 _23361_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_165_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22312_ _22314_/A _22314_/B _22323_/B vssd1 vssd1 vccd1 vccd1 _22312_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_191_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23292_ _23296_/CLK _23292_/D vssd1 vssd1 vccd1 vccd1 _23292_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__22970__A _23038_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13369__A _23471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22243_ _22439_/D _22118_/Y _22439_/C _22439_/B vssd1 vssd1 vccd1 vccd1 _22243_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_30_1166 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22174_ _22012_/Y _22171_/Y _22276_/A _22173_/Y _22487_/A vssd1 vssd1 vccd1 vccd1
+ _22174_/Y sky130_fd_sc_hd__o2111ai_4
XANTENNA__19680__B2 _19482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20921__C _21036_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21125_ _21125_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _21134_/C sky130_fd_sc_hd__nor2_1
XFILLER_105_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21056_ _21202_/B _21056_/B vssd1 vssd1 vccd1 vccd1 _21084_/C sky130_fd_sc_hd__nor2_1
XFILLER_87_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15734__D _15964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21775__C1 _22028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20007_ _20007_/A _20011_/C vssd1 vssd1 vccd1 vccd1 _20007_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19503__B _20369_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12760_ _12929_/A _20801_/C _20681_/C _12930_/A vssd1 vssd1 vccd1 vccd1 _12760_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15750__C _15860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21958_ _21820_/A _21817_/Y _21819_/B _21964_/A _21964_/B vssd1 vssd1 vccd1 vccd1
+ _21961_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18943__B1 _18755_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11918_/A _11711_/B _11711_/C vssd1 vssd1 vccd1 vccd1 _12036_/A sky130_fd_sc_hd__nand3_2
XFILLER_187_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _20906_/X _20907_/X _21054_/B _20908_/X vssd1 vssd1 vccd1 vccd1 _20909_/X
+ sky130_fd_sc_hd__o211a_1
X_12691_ _23292_/Q vssd1 vssd1 vccd1 vccd1 _20639_/D sky130_fd_sc_hd__clkinv_2
XFILLER_187_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21889_ _21984_/A _21984_/B _21984_/C _21984_/D vssd1 vssd1 vccd1 vccd1 _21893_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_43_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14430_/A _15094_/C _15238_/C _14430_/D vssd1 vssd1 vccd1 vccd1 _14456_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20727__A2_N _20726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11642_ _23583_/Q vssd1 vssd1 vccd1 vccd1 _11644_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _14361_/A _14980_/A _14361_/C _14819_/A vssd1 vssd1 vccd1 vccd1 _14361_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_35_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11573_ _11634_/A vssd1 vssd1 vccd1 vccd1 _12497_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20502__B1 _14615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23559_ _23559_/CLK _23559_/D vssd1 vssd1 vccd1 vccd1 _23559_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18171__A1 _17959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16100_ _16297_/A _16297_/B _16425_/A _16099_/Y vssd1 vssd1 vccd1 vccd1 _16340_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_7_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 wb_dat_i[1] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_4
XFILLER_161_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13312_ _13312_/A vssd1 vssd1 vccd1 vccd1 _13466_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_110 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17080_ _17221_/A _17221_/B _17221_/C vssd1 vssd1 vccd1 vccd1 _17125_/A sky130_fd_sc_hd__nand3_2
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 wb_dat_i[2] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_4
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14292_ _14292_/A _14292_/B _14292_/C vssd1 vssd1 vccd1 vccd1 _14367_/C sky130_fd_sc_hd__nand3_2
XANTENNA__15478__B _15527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_0_0_bq_clk_i_A clkbuf_2_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16031_ _16464_/A _16058_/A _16028_/A _16028_/B vssd1 vssd1 vccd1 vccd1 _16089_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__17974__A _19967_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14732__A1 _18435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ _13563_/A _21883_/B _13563_/C vssd1 vssd1 vccd1 vccd1 _13243_/Y sky130_fd_sc_hd__nand3_2
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12743__B1 _23301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19671__A1 _17643_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ _13174_/A _13174_/B vssd1 vssd1 vccd1 vccd1 _13174_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12125_ _11686_/B _11841_/Y _15905_/A _15904_/A _12118_/A vssd1 vssd1 vccd1 vccd1
+ _12125_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_151_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17982_ _17982_/A _17982_/B vssd1 vssd1 vccd1 vccd1 _17988_/D sky130_fd_sc_hd__nand2_1
XFILLER_97_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19721_ _19698_/C _19903_/A _12324_/X _18097_/A vssd1 vssd1 vccd1 vccd1 _19722_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_81_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16933_ _16924_/Y _17166_/B _16931_/X _16932_/Y vssd1 vssd1 vccd1 vccd1 _16948_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ _11998_/Y _12008_/X _12055_/Y _12033_/Y vssd1 vssd1 vccd1 vccd1 _12057_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19652_ _19652_/A vssd1 vssd1 vccd1 vccd1 _19862_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_78_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16864_ _16864_/A vssd1 vssd1 vccd1 vccd1 _16893_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18603_ _18537_/Y _18932_/A _18602_/Y vssd1 vssd1 vccd1 vccd1 _18603_/X sky130_fd_sc_hd__a21o_1
X_15815_ _15815_/A vssd1 vssd1 vccd1 vccd1 _16314_/C sky130_fd_sc_hd__buf_2
X_19583_ _19735_/A _19734_/A _19734_/B _19735_/B vssd1 vssd1 vccd1 vccd1 _19583_/Y
+ sky130_fd_sc_hd__nand4_4
X_16795_ _16795_/A _16795_/B _16795_/C _17963_/C vssd1 vssd1 vccd1 vccd1 _16808_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA__19187__B1 _19185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18534_ _11815_/A _17456_/A _18599_/A vssd1 vssd1 vccd1 vccd1 _18534_/Y sky130_fd_sc_hd__o21ai_2
X_15746_ _16070_/C _15746_/B vssd1 vssd1 vccd1 vccd1 _15746_/Y sky130_fd_sc_hd__nand2_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12958_ _12957_/Y _13151_/B _12714_/X _12950_/X vssd1 vssd1 vccd1 vccd1 _12958_/Y
+ sky130_fd_sc_hd__o31ai_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18934__B1 _17593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11909_ _12251_/A vssd1 vssd1 vccd1 vccd1 _12391_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18465_ _18465_/A vssd1 vssd1 vccd1 vccd1 _18465_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15677_ _23416_/Q vssd1 vssd1 vccd1 vccd1 _15677_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15748__B1 _15662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12358__A _12508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12889_ _12900_/A _13034_/A _12887_/X _12888_/Y vssd1 vssd1 vccd1 vccd1 _12896_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17416_ _17406_/Y _17407_/Y _17885_/A _17411_/Y _17723_/C vssd1 vssd1 vccd1 vccd1
+ _17557_/A sky130_fd_sc_hd__o2111ai_1
X_14628_ _14633_/A _18799_/B _14633_/C _14633_/B _14519_/D vssd1 vssd1 vccd1 vccd1
+ _14628_/X sky130_fd_sc_hd__a2111o_1
X_18396_ _18400_/A _18414_/C _18400_/C vssd1 vssd1 vccd1 vccd1 _18417_/A sky130_fd_sc_hd__a21o_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17347_ _17347_/A _17347_/B _17347_/C vssd1 vssd1 vccd1 vccd1 _17361_/B sky130_fd_sc_hd__nand3_4
XANTENNA__15669__A _17233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14559_ _23264_/Q _14551_/X _14698_/A _15662_/C vssd1 vssd1 vccd1 vccd1 _14559_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _17089_/A _17079_/C _17079_/D _17277_/Y vssd1 vssd1 vccd1 vccd1 _17278_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_146_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19017_ _19017_/A _19703_/D _19364_/A _19017_/D vssd1 vssd1 vccd1 vccd1 _19018_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12329__A3 _18755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16229_ _16049_/D _17625_/B _17625_/C _17420_/B _19503_/C vssd1 vssd1 vccd1 vccd1
+ _16749_/A sky130_fd_sc_hd__a32o_1
XANTENNA__13526__A2 _22558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17884__A _19951_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23594__CLK _23598_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22014__B _22364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18211__C _18211_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19919_ _19919_/A _23548_/Q _19919_/C vssd1 vssd1 vccd1 vccd1 _19923_/B sky130_fd_sc_hd__nand3_1
XFILLER_87_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17108__B _17108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18768__A3 _17444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22930_ _22930_/A vssd1 vssd1 vccd1 vccd1 _23300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21853__B _23482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16779__A2 _16278_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19323__B _20046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22861_ _22861_/A _22861_/B _22861_/C vssd1 vssd1 vccd1 vccd1 _22861_/X sky130_fd_sc_hd__and3_1
XFILLER_25_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21812_ _13834_/C _13834_/A _13834_/B _13842_/B vssd1 vssd1 vccd1 vccd1 _21812_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_37_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22792_ _22800_/A _22861_/B _22792_/C vssd1 vssd1 vccd1 vccd1 _22792_/X sky130_fd_sc_hd__and3_1
XFILLER_52_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15739__B1 _16122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21743_ _13791_/A _21896_/A _21742_/Y vssd1 vssd1 vccd1 vccd1 _21754_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12268__A _19323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21674_ _21666_/Y _21647_/Y _21646_/A _21673_/Y vssd1 vssd1 vccd1 vccd1 _21694_/A
+ sky130_fd_sc_hd__a211o_1
X_23413_ _23445_/CLK _23413_/D vssd1 vssd1 vccd1 vccd1 _23413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_983 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22485__B1 _22644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20625_ _20625_/A _20625_/B vssd1 vssd1 vccd1 vccd1 _20625_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18153__A1 _23531_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11776__A1 _11738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11900__A _18849_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23344_ _23347_/CLK _23344_/D vssd1 vssd1 vccd1 vccd1 _23344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15298__B _15298_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20556_ _20556_/A _20556_/B _20556_/C vssd1 vssd1 vccd1 vccd1 _20556_/X sky130_fd_sc_hd__and3_1
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23275_ _23559_/CLK _23275_/D vssd1 vssd1 vccd1 vccd1 _23275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20487_ _12932_/A _21061_/A _12849_/A _12571_/A vssd1 vssd1 vccd1 vccd1 _20487_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22226_ _22670_/D _22226_/B _22226_/C vssd1 vssd1 vccd1 vccd1 _22226_/X sky130_fd_sc_hd__and3_1
XFILLER_105_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22157_ _22149_/Y _22151_/Y _22154_/Y _22156_/Y vssd1 vssd1 vccd1 vccd1 _22158_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_106_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21108_ _21159_/A _21109_/A _21110_/C vssd1 vssd1 vccd1 vccd1 _21113_/A sky130_fd_sc_hd__a21o_1
XFILLER_191_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22088_ _22089_/A _22089_/B _22088_/C _22088_/D vssd1 vssd1 vccd1 vccd1 _22099_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_154_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17416__B1 _17885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13930_ _23499_/Q vssd1 vssd1 vccd1 vccd1 _14312_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21039_ _21174_/A _21039_/B _21174_/C vssd1 vssd1 vccd1 vccd1 _21040_/B sky130_fd_sc_hd__and3_1
XANTENNA__17960__C _18016_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22960__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_536 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13861_ _13861_/A _13861_/B _13861_/C vssd1 vssd1 vccd1 vccd1 _21840_/A sky130_fd_sc_hd__nand3_2
XFILLER_16_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15600_ _23420_/Q _23421_/Q vssd1 vssd1 vccd1 vccd1 _15615_/A sky130_fd_sc_hd__nor2_1
XANTENNA__17034__A _18163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ _12812_/A _12812_/B vssd1 vssd1 vccd1 vccd1 _12812_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16580_ _16581_/A _16581_/B _16581_/C vssd1 vssd1 vccd1 vccd1 _16582_/A sky130_fd_sc_hd__a21o_1
X_13792_ _22064_/A _22064_/B _21905_/B vssd1 vssd1 vccd1 vccd1 _13793_/B sky130_fd_sc_hd__nand3_2
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14377__B _15082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_bq_clk_i clkbuf_3_6_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _23566_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15531_ _15531_/A vssd1 vssd1 vccd1 vccd1 _23282_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12601_/A _12748_/A _23301_/Q vssd1 vssd1 vccd1 vccd1 _12756_/A sky130_fd_sc_hd__o21ai_1
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18250_ _18296_/A _18295_/A vssd1 vssd1 vccd1 vccd1 _18251_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _15462_/A _15462_/B _15462_/C vssd1 vssd1 vccd1 vccd1 _15467_/C sky130_fd_sc_hd__or3_1
XFILLER_30_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12674_/A vssd1 vssd1 vccd1 vccd1 _12674_/X sky130_fd_sc_hd__buf_2
XFILLER_30_425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16592__B _16592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17201_ _16663_/X _16704_/A _16969_/B vssd1 vssd1 vccd1 vccd1 _17202_/B sky130_fd_sc_hd__o21ai_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14420_/A _14352_/B _14416_/A vssd1 vssd1 vccd1 vccd1 _14415_/B sky130_fd_sc_hd__o21ai_1
X_18181_ _18182_/B _18182_/A vssd1 vssd1 vccd1 vccd1 _18185_/C sky130_fd_sc_hd__nor2_1
X_11625_ _11625_/A _11711_/B _16802_/B vssd1 vssd1 vccd1 vccd1 _12174_/A sky130_fd_sc_hd__and3_1
XFILLER_168_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15393_ _15221_/Y _15222_/Y _15282_/Y vssd1 vssd1 vccd1 vccd1 _15393_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11767__A1 _16497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17132_ _16480_/A _17304_/A _17303_/A _12311_/A vssd1 vssd1 vccd1 vccd1 _17156_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14344_ _14355_/A _14344_/B _14407_/C vssd1 vssd1 vccd1 vccd1 _14403_/D sky130_fd_sc_hd__nand3_1
XFILLER_7_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18695__A2 _17643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17063_ _17592_/A _17590_/A _16840_/A _19364_/C vssd1 vssd1 vccd1 vccd1 _17260_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14275_ _14911_/A vssd1 vssd1 vccd1 vccd1 _15225_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_170_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16014_ _16078_/A _16078_/B _16078_/C _15896_/X vssd1 vssd1 vccd1 vccd1 _16017_/B
+ sky130_fd_sc_hd__a31oi_1
X_13226_ _13259_/A vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__buf_4
XFILLER_171_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13157_ _21279_/D _13157_/B vssd1 vssd1 vccd1 vccd1 _13157_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12108_ _11844_/B _12093_/X _12103_/X _12104_/X _12107_/X vssd1 vssd1 vccd1 vccd1
+ _12491_/A sky130_fd_sc_hd__o311a_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13456__B _13456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17965_ _14729_/A _17964_/Y _17963_/C vssd1 vssd1 vccd1 vccd1 _17966_/B sky130_fd_sc_hd__o21bai_2
X_13088_ _13101_/C _13088_/B vssd1 vssd1 vccd1 vccd1 _13088_/X sky130_fd_sc_hd__and2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19704_ _19708_/B vssd1 vssd1 vccd1 vccd1 _19820_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17407__B1 _11951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21203__A1 _12785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ _15682_/A vssd1 vssd1 vccd1 vccd1 _18481_/B sky130_fd_sc_hd__clkbuf_4
X_16916_ _11871_/A _17142_/A _12051_/A _16928_/A vssd1 vssd1 vccd1 vccd1 _16923_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_78_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21203__B2 _21545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17896_ _17896_/A _17896_/B _17896_/C vssd1 vssd1 vccd1 vccd1 _17896_/Y sky130_fd_sc_hd__nand3_1
XFILLER_78_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23591__D _23591_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22951__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19635_ _19635_/A _19635_/B vssd1 vssd1 vccd1 vccd1 _23526_/D sky130_fd_sc_hd__xnor2_4
X_16847_ _17060_/A vssd1 vssd1 vccd1 vccd1 _18607_/A sky130_fd_sc_hd__buf_2
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19566_ _19528_/Y _19333_/Y _19340_/A _19345_/C vssd1 vssd1 vccd1 vccd1 _19567_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16778_ _16778_/A _16792_/A vssd1 vssd1 vccd1 vccd1 _16989_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18517_ _12465_/X _18501_/X _12463_/Y vssd1 vssd1 vccd1 vccd1 _18520_/B sky130_fd_sc_hd__o21ai_1
XFILLER_80_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15729_ _15729_/A vssd1 vssd1 vccd1 vccd1 _15729_/X sky130_fd_sc_hd__buf_2
X_19497_ _19577_/B vssd1 vssd1 vccd1 vccd1 _19521_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_80_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15197__A1 _14834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18448_ _18448_/A _18448_/B vssd1 vssd1 vccd1 vccd1 _18456_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17598__B _18093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18379_ _18378_/C _18378_/B _18378_/A vssd1 vssd1 vccd1 vccd1 _18411_/A sky130_fd_sc_hd__a21oi_1
XFILLER_175_920 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23112__C input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20410_ _20396_/Y _20397_/Y _20411_/C vssd1 vssd1 vccd1 vccd1 _20431_/B sky130_fd_sc_hd__o21bai_2
XFILLER_159_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21390_ _21391_/A _21465_/A _21391_/C vssd1 vssd1 vccd1 vccd1 _21390_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18686__A2 _17627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_986 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20341_ _20341_/A vssd1 vssd1 vccd1 vccd1 _20341_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21848__B _23482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18503__A _18503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20272_ _20269_/X _20270_/X _20271_/C _20271_/Y vssd1 vssd1 vccd1 vccd1 _20274_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_175_1029 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23060_ _14070_/X input37/X _23062_/S vssd1 vssd1 vccd1 vccd1 _23061_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22011_ _22064_/B vssd1 vssd1 vccd1 vccd1 _22564_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__13380__B1 _13379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_758 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23195__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19334__A _19334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15862__A _15862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22913_ _22913_/A vssd1 vssd1 vccd1 vccd1 _23292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13382__A _23473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22844_ _22788_/X _22805_/X _22789_/X _22812_/A vssd1 vssd1 vccd1 vccd1 _22849_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22775_ _22774_/A _22734_/A _22774_/B _22808_/A vssd1 vssd1 vccd1 vccd1 _22775_/Y
+ sky130_fd_sc_hd__o22ai_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22170__A2 _22484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11997__A1 _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21726_ _21726_/A _21726_/B vssd1 vssd1 vccd1 vccd1 _23557_/D sky130_fd_sc_hd__xnor2_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_734 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21657_ _21615_/X _21618_/Y _21619_/Y vssd1 vssd1 vccd1 vccd1 _21657_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11630__A _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20608_ _20608_/A _20608_/B _20608_/C vssd1 vssd1 vccd1 vccd1 _20610_/A sky130_fd_sc_hd__and3_1
XFILLER_177_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18677__A2 _15882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12390_ _12388_/C _12388_/A _12388_/B vssd1 vssd1 vccd1 vccd1 _12391_/A sky130_fd_sc_hd__o21ai_1
XFILLER_21_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21588_ _21521_/B _21521_/A _21568_/B vssd1 vssd1 vccd1 vccd1 _21588_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22861__C _22861_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16688__A1 _11766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23327_ _23327_/CLK _23327_/D vssd1 vssd1 vccd1 vccd1 _23327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20539_ _13051_/X _13054_/Y _20529_/A _12828_/Y vssd1 vssd1 vccd1 vccd1 _20547_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14060_ _14026_/X _14121_/A _14009_/X _14020_/Y _14039_/Y vssd1 vssd1 vccd1 vccd1
+ _14064_/B sky130_fd_sc_hd__o221ai_1
X_23258_ _23260_/A _23258_/B vssd1 vssd1 vccd1 vccd1 _23259_/A sky130_fd_sc_hd__and2_1
XANTENNA__15360__A1 _14184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13011_ _13011_/A _20798_/C _13011_/C _13011_/D vssd1 vssd1 vccd1 vccd1 _20479_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_106_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22209_ _22076_/X _22077_/Y _22074_/X vssd1 vssd1 vccd1 vccd1 _22209_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23189_ _14553_/X input18/X _23195_/S vssd1 vssd1 vccd1 vccd1 _23190_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input43_A x[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21774__A _22014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17750_ _17750_/A _17750_/B vssd1 vssd1 vccd1 vccd1 _17751_/C sky130_fd_sc_hd__nand2_1
XANTENNA__21493__B _21493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14962_ _14962_/A _14965_/B _15289_/C vssd1 vssd1 vccd1 vccd1 _14964_/A sky130_fd_sc_hd__and3_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14871__B1 _14089_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701_ _16174_/B _16168_/C _16696_/Y vssd1 vssd1 vccd1 vccd1 _16709_/A sky130_fd_sc_hd__a21oi_1
X_13913_ _14795_/A _14795_/B vssd1 vssd1 vccd1 vccd1 _13914_/A sky130_fd_sc_hd__nand2_1
X_17681_ _17523_/B _17540_/X _17686_/A vssd1 vssd1 vccd1 vccd1 _17682_/B sky130_fd_sc_hd__a21o_1
X_14893_ _14893_/A _14893_/B vssd1 vssd1 vccd1 vccd1 _14896_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19420_ _19420_/A vssd1 vssd1 vccd1 vccd1 _19420_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13292__A _23477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16632_ _15731_/A _15731_/B _16627_/A vssd1 vssd1 vccd1 vccd1 _16632_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13844_ _23480_/Q vssd1 vssd1 vccd1 vccd1 _22420_/A sky130_fd_sc_hd__clkinv_2
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15820__C1 _17259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19351_ _19339_/X _19342_/Y _19735_/A _19325_/Y vssd1 vssd1 vccd1 vccd1 _19353_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_90_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16563_ _16519_/Y _16522_/Y _16534_/Y vssd1 vssd1 vccd1 vccd1 _16565_/A sky130_fd_sc_hd__o21ai_1
X_13775_ _13768_/Y _13771_/Y _13774_/X _13632_/X vssd1 vssd1 vccd1 vccd1 _13776_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_188_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18302_ _18302_/A _18302_/B _18302_/C vssd1 vssd1 vccd1 vccd1 _18302_/Y sky130_fd_sc_hd__nand3_1
X_15514_ _15514_/A vssd1 vssd1 vccd1 vccd1 _15540_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12726_ _12644_/X _12711_/Y _12932_/A vssd1 vssd1 vccd1 vccd1 _12726_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_188_544 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19282_ _20120_/A _19924_/A _18919_/X _19443_/B _19106_/A vssd1 vssd1 vccd1 vccd1
+ _19282_/Y sky130_fd_sc_hd__o221ai_1
X_16494_ _16495_/C _16495_/B _16493_/X _16481_/X vssd1 vssd1 vccd1 vccd1 _16566_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_128_1064 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16915__A2 _16669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14835__B _15298_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18233_ _18233_/A vssd1 vssd1 vccd1 vccd1 _18233_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ _15446_/C _15370_/A _15488_/C _15488_/B vssd1 vssd1 vccd1 vccd1 _15445_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_12657_ _12724_/A vssd1 vssd1 vccd1 vccd1 _20966_/A sky130_fd_sc_hd__buf_2
XANTENNA__19314__B1 _18656_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23110__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11608_ _11608_/A vssd1 vssd1 vccd1 vccd1 _11828_/B sky130_fd_sc_hd__clkbuf_2
X_18164_ _18163_/A _18163_/B _18163_/C _18163_/D vssd1 vssd1 vccd1 vccd1 _18165_/B
+ sky130_fd_sc_hd__a22oi_1
X_15376_ _15171_/Y _15321_/B _15001_/X _15536_/B vssd1 vssd1 vccd1 vccd1 _15377_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12588_ _20493_/B _12618_/A _20493_/D _12678_/C _14655_/A vssd1 vssd1 vccd1 vccd1
+ _20532_/B sky130_fd_sc_hd__o311ai_4
XFILLER_11_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17115_ _16894_/A _16884_/Y _16878_/Y _16877_/X vssd1 vssd1 vccd1 vccd1 _17120_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_14327_ _14203_/A _14203_/B _14181_/A vssd1 vssd1 vccd1 vccd1 _14329_/A sky130_fd_sc_hd__a21o_1
X_18095_ _18101_/D _18101_/B _17752_/X _20210_/D vssd1 vssd1 vccd1 vccd1 _18095_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23586__D _23586_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17046_ _16811_/X _16814_/X _17039_/A _16627_/X vssd1 vssd1 vccd1 vccd1 _17047_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_171_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14258_ _14795_/A _14795_/B _14384_/A vssd1 vssd1 vccd1 vccd1 _14260_/A sky130_fd_sc_hd__nand3_2
XFILLER_172_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21387__C _21387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17628__B1 _17625_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11988__A1_N _15699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13467__A _13660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ _23559_/Q vssd1 vssd1 vccd1 vccd1 _13210_/C sky130_fd_sc_hd__clkinv_2
XFILLER_87_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _14189_/A _14864_/B _14864_/C _14191_/C vssd1 vssd1 vccd1 vccd1 _14199_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21975__A2 _21976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13186__B _20726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _18997_/A _18997_/B _23394_/Q _12410_/C vssd1 vssd1 vccd1 vccd1 _18998_/B
+ sky130_fd_sc_hd__nor4b_1
XANTENNA__16778__A _16778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15682__A _15682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _18058_/A _17703_/B _17703_/C _18154_/A vssd1 vssd1 vccd1 vccd1 _17948_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12468__A2 _11926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17879_ _17773_/B _17878_/Y _17747_/X vssd1 vssd1 vccd1 vccd1 _17881_/B sky130_fd_sc_hd__a21oi_1
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19618_ _19613_/Y _19615_/X _19617_/Y vssd1 vssd1 vccd1 vccd1 _19768_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__11614__B1_N _11604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20890_ _20890_/A _20890_/B _21124_/A vssd1 vssd1 vccd1 vccd1 _20989_/A sky130_fd_sc_hd__and3_1
XFILLER_0_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19002__C1 _18788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19549_ _19547_/X _19537_/X _19542_/X _19967_/A _19705_/A vssd1 vssd1 vccd1 vccd1
+ _19552_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13930__A _23499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16367__B1 _15860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22560_ _22560_/A _22560_/B vssd1 vssd1 vccd1 vccd1 _22800_/B sky130_fd_sc_hd__nand2_2
XFILLER_179_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21511_ _21463_/A _21463_/C _21463_/D _21510_/X vssd1 vssd1 vccd1 vccd1 _21512_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_55_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22491_ _21891_/A _22558_/A _22670_/A _22716_/A _22372_/X vssd1 vssd1 vccd1 vccd1
+ _22493_/C sky130_fd_sc_hd__a41o_1
XANTENNA__19305__B1 _19651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21442_ _21442_/A _21442_/B _21442_/C vssd1 vssd1 vccd1 vccd1 _21561_/A sky130_fd_sc_hd__nand3_2
XANTENNA__17316__C1 _17307_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18659__A2 _18656_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22860__B1 _22237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21373_ _20957_/X _21371_/Y _21372_/X vssd1 vssd1 vccd1 vccd1 _21373_/Y sky130_fd_sc_hd__o21ai_1
X_23112_ input40/X _23184_/B input6/X _23112_/D vssd1 vssd1 vccd1 vccd1 _23169_/A
+ sky130_fd_sc_hd__and4_1
X_20324_ _20400_/A _20400_/B _20323_/C vssd1 vssd1 vccd1 vccd1 _20376_/A sky130_fd_sc_hd__a21oi_1
XFILLER_190_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23043_ _14298_/C input7/X _23051_/S vssd1 vssd1 vccd1 vccd1 _23044_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14911__D _15075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20255_ _20255_/A _20255_/B _20255_/C vssd1 vssd1 vccd1 vccd1 _20311_/B sky130_fd_sc_hd__nand3_1
XFILLER_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21966__A2 _21981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20186_ _20186_/A _20186_/B vssd1 vssd1 vccd1 vccd1 _20189_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16842__A1 _12509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20386__B1_N _20384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13120__A3 _20905_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20003__A _20003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11890_ _19363_/A _19363_/B _16049_/D vssd1 vssd1 vccd1 vccd1 _11891_/B sky130_fd_sc_hd__and3_1
XFILLER_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22827_ _22827_/A vssd1 vssd1 vccd1 vccd1 _23571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14936__A _15044_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22143__A2 _23331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13560_ _22159_/C vssd1 vssd1 vccd1 vccd1 _21778_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_198_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22758_ _22700_/C _22566_/A _22566_/B _22701_/C _22790_/A vssd1 vssd1 vccd1 vccd1
+ _22759_/B sky130_fd_sc_hd__a32o_1
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _12511_/A vssd1 vssd1 vccd1 vccd1 _17592_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_198_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21709_ _21721_/B _21709_/B vssd1 vssd1 vccd1 vccd1 _21723_/D sky130_fd_sc_hd__nand2_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ _13491_/A vssd1 vssd1 vccd1 vccd1 _13492_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_197_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22689_ _22630_/X _22617_/A _22687_/Y vssd1 vssd1 vccd1 vccd1 _22690_/C sky130_fd_sc_hd__a21o_1
XFILLER_185_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16373__A3 _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15230_ _14834_/A _15388_/C _15228_/A _15228_/B _15227_/Y vssd1 vssd1 vccd1 vccd1
+ _15231_/C sky130_fd_sc_hd__a221oi_2
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12442_ _12130_/X _12103_/X _12425_/X _12427_/X _12429_/Y vssd1 vssd1 vccd1 vccd1
+ _12443_/C sky130_fd_sc_hd__o221ai_4
XFILLER_138_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17858__B1 _17766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15161_ _15162_/A _15228_/B vssd1 vssd1 vccd1 vccd1 _15191_/A sky130_fd_sc_hd__nor2_1
X_12373_ _12373_/A vssd1 vssd1 vccd1 vccd1 _16480_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_165_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14112_ _14858_/A _14276_/A vssd1 vssd1 vccd1 vccd1 _14112_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15092_ _15092_/A _15092_/B vssd1 vssd1 vccd1 vccd1 _15093_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_80 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18920_ _20031_/A _19107_/B _18921_/A _18919_/X vssd1 vssd1 vccd1 vccd1 _18925_/A
+ sky130_fd_sc_hd__o211ai_1
X_14043_ _23356_/Q vssd1 vssd1 vccd1 vccd1 _14193_/D sky130_fd_sc_hd__inv_2
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18851_ _18958_/B _18856_/A _18675_/B _17642_/A vssd1 vssd1 vccd1 vccd1 _18959_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_122_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23159__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17802_ _17779_/Y _17786_/Y _17796_/Y vssd1 vssd1 vccd1 vccd1 _17802_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18782_ _18627_/Y _18628_/X _18665_/Y _18666_/X vssd1 vssd1 vccd1 vccd1 _18782_/X
+ sky130_fd_sc_hd__o211a_2
X_15994_ _15995_/A _16181_/A _15993_/X _15969_/X vssd1 vssd1 vccd1 vccd1 _16000_/B
+ sky130_fd_sc_hd__o2bb2ai_2
X_17733_ _17733_/A vssd1 vssd1 vccd1 vccd1 _17980_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__13111__A3 _21177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14945_ _14947_/A _14945_/B _14945_/C vssd1 vssd1 vccd1 vccd1 _14945_/Y sky130_fd_sc_hd__nand3_1
XFILLER_85_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17664_ _17663_/Y _17497_/D _17497_/C vssd1 vssd1 vccd1 vccd1 _17670_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__21951__B _22089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14876_ _14886_/A _14876_/B _14886_/C vssd1 vssd1 vccd1 vccd1 _15000_/A sky130_fd_sc_hd__nand3_2
XFILLER_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12870__A2 _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19403_ _19401_/A _19398_/B _19402_/Y vssd1 vssd1 vccd1 vccd1 _19403_/X sky130_fd_sc_hd__a21o_1
XFILLER_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16615_ _16152_/A _16832_/A _16614_/Y vssd1 vssd1 vccd1 vccd1 _16635_/A sky130_fd_sc_hd__o21ai_1
XFILLER_51_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13827_ _13495_/X _13431_/A _13825_/Y _13818_/A _13826_/X vssd1 vssd1 vccd1 vccd1
+ _21786_/A sky130_fd_sc_hd__o311a_1
X_17595_ _17595_/A vssd1 vssd1 vccd1 vccd1 _17595_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__14072__A1 _14070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19535__B1 _11849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19334_ _19334_/A _19539_/A _19539_/B vssd1 vssd1 vccd1 vccd1 _19335_/B sky130_fd_sc_hd__and3_1
X_13758_ _13593_/X _13698_/Y _13754_/Y _13757_/Y vssd1 vssd1 vccd1 vccd1 _13759_/B
+ sky130_fd_sc_hd__o211ai_1
X_16546_ _11726_/A _11726_/B _15731_/A _15731_/B vssd1 vssd1 vccd1 vccd1 _16546_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12709_ _12709_/A vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__clkbuf_4
X_19265_ _19082_/B _20366_/B _12353_/X _20368_/A vssd1 vssd1 vccd1 vccd1 _19265_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_188_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16477_ _16471_/Y _16477_/B _16477_/C vssd1 vssd1 vccd1 vccd1 _16495_/C sky130_fd_sc_hd__nand3b_1
X_13689_ _22508_/C vssd1 vssd1 vccd1 vccd1 _22713_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18216_ _17959_/A _17959_/B _18218_/A _20212_/D _18219_/D vssd1 vssd1 vccd1 vccd1
+ _18279_/A sky130_fd_sc_hd__a32o_1
XFILLER_15_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15428_ _15463_/B _15463_/A vssd1 vssd1 vccd1 vccd1 _15429_/B sky130_fd_sc_hd__xnor2_1
X_19196_ _19196_/A _19196_/B _19196_/C vssd1 vssd1 vccd1 vccd1 _19196_/Y sky130_fd_sc_hd__nor3_2
XANTENNA__11701__C _16674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20583__A _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16780__B _16780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17849__B1 _17605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18147_ _17942_/A _23529_/Q _17942_/C _18145_/Y _18146_/Y vssd1 vssd1 vccd1 vccd1
+ _18149_/A sky130_fd_sc_hd__a32oi_1
XFILLER_156_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15359_ _15488_/A vssd1 vssd1 vccd1 vccd1 _15536_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18078_ _20217_/A vssd1 vssd1 vccd1 vccd1 _20269_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_116_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17029_ _17029_/A vssd1 vssd1 vccd1 vccd1 _17029_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20040_ _20201_/B _20040_/B vssd1 vssd1 vccd1 vccd1 _20041_/A sky130_fd_sc_hd__and2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16824__A1 _16447_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15627__A2 _15621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21991_ _21829_/A _13553_/X _21983_/X _21893_/A _21984_/Y vssd1 vssd1 vccd1 vccd1
+ _22090_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16037__C1 _15704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14459__C _15233_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20942_ _20947_/B vssd1 vssd1 vccd1 vccd1 _21057_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16588__B1 _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20873_ _20751_/B _20751_/A _21157_/C _21157_/D _21157_/B vssd1 vssd1 vccd1 vccd1
+ _21017_/C sky130_fd_sc_hd__o2111ai_4
XANTENNA__22125__A2 _13431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16674__C _17108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13660__A _13660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22612_ _22631_/A _22631_/B _22611_/X vssd1 vssd1 vccd1 vccd1 _22615_/B sky130_fd_sc_hd__o21ai_2
X_23592_ _23598_/CLK _23592_/D vssd1 vssd1 vccd1 vccd1 _23592_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__17001__A1 _17217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22543_ _13547_/X _22484_/X _22362_/B _22496_/B vssd1 vssd1 vccd1 vccd1 _22544_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_167_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13810__D _22159_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23528__CLK _23538_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22474_ _22474_/A _22757_/B _22474_/C vssd1 vssd1 vccd1 vccd1 _22475_/A sky130_fd_sc_hd__or3_1
XFILLER_148_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12377__A1 _11931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12377__B2 _11792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21425_ _21397_/A _21397_/B _21424_/X vssd1 vssd1 vccd1 vccd1 _21425_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18501__A1 _11760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21356_ _21356_/A vssd1 vssd1 vccd1 vccd1 _21635_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20307_ _20307_/A _20307_/B _20307_/C _20452_/B vssd1 vssd1 vccd1 vccd1 _20354_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_190_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21287_ _21187_/A _21173_/X _21210_/B vssd1 vssd1 vccd1 vccd1 _21290_/B sky130_fd_sc_hd__o21ai_1
XFILLER_146_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23026_ _23343_/Q input24/X _23034_/S vssd1 vssd1 vccd1 vccd1 _23027_/A sky130_fd_sc_hd__mux2_1
X_20238_ _20151_/D _20158_/C _20236_/X _20237_/Y vssd1 vssd1 vccd1 vccd1 _20290_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15079__B1 _15054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20169_ _20171_/B vssd1 vssd1 vccd1 vccd1 _20283_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _12991_/A _12991_/B _12991_/C vssd1 vssd1 vccd1 vccd1 _20585_/B sky130_fd_sc_hd__nand3_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14730_ _16800_/D _16807_/B _16815_/D _14730_/D vssd1 vssd1 vccd1 vccd1 _14731_/A
+ sky130_fd_sc_hd__and4_1
X_11942_ _12167_/A _12168_/A _18503_/A _18503_/B vssd1 vssd1 vccd1 vccd1 _11942_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_55_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19053__A2_N _18840_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12852__A2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _23334_/Q _14636_/X _14642_/X _23302_/Q _14657_/X vssd1 vssd1 vccd1 vccd1
+ _14661_/X sky130_fd_sc_hd__a221o_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11873_ _11887_/A vssd1 vssd1 vccd1 vccd1 _18503_/D sky130_fd_sc_hd__clkbuf_4
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22116__A2 _22112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _12279_/A _16398_/X _16364_/X _16399_/X vssd1 vssd1 vccd1 vccd1 _16403_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_13612_ _13552_/A _13599_/X _13627_/A vssd1 vssd1 vccd1 vccd1 _13619_/A sky130_fd_sc_hd__o21ai_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _23525_/Q _17380_/B vssd1 vssd1 vccd1 vccd1 _17533_/A sky130_fd_sc_hd__nand2_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _23422_/Q vssd1 vssd1 vccd1 vccd1 _15664_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16331_ _16331_/A _16331_/B vssd1 vssd1 vccd1 vccd1 _16331_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13543_ _13541_/X _13542_/Y _13540_/B vssd1 vssd1 vccd1 vccd1 _13543_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__11958__A4 _16141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19050_ _19041_/X _19042_/X _19052_/A vssd1 vssd1 vccd1 vccd1 _19066_/B sky130_fd_sc_hd__o21ai_1
X_16262_ _15946_/Y _15947_/X _15950_/Y _16268_/A vssd1 vssd1 vccd1 vccd1 _16262_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_146_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13474_ _13474_/A _13474_/B vssd1 vssd1 vccd1 vccd1 _13474_/Y sky130_fd_sc_hd__nand2_1
X_18001_ _20081_/B vssd1 vssd1 vccd1 vccd1 _18001_/X sky130_fd_sc_hd__clkbuf_2
X_15213_ _15214_/B _15214_/A vssd1 vssd1 vccd1 vccd1 _15213_/Y sky130_fd_sc_hd__nor2_1
X_12425_ _12425_/A vssd1 vssd1 vccd1 vccd1 _12425_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16193_ _12373_/A _16662_/A _16194_/C _16192_/X vssd1 vssd1 vccd1 vccd1 _16193_/Y
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__19296__A2 _20320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15928__C _15928_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15144_ _15144_/A _15144_/B vssd1 vssd1 vccd1 vccd1 _15144_/X sky130_fd_sc_hd__or2_1
X_12356_ _14735_/A _11747_/X _11749_/X _12355_/Y vssd1 vssd1 vccd1 vccd1 _12363_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19952_ _19952_/A vssd1 vssd1 vccd1 vccd1 _20043_/A sky130_fd_sc_hd__clkbuf_2
X_15075_ _15075_/A _15075_/B vssd1 vssd1 vccd1 vccd1 _15077_/C sky130_fd_sc_hd__nand2_1
X_12287_ _12297_/B _12297_/C _12287_/C vssd1 vssd1 vccd1 vccd1 _12288_/C sky130_fd_sc_hd__nand3_1
XFILLER_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18903_ _18903_/A _18903_/B vssd1 vssd1 vccd1 vccd1 _18903_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14026_ _14054_/A vssd1 vssd1 vccd1 vccd1 _14026_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_output74_A _14711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23219__A _23241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19883_ _19827_/A _19830_/A _19882_/X vssd1 vssd1 vccd1 vccd1 _19883_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18958__D _19674_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20063__B1 _17565_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13167__D _21279_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16806__A1 _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17217__A _17217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_823 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18834_ _11822_/X _19196_/B _18825_/A vssd1 vssd1 vccd1 vccd1 _18841_/A sky130_fd_sc_hd__o21ai_1
XFILLER_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23001__A0 _22142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21962__A _22118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18765_ _18765_/A _18765_/B vssd1 vssd1 vccd1 vccd1 _18767_/B sky130_fd_sc_hd__nand2_1
X_15977_ _15843_/B _16123_/A _16172_/A vssd1 vssd1 vccd1 vccd1 _15982_/A sky130_fd_sc_hd__o21ai_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17716_ _17628_/Y _17712_/Y _17714_/A vssd1 vssd1 vccd1 vccd1 _17724_/A sky130_fd_sc_hd__o21ai_1
X_14928_ _14928_/A _14928_/B vssd1 vssd1 vccd1 vccd1 _14928_/X sky130_fd_sc_hd__xor2_1
X_18696_ _18880_/A _18773_/A _18753_/B vssd1 vssd1 vccd1 vccd1 _18696_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17647_ _12237_/X _18276_/C _17646_/X _17420_/Y vssd1 vssd1 vccd1 vccd1 _17649_/C
+ sky130_fd_sc_hd__o31ai_2
XFILLER_91_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14859_ _15155_/A _14980_/A vssd1 vssd1 vccd1 vccd1 _14874_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17578_ _17578_/A _17578_/B _17578_/C vssd1 vssd1 vccd1 vccd1 _17609_/A sky130_fd_sc_hd__nand3_4
XANTENNA__13911__C _13911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12808__B _20969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19317_ _19320_/A _19321_/A _19517_/B vssd1 vssd1 vccd1 vccd1 _19317_/X sky130_fd_sc_hd__and3_1
X_16529_ _16529_/A _16549_/A _16529_/C _16544_/B vssd1 vssd1 vccd1 vccd1 _16530_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_17_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16791__A _16988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19248_ _19236_/Y _19245_/X _19254_/A vssd1 vssd1 vccd1 vccd1 _19434_/A sky130_fd_sc_hd__a21o_1
XFILLER_192_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12359__A1 _14735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19179_ _19007_/Y _19177_/Y _19047_/C _19178_/Y vssd1 vssd1 vccd1 vccd1 _19179_/Y
+ sky130_fd_sc_hd__o211ai_4
X_21210_ _21290_/C _21210_/B vssd1 vssd1 vccd1 vccd1 _21211_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22190_ _21902_/B _22028_/A _22141_/D _21853_/A vssd1 vssd1 vccd1 vccd1 _22191_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__19029__D _19029_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21141_ _21414_/A _21415_/A _21344_/A _21344_/B vssd1 vssd1 vccd1 vccd1 _21141_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18511__A _18511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12262__C _12306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21072_ _21072_/A vssd1 vssd1 vccd1 vccd1 _21500_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20023_ _20113_/A vssd1 vssd1 vccd1 vccd1 _20023_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22968__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21974_ _22107_/B _22107_/C _21973_/C _21980_/A vssd1 vssd1 vccd1 vccd1 _21976_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_656 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20925_ _21281_/A _21282_/A _21174_/B vssd1 vssd1 vccd1 vccd1 _20940_/B sky130_fd_sc_hd__and3_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20856_ _20856_/A _20856_/B _20856_/C vssd1 vssd1 vccd1 vccd1 _20860_/A sky130_fd_sc_hd__nand3_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23575_ _23575_/CLK _23575_/D vssd1 vssd1 vccd1 vccd1 _23575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20787_ _20783_/A _20783_/B _20920_/A _20778_/A vssd1 vssd1 vccd1 vccd1 _20790_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_195_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22526_ _22538_/B _22443_/B _22729_/B vssd1 vssd1 vccd1 vccd1 _22528_/A sky130_fd_sc_hd__a21o_1
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14933__B _23505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22457_ _22457_/A _22457_/B vssd1 vssd1 vccd1 vccd1 _22524_/B sky130_fd_sc_hd__nand2_1
XFILLER_148_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12210_ _12211_/A _18559_/A _12211_/C vssd1 vssd1 vccd1 vccd1 _12210_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21408_ _21411_/A _21411_/B vssd1 vssd1 vccd1 vccd1 _21528_/C sky130_fd_sc_hd__or2_1
XFILLER_109_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13190_ _13174_/A _13169_/C _13169_/D _13169_/B vssd1 vssd1 vccd1 vccd1 _13191_/B
+ sky130_fd_sc_hd__a22o_1
X_22388_ _22553_/A _22388_/B _22388_/C vssd1 vssd1 vccd1 vccd1 _22463_/C sky130_fd_sc_hd__and3_1
XANTENNA__13562__A3 _21778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20951__A _20984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12141_ _11998_/Y _12008_/X _12033_/Y vssd1 vssd1 vccd1 vccd1 _12141_/Y sky130_fd_sc_hd__o21ai_1
X_21339_ _21404_/A _21402_/A _21264_/Y _21342_/C vssd1 vssd1 vccd1 vccd1 _21340_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_190_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12072_ _23256_/B _11947_/A _12070_/Y _15957_/C vssd1 vssd1 vccd1 vccd1 _12222_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20045__B1 _17414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23009_ _23009_/A vssd1 vssd1 vccd1 vccd1 _23335_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18789__B2 _18484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15900_ _11853_/A _11807_/X _15682_/B _15798_/A _15799_/A vssd1 vssd1 vccd1 vccd1
+ _16209_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16880_ _16319_/A _12208_/A _16592_/B _16128_/X vssd1 vssd1 vccd1 vccd1 _16880_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_103_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22878__A _22878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__C1 _11960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17461__A1 _17610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15831_ _15831_/A vssd1 vssd1 vccd1 vccd1 _16634_/C sky130_fd_sc_hd__clkbuf_2
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _18528_/Y _18529_/Y _18526_/Y _18519_/Y vssd1 vssd1 vccd1 vccd1 _18550_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15762_ _15762_/A _15921_/B vssd1 vssd1 vccd1 vccd1 _15762_/Y sky130_fd_sc_hd__nand2_2
X_12974_ _13141_/B _13141_/C _12973_/Y vssd1 vssd1 vccd1 vccd1 _12977_/A sky130_fd_sc_hd__a21o_1
XFILLER_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _17502_/A _17502_/B _17502_/C vssd1 vssd1 vccd1 vccd1 _17513_/A sky130_fd_sc_hd__a21o_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _23379_/Q _14635_/A _14712_/X vssd1 vssd1 vccd1 vccd1 _14713_/X sky130_fd_sc_hd__o21a_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _17626_/A vssd1 vssd1 vccd1 vccd1 _11926_/A sky130_fd_sc_hd__clkbuf_4
X_18481_ _18859_/B _18481_/B _18481_/C vssd1 vssd1 vccd1 vccd1 _18481_/X sky130_fd_sc_hd__and3_1
XFILLER_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15693_ _15686_/A _15686_/B _15672_/C _15692_/Y vssd1 vssd1 vccd1 vccd1 _15693_/Y
+ sky130_fd_sc_hd__a31oi_2
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17764__A2 _17613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17432_ _16370_/X _17733_/A _17039_/B _17439_/A vssd1 vssd1 vccd1 vccd1 _17432_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11813__A _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11856_ _12378_/A _12378_/B _11807_/X _14729_/A _18481_/C vssd1 vssd1 vccd1 vccd1
+ _11856_/X sky130_fd_sc_hd__o221a_2
X_14644_ _23364_/Q _14635_/X _14643_/X vssd1 vssd1 vccd1 vccd1 _14644_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15775__A1 _16480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17363_ _17353_/Y _17357_/Y _17362_/Y vssd1 vssd1 vccd1 vccd1 _17832_/A sky130_fd_sc_hd__o21ai_4
X_14575_ _14647_/A vssd1 vssd1 vccd1 vccd1 _14575_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11787_ _12145_/B vssd1 vssd1 vccd1 vccd1 _18755_/B sky130_fd_sc_hd__clkbuf_4
X_19102_ _18926_/A _18927_/A _19288_/C vssd1 vssd1 vccd1 vccd1 _19104_/C sky130_fd_sc_hd__o21ai_1
XFILLER_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12347__C _19261_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16314_ _19161_/A _16314_/B _16314_/C _17133_/C vssd1 vssd1 vccd1 vccd1 _16384_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_119_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13526_ _13712_/A _22558_/A _13736_/B _21891_/A vssd1 vssd1 vccd1 vccd1 _13544_/B
+ sky130_fd_sc_hd__a22o_1
X_17294_ _17397_/A _17239_/X _17397_/B vssd1 vssd1 vccd1 vccd1 _17477_/A sky130_fd_sc_hd__a21o_1
XFILLER_174_815 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22118__A _22118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18315__B _23534_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19033_ _19033_/A _19138_/B vssd1 vssd1 vccd1 vccd1 _19036_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13457_ _13425_/Y _13599_/A _22269_/C _13443_/B _21877_/A vssd1 vssd1 vccd1 vccd1
+ _13458_/B sky130_fd_sc_hd__o2111ai_1
X_16245_ _16251_/B _16246_/B _16246_/C _16725_/A vssd1 vssd1 vccd1 vccd1 _16247_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15020__A _15075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ _19155_/B _19155_/C _12410_/C _18440_/A vssd1 vssd1 vccd1 vccd1 _12409_/A
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__12210__B1 _12211_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16176_ _16139_/Y _16169_/Y _16179_/B vssd1 vssd1 vccd1 vccd1 _16176_/Y sky130_fd_sc_hd__o21ai_4
X_13388_ _22039_/C vssd1 vssd1 vccd1 vccd1 _22145_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_154_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15955__A _23589_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12339_ _12339_/A _12339_/B _12339_/C vssd1 vssd1 vccd1 vccd1 _12339_/Y sky130_fd_sc_hd__nand3_1
XFILLER_5_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15127_ _15127_/A _15188_/B _15127_/C vssd1 vssd1 vccd1 vccd1 _15130_/C sky130_fd_sc_hd__nand3_1
XFILLER_47_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18331__A _19900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18492__A3 _19670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23594__D _23594_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19935_ _19928_/B _19934_/Y _19928_/D vssd1 vssd1 vccd1 vccd1 _19935_/Y sky130_fd_sc_hd__o21ai_1
X_15058_ _15408_/A vssd1 vssd1 vccd1 vccd1 _15538_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_142_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14009_ _14135_/A vssd1 vssd1 vccd1 vccd1 _14009_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19866_ _19685_/A _19685_/B _19685_/C _19654_/X vssd1 vssd1 vccd1 vccd1 _19867_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_110_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_854 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18817_ _12432_/A _18813_/A _18998_/D vssd1 vssd1 vccd1 vccd1 _18818_/A sky130_fd_sc_hd__o21ai_1
XFILLER_110_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19797_ _19880_/A _19880_/B _19893_/B _19796_/Y vssd1 vssd1 vccd1 vccd1 _19879_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18748_ _19288_/A _19288_/B vssd1 vssd1 vccd1 vccd1 _18927_/A sky130_fd_sc_hd__and2_1
XFILLER_23_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_280 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18401__B1 _23536_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18679_ _12343_/A _19334_/A _18677_/Y _18678_/Y vssd1 vssd1 vccd1 vccd1 _18681_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20710_ _20618_/Y _20697_/Y _20700_/X _20853_/B vssd1 vssd1 vccd1 vccd1 _20717_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_91_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11723__A _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21690_ _21690_/A vssd1 vssd1 vccd1 vccd1 _23553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14456__D _15175_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20641_ _20641_/A _20660_/A vssd1 vssd1 vccd1 vccd1 _20916_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18506__A _18506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23360_ _23363_/CLK _23360_/D vssd1 vssd1 vccd1 vccd1 _23360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20572_ _20562_/B _20726_/D _20769_/A _20566_/B vssd1 vssd1 vccd1 vccd1 _20572_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_177_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22311_ _22310_/Y _22199_/A _22288_/Y _22289_/Y vssd1 vssd1 vccd1 vccd1 _22323_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_176_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12472__A1_N _12104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23291_ _23296_/CLK _23291_/D vssd1 vssd1 vccd1 vccd1 _23291_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_192_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22242_ _22242_/A _22242_/B _22242_/C vssd1 vssd1 vccd1 vccd1 _22439_/B sky130_fd_sc_hd__nand3_2
XFILLER_127_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12273__B _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19337__A _19709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22173_ _22173_/A _22279_/A vssd1 vssd1 vccd1 vccd1 _22173_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19680__A2 _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21124_ _21124_/A _21124_/B _21514_/A vssd1 vssd1 vccd1 vccd1 _21125_/B sky130_fd_sc_hd__and3_1
XANTENNA__23213__A0 _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19968__B1 _19203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21055_ _21054_/C _21169_/A _13122_/B _20471_/Y vssd1 vssd1 vccd1 vccd1 _21056_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13816__C _23475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20006_ _19876_/B _19833_/X _19939_/Y vssd1 vssd1 vccd1 vccd1 _20011_/C sky130_fd_sc_hd__a21oi_1
XFILLER_189_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19503__C _19503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22724__C1 _22237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21957_ _21957_/A _21957_/B _21957_/C vssd1 vssd1 vccd1 vccd1 _21964_/B sky130_fd_sc_hd__nand3_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15750__D _15968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11633__A _23590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _23587_/Q vssd1 vssd1 vccd1 vccd1 _11711_/C sky130_fd_sc_hd__inv_2
XFILLER_188_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19800__A _19900_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _20908_/A vssd1 vssd1 vccd1 vccd1 _20908_/X sky130_fd_sc_hd__buf_2
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20368__D _20368_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12683_/B _12712_/A _23293_/Q vssd1 vssd1 vccd1 vccd1 _12850_/B sky130_fd_sc_hd__a21oi_4
XFILLER_188_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21888_ _21984_/A _21984_/B _21984_/C _21984_/D vssd1 vssd1 vccd1 vccd1 _21893_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _12281_/A _18675_/A _11915_/A _19196_/A vssd1 vssd1 vccd1 vccd1 _11907_/B
+ sky130_fd_sc_hd__o22a_1
X_20839_ _20839_/A _20839_/B _20839_/C vssd1 vssd1 vccd1 vccd1 _20840_/A sky130_fd_sc_hd__nand3_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14360_ _14360_/A vssd1 vssd1 vccd1 vccd1 _14819_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23558_ _23558_/CLK _23558_/D vssd1 vssd1 vccd1 vccd1 _23558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11572_ _11648_/A _11918_/B _11624_/A vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__nand3_1
XFILLER_11_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20502__A1 _12601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ _21882_/C _21882_/A vssd1 vssd1 vccd1 vccd1 _13312_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20384__C _20384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 wb_dat_i[20] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22509_ _22509_/A _22509_/B _22509_/C vssd1 vssd1 vccd1 vccd1 _22509_/X sky130_fd_sc_hd__and3_1
XFILLER_196_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ _14279_/C _14279_/A _14279_/B _14358_/A _14358_/B vssd1 vssd1 vccd1 vccd1
+ _14292_/C sky130_fd_sc_hd__a32o_1
XANTENNA__16182__A1 _19161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23489_ _23499_/CLK _23501_/Q vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
XFILLER_182_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16182__B2 _12306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13242_ _23477_/Q vssd1 vssd1 vccd1 vccd1 _21883_/B sky130_fd_sc_hd__buf_2
X_16030_ _16030_/A vssd1 vssd1 vccd1 vccd1 _16058_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17974__B _20133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20681__A _21431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12183__B _12187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20266__B1 _19425_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13173_ _13171_/A _13172_/X _13169_/B _13191_/A vssd1 vssd1 vccd1 vccd1 _13174_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22007__A1 _21997_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23204__A0 _15664_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ _12022_/X _12025_/X _12029_/B _12011_/X vssd1 vssd1 vccd1 vccd1 _12399_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_124_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17981_ _17611_/X _20210_/D _17986_/D _17986_/B vssd1 vssd1 vccd1 vccd1 _17994_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19720_ _12324_/X _18097_/A _19698_/C _19903_/A vssd1 vssd1 vccd1 vccd1 _19722_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__13295__A _23478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16932_ _16590_/A _16590_/B _16600_/Y _16601_/Y vssd1 vssd1 vccd1 vccd1 _16932_/Y
+ sky130_fd_sc_hd__a22oi_4
X_12055_ _12016_/Y _12023_/Y _12054_/Y _12026_/Y vssd1 vssd1 vccd1 vccd1 _12055_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_2_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19651_ _19651_/A vssd1 vssd1 vccd1 vccd1 _19862_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16863_ _16879_/A _16879_/B _16879_/C vssd1 vssd1 vccd1 vccd1 _16864_/A sky130_fd_sc_hd__nand3_1
XANTENNA__14248__A1 _14245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18602_ _12167_/X _12168_/X _17761_/A _17761_/B vssd1 vssd1 vccd1 vccd1 _18602_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15814_ _15814_/A vssd1 vssd1 vccd1 vccd1 _16314_/B sky130_fd_sc_hd__buf_2
X_19582_ _19580_/Y _19581_/X _19476_/Y _19477_/Y vssd1 vssd1 vccd1 vccd1 _19735_/B
+ sky130_fd_sc_hd__o2bb2ai_2
X_16794_ _16817_/A _16794_/B vssd1 vssd1 vccd1 vccd1 _17043_/A sky130_fd_sc_hd__nand2_1
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18533_ _11851_/A _11852_/A _18755_/C _18755_/D vssd1 vssd1 vccd1 vccd1 _18599_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _15742_/X _16447_/B _12174_/X _12173_/X _12175_/X vssd1 vssd1 vccd1 vccd1
+ _15746_/B sky130_fd_sc_hd__o221a_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _13019_/C _12678_/Y _12640_/A vssd1 vssd1 vccd1 vccd1 _12957_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18934__A1 _12246_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18934__B2 _17591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_918 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11908_ _11908_/A _11908_/B vssd1 vssd1 vccd1 vccd1 _12251_/A sky130_fd_sc_hd__nor2_1
X_18464_ _18464_/A _18464_/B _18464_/C vssd1 vssd1 vccd1 vccd1 _18465_/A sky130_fd_sc_hd__nand3_2
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ _15712_/A vssd1 vssd1 vccd1 vccd1 _16187_/A sky130_fd_sc_hd__buf_2
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12899_/B _12899_/C _12887_/C vssd1 vssd1 vccd1 vccd1 _12888_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12358__B _16549_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _17265_/Y _17414_/X _17260_/Y vssd1 vssd1 vccd1 vccd1 _17417_/B sky130_fd_sc_hd__a21o_1
XFILLER_33_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14627_ _23394_/Q vssd1 vssd1 vccd1 vccd1 _18799_/B sky130_fd_sc_hd__clkbuf_2
X_18395_ _18395_/A _18395_/B vssd1 vssd1 vccd1 vccd1 _18400_/C sky130_fd_sc_hd__nand2_1
X_11839_ _11834_/A _11834_/B _12241_/A vssd1 vssd1 vccd1 vccd1 _11844_/A sky130_fd_sc_hd__a21o_1
XFILLER_53_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18326__A _20368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23589__D _23589_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17230__A _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17346_ _17346_/A _17346_/B vssd1 vssd1 vccd1 vccd1 _17347_/C sky130_fd_sc_hd__nand2_1
X_14558_ _23416_/Q vssd1 vssd1 vccd1 vccd1 _15662_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__15669__B _16198_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18162__A2 _17723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _21793_/A vssd1 vssd1 vccd1 vccd1 _13650_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17277_ _17047_/A _17047_/B _17047_/C vssd1 vssd1 vccd1 vccd1 _17277_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__12374__A _12374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14489_ _14486_/A _14486_/B _14486_/C _14487_/A _14487_/B vssd1 vssd1 vccd1 vccd1
+ _14496_/B sky130_fd_sc_hd__a32o_1
XANTENNA__12286__A2_N _12297_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19016_ _19148_/A _19148_/B _19148_/C vssd1 vssd1 vccd1 vccd1 _19037_/A sky130_fd_sc_hd__nand3_2
XANTENNA__21049__A2 _21174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16228_ _16662_/A vssd1 vssd1 vccd1 vccd1 _16741_/A sky130_fd_sc_hd__buf_2
XFILLER_173_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1000 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ _12086_/A _15884_/X _16157_/A vssd1 vssd1 vccd1 vccd1 _16641_/A sky130_fd_sc_hd__o21ai_1
XFILLER_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11942__C1 _18503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22014__C _22380_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18211__D _18211_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19918_ _19919_/C _19919_/A _23548_/Q vssd1 vssd1 vccd1 vccd1 _19920_/A sky130_fd_sc_hd__a21o_1
XANTENNA__17108__C _19485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19849_ _19659_/Y _20079_/A _19847_/X _19848_/Y vssd1 vssd1 vccd1 vccd1 _19855_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_110_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22860_ _22187_/A _22187_/B _22237_/X vssd1 vssd1 vccd1 vccd1 _22860_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15987__A1 _15858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19323__C _20047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21811_ _13822_/Y _13824_/Y _21807_/Y _13829_/Y vssd1 vssd1 vccd1 vccd1 _21811_/X
+ sky130_fd_sc_hd__o211a_1
X_22791_ _22800_/A _22861_/B _22762_/B _22762_/A vssd1 vssd1 vccd1 vccd1 _22791_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__22182__B1 _13430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15739__A1 _15862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21742_ _22014_/A _13804_/B _21896_/A _13791_/A vssd1 vssd1 vccd1 vccd1 _21742_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_52_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21673_ _21673_/A vssd1 vssd1 vccd1 vccd1 _21673_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17140__A _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23412_ _23444_/CLK _23412_/D vssd1 vssd1 vccd1 vccd1 _23412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20624_ _20624_/A vssd1 vssd1 vccd1 vccd1 _20624_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22981__A _23038_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23269__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11776__A2 _11740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23343_ _23343_/CLK _23343_/D vssd1 vssd1 vccd1 vccd1 _23343_/Q sky130_fd_sc_hd__dfxtp_1
X_20555_ _20547_/X _20549_/Y _20516_/A _20524_/A vssd1 vssd1 vccd1 vccd1 _20578_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_165_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14714__A2 _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23274_ _23492_/CLK _23274_/D vssd1 vssd1 vccd1 vccd1 _23274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20486_ _20625_/A _20621_/A _20485_/Y vssd1 vssd1 vccd1 vccd1 _20634_/B sky130_fd_sc_hd__o21ai_2
XFILLER_180_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22225_ _22225_/A _22231_/B _22225_/C vssd1 vssd1 vccd1 vccd1 _22225_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__18310__C1 _18417_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22156_ _13732_/A _22164_/A _22151_/Y _22155_/Y vssd1 vssd1 vccd1 vccd1 _22156_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_191_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21107_ _21115_/A _21115_/B vssd1 vssd1 vccd1 vccd1 _21110_/C sky130_fd_sc_hd__xnor2_1
XFILLER_105_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12489__B1 _12478_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22087_ _22093_/C _22093_/D _22086_/Y vssd1 vssd1 vccd1 vccd1 _22088_/D sky130_fd_sc_hd__a21bo_1
XFILLER_120_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21038_ _20934_/B _21176_/C _21184_/A vssd1 vssd1 vccd1 vccd1 _21040_/A sky130_fd_sc_hd__o21ai_1
XFILLER_75_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13860_ _13676_/A _13676_/B _13676_/C _13692_/B _13692_/C vssd1 vssd1 vccd1 vccd1
+ _13861_/C sky130_fd_sc_hd__a32o_1
XFILLER_47_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19169__A1 _11898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ _12812_/A _12812_/B _12810_/Y vssd1 vssd1 vccd1 vccd1 _12816_/B sky130_fd_sc_hd__a21oi_1
X_13791_ _13791_/A vssd1 vssd1 vccd1 vccd1 _21916_/A sky130_fd_sc_hd__clkbuf_2
X_22989_ _22989_/A vssd1 vssd1 vccd1 vccd1 _23326_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17719__A2 _17644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _15530_/A _15530_/B vssd1 vssd1 vccd1 vccd1 _15531_/A sky130_fd_sc_hd__and2_1
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12742_/A _20639_/D _20639_/C vssd1 vssd1 vccd1 vccd1 _12748_/A sky130_fd_sc_hd__nand3_1
XFILLER_16_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15461_ _15462_/A _15462_/B _15462_/C vssd1 vssd1 vccd1 vccd1 _15467_/B sky130_fd_sc_hd__o21ai_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _23451_/Q vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__inv_2
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18146__A _23530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17200_ _17200_/A _17200_/B _17200_/C vssd1 vssd1 vccd1 vccd1 _17200_/Y sky130_fd_sc_hd__nand3_1
X_11624_ _11624_/A vssd1 vssd1 vccd1 vccd1 _16802_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14412_ _14414_/A _14414_/B vssd1 vssd1 vccd1 vccd1 _14416_/A sky130_fd_sc_hd__nand2_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ _18180_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _18182_/A sky130_fd_sc_hd__nand2_1
XFILLER_175_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15392_ _15392_/A _15392_/B vssd1 vssd1 vccd1 vccd1 _15392_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17131_ _17133_/A _17133_/B vssd1 vssd1 vccd1 vccd1 _17303_/A sky130_fd_sc_hd__nand2_2
XANTENNA__17985__A _20133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16155__A1 _15971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14343_ _14407_/B _14355_/C _14355_/A vssd1 vssd1 vccd1 vccd1 _14403_/C sky130_fd_sc_hd__a21o_1
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17062_ _17761_/B _17062_/B _17761_/A vssd1 vssd1 vccd1 vccd1 _17069_/A sky130_fd_sc_hd__nand3_2
XFILLER_13_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14274_ _15231_/A _14009_/X _14269_/Y _14054_/Y vssd1 vssd1 vccd1 vccd1 _14279_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_156_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13225_ _13732_/B _13732_/C vssd1 vssd1 vccd1 vccd1 _13299_/A sky130_fd_sc_hd__nor2_1
X_16013_ _16004_/X _16005_/Y _16012_/Y vssd1 vssd1 vccd1 vccd1 _16017_/A sky130_fd_sc_hd__o21ai_1
XFILLER_83_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12192__A2 _17642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ _13156_/A vssd1 vssd1 vccd1 vccd1 _21279_/D sky130_fd_sc_hd__buf_2
XFILLER_88_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12107_ _12107_/A vssd1 vssd1 vccd1 vccd1 _12107_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17964_ _17964_/A _23260_/B _17964_/C vssd1 vssd1 vccd1 vccd1 _17964_/Y sky130_fd_sc_hd__nor3_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13087_ _20594_/A _20594_/B _13087_/C vssd1 vssd1 vccd1 vccd1 _13205_/C sky130_fd_sc_hd__nand3_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21954__B _22089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17407__A1 _16684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19703_ _19703_/A _19703_/B _19703_/C _19703_/D vssd1 vssd1 vccd1 vccd1 _19708_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__17407__B2 _11948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16915_ _16669_/A _16669_/B _16662_/B vssd1 vssd1 vccd1 vccd1 _16923_/C sky130_fd_sc_hd__a21o_1
XFILLER_66_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12038_ _15706_/A vssd1 vssd1 vccd1 vccd1 _15682_/A sky130_fd_sc_hd__buf_2
XANTENNA__21203__A2 _21061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17895_ _20217_/D _17969_/D _17754_/Y _17760_/Y vssd1 vssd1 vccd1 vccd1 _17896_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19634_ _19636_/B _19788_/A vssd1 vssd1 vccd1 vccd1 _19635_/B sky130_fd_sc_hd__or2b_1
XANTENNA__17225__A _18506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16846_ _17061_/A vssd1 vssd1 vccd1 vccd1 _18607_/C sky130_fd_sc_hd__buf_2
XFILLER_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19565_ _19555_/Y _19556_/X _19546_/Y _19552_/Y vssd1 vssd1 vccd1 vccd1 _19567_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16777_ _16584_/A _16762_/Y _16776_/Y vssd1 vssd1 vccd1 vccd1 _16777_/Y sky130_fd_sc_hd__a21oi_2
X_13989_ _14360_/A _14791_/B _14806_/C _14911_/B vssd1 vssd1 vccd1 vccd1 _13989_/Y
+ sky130_fd_sc_hd__a22oi_1
X_18516_ _12353_/X _17643_/X _18501_/X _12463_/Y _18520_/A vssd1 vssd1 vccd1 vccd1
+ _18516_/X sky130_fd_sc_hd__o311a_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ _23414_/Q vssd1 vssd1 vccd1 vccd1 _15864_/A sky130_fd_sc_hd__inv_2
X_19496_ _19522_/A _19577_/B _19577_/C vssd1 vssd1 vccd1 vccd1 _19575_/A sky130_fd_sc_hd__a21o_2
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19580__A1 _19207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18447_ _19010_/A _18447_/B _19157_/C vssd1 vssd1 vccd1 vccd1 _18448_/B sky130_fd_sc_hd__nand3_1
XANTENNA__15197__A2 _14777_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15659_ _15659_/A vssd1 vssd1 vccd1 vccd1 _15660_/A sky130_fd_sc_hd__buf_2
XFILLER_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22467__A1 _13495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18378_ _18378_/A _18378_/B _18378_/C vssd1 vssd1 vccd1 vccd1 _18410_/A sky130_fd_sc_hd__and3_1
XFILLER_147_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17329_ _17330_/A _17330_/B _17330_/C vssd1 vssd1 vccd1 vccd1 _17331_/A sky130_fd_sc_hd__a21oi_2
XFILLER_18_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22009__C _22218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_902 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20340_ _19785_/X _20205_/X _20293_/X _20294_/X _20343_/A vssd1 vssd1 vccd1 vccd1
+ _20340_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__22219__A1 _22508_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18503__B _18503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20271_ _20271_/A _20371_/C _20271_/C _20271_/D vssd1 vssd1 vccd1 vccd1 _20271_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_162_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12832__A _20532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22010_ _22064_/A vssd1 vssd1 vccd1 vccd1 _22564_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__17646__A1 _17643_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17646__B2 _20081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15862__B _15862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19334__B _19539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13663__A _13663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22912_ _12712_/X input35/X _22918_/S vssd1 vssd1 vccd1 vccd1 _22913_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20953__A1 _12675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22843_ _22843_/A _22843_/B vssd1 vssd1 vccd1 vccd1 _22849_/A sky130_fd_sc_hd__nand2_2
XANTENNA__12279__A _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_732 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22774_ _22774_/A _22774_/B _22808_/A vssd1 vssd1 vccd1 vccd1 _22774_/X sky130_fd_sc_hd__or3_1
XFILLER_197_512 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21725_ _21723_/Y _21717_/Y _21728_/B vssd1 vssd1 vccd1 vccd1 _21726_/B sky130_fd_sc_hd__o21ai_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11997__A2 _11713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21656_ _21627_/B _21540_/X _21627_/C _21625_/X vssd1 vssd1 vccd1 vccd1 _21656_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14935__A2 _15044_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20607_ _20607_/A _20607_/B _20607_/C vssd1 vssd1 vccd1 vccd1 _20608_/C sky130_fd_sc_hd__nand3_1
X_21587_ _21540_/X _21585_/X _21586_/X vssd1 vssd1 vccd1 vccd1 _23550_/D sky130_fd_sc_hd__a21bo_1
XFILLER_123_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23326_ _23327_/CLK _23326_/D vssd1 vssd1 vccd1 vccd1 _23326_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_193_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16688__A2 _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20538_ _20957_/A _12936_/X _12952_/X _13025_/X vssd1 vssd1 vccd1 vccd1 _20542_/C
+ sky130_fd_sc_hd__o22ai_2
XFILLER_125_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21120__A _21387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23257_ _23257_/A vssd1 vssd1 vccd1 vccd1 _23579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15360__A2 _14184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20469_ _20628_/A vssd1 vssd1 vccd1 vccd1 _21493_/A sky130_fd_sc_hd__buf_2
XFILLER_181_979 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13010_ _23294_/Q _23295_/Q vssd1 vssd1 vccd1 vccd1 _20798_/C sky130_fd_sc_hd__nor2_4
XFILLER_165_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22208_ _22208_/A _22208_/B _22208_/C vssd1 vssd1 vccd1 vccd1 _22208_/X sky130_fd_sc_hd__and3_1
X_23188_ _23188_/A vssd1 vssd1 vccd1 vccd1 _23414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22139_ _22139_/A _22139_/B _22139_/C vssd1 vssd1 vccd1 vccd1 _22215_/B sky130_fd_sc_hd__and3_1
XFILLER_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input36_A wb_dat_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14961_ _14961_/A vssd1 vssd1 vccd1 vccd1 _15289_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_48_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_770 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16700_ _16700_/A vssd1 vssd1 vccd1 vccd1 _16957_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18062__A1 _23528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13912_ _14069_/A vssd1 vssd1 vccd1 vccd1 _14795_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17680_ _17700_/A _17680_/B _17680_/C vssd1 vssd1 vccd1 vccd1 _17686_/A sky130_fd_sc_hd__nand3_2
X_14892_ _15004_/B _14884_/X _14885_/Y _14891_/Y vssd1 vssd1 vccd1 vccd1 _14908_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__12882__B1 _12875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16631_ _16649_/A vssd1 vssd1 vccd1 vccd1 _16853_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13843_ _13843_/A _13843_/B _13843_/C vssd1 vssd1 vccd1 vccd1 _13853_/B sky130_fd_sc_hd__nand3_2
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19260__A _20320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19350_ _19350_/A vssd1 vssd1 vccd1 vccd1 _19735_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16562_ _16562_/A _16562_/B vssd1 vssd1 vccd1 vccd1 _16567_/A sky130_fd_sc_hd__nand2_1
XFILLER_74_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13774_ _13642_/A _13492_/A _13630_/A _13630_/B vssd1 vssd1 vccd1 vccd1 _13774_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_90_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18301_ _18301_/A _18301_/B vssd1 vssd1 vccd1 vccd1 _18314_/C sky130_fd_sc_hd__nand2_1
XFILLER_188_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15513_ _15536_/B _15513_/B _15513_/C _15513_/D vssd1 vssd1 vccd1 vccd1 _15514_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_71_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19281_ _20120_/A _19924_/A _19107_/C _19107_/B vssd1 vssd1 vccd1 vccd1 _19281_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12725_ _12725_/A vssd1 vssd1 vccd1 vccd1 _12725_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16493_ _16356_/X _16384_/X _16458_/X _16478_/X vssd1 vssd1 vccd1 vccd1 _16493_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_188_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12917__A _23456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18232_ _18098_/X _18094_/X _18095_/X _18179_/B vssd1 vssd1 vccd1 vccd1 _18233_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_128_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23584__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11821__A _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15444_ _15430_/B _15430_/A _15431_/A _15431_/B vssd1 vssd1 vccd1 vccd1 _15474_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12656_ _12652_/X _12651_/X _12654_/Y vssd1 vssd1 vccd1 vccd1 _12661_/A sky130_fd_sc_hd__o21ai_1
XFILLER_90_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19314__A1 _11822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18163_ _18163_/A _18163_/B _18163_/C _18163_/D vssd1 vssd1 vccd1 vccd1 _18165_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_175_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ _23397_/Q vssd1 vssd1 vccd1 vccd1 _11608_/A sky130_fd_sc_hd__buf_2
X_15375_ _15375_/A vssd1 vssd1 vccd1 vccd1 _15536_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12587_ _12875_/C vssd1 vssd1 vccd1 vccd1 _14655_/A sky130_fd_sc_hd__buf_2
X_17114_ _17125_/A _17298_/A _17109_/X _17113_/X vssd1 vssd1 vccd1 vccd1 _17120_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_117_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14326_ _14367_/C _14367_/B _14325_/B vssd1 vssd1 vccd1 vccd1 _14365_/B sky130_fd_sc_hd__a21o_1
X_18094_ _18169_/A _18101_/B _18100_/A _18101_/D vssd1 vssd1 vccd1 vccd1 _18094_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_8_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17045_ _16625_/X _17252_/A _19381_/B _17039_/Y _16499_/A vssd1 vssd1 vccd1 vccd1
+ _17047_/B sky130_fd_sc_hd__o2111ai_4
X_14257_ _14796_/A _14276_/A _14790_/C vssd1 vssd1 vccd1 vccd1 _14340_/B sky130_fd_sc_hd__and3_1
XFILLER_125_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17628__A1 _16781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13208_ _13208_/A _13208_/B vssd1 vssd1 vccd1 vccd1 _20465_/D sky130_fd_sc_hd__nand2_1
XANTENNA__13467__B _21925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14188_ _14188_/A _23354_/Q _14188_/C vssd1 vssd1 vccd1 vccd1 _14864_/C sky130_fd_sc_hd__nor3_2
XFILLER_140_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13139_ _13138_/A _13138_/B _13138_/C _13138_/D vssd1 vssd1 vccd1 vccd1 _13140_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_854 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ _18996_/A _18996_/B _18996_/C vssd1 vssd1 vccd1 vccd1 _19163_/A sky130_fd_sc_hd__nand3_4
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16778__B _16792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13114__A1 _21050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13114__B2 _21050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17947_ _17820_/Y _17825_/Y _17946_/X vssd1 vssd1 vccd1 vccd1 _18148_/B sky130_fd_sc_hd__o21ai_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17878_ _17878_/A _17878_/B vssd1 vssd1 vccd1 vccd1 _17878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14298__B _14834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19617_ _19638_/A _19638_/C vssd1 vssd1 vccd1 vccd1 _19617_/Y sky130_fd_sc_hd__nand2_1
X_16829_ _12511_/A _12513_/A _15855_/Y _15856_/Y _17594_/A vssd1 vssd1 vccd1 vccd1
+ _17068_/A sky130_fd_sc_hd__o221ai_4
XFILLER_0_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15811__B1 _15974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19548_ _19548_/A vssd1 vssd1 vccd1 vccd1 _19967_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14090__A2 _14203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19479_ _18476_/A _18484_/A _18503_/B _18503_/A _18479_/A vssd1 vssd1 vccd1 vccd1
+ _19480_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21510_ _21510_/A _21510_/B _21510_/C vssd1 vssd1 vccd1 vccd1 _21510_/X sky130_fd_sc_hd__and3_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22490_ _22493_/B vssd1 vssd1 vccd1 vccd1 _22544_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19305__A1 _11799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21441_ _21359_/B _21635_/C _21314_/A _21433_/Y _21552_/A vssd1 vssd1 vccd1 vccd1
+ _21442_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17316__B1 _17140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18513__C1 _19534_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21372_ _21371_/C _21440_/B _21371_/B _21546_/A _21448_/B vssd1 vssd1 vccd1 vccd1
+ _21372_/X sky130_fd_sc_hd__a32o_1
XFILLER_107_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_795 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15878__B1 _15866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23111_ _23111_/A vssd1 vssd1 vccd1 vccd1 _23381_/D sky130_fd_sc_hd__clkbuf_1
X_20323_ _20400_/A _20400_/B _20323_/C vssd1 vssd1 vccd1 vccd1 _20325_/A sky130_fd_sc_hd__and3_1
XANTENNA__13658__A _13660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23042_ _23110_/S vssd1 vssd1 vccd1 vccd1 _23051_/S sky130_fd_sc_hd__clkbuf_2
X_20254_ _20118_/X _20307_/A _20252_/X _20253_/Y vssd1 vssd1 vccd1 vccd1 _20255_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__13377__B _13377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15873__A _19700_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20185_ _20185_/A _20185_/B vssd1 vssd1 vccd1 vccd1 _20186_/B sky130_fd_sc_hd__nor2_1
XFILLER_153_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16842__A2 _15972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20139__C1 _17414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22826_ _22824_/Y _22854_/B vssd1 vssd1 vccd1 vccd1 _22827_/A sky130_fd_sc_hd__and2b_1
XFILLER_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16358__A1 _12379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22757_ _22830_/A _22757_/B _22830_/D vssd1 vssd1 vccd1 vccd1 _22759_/A sky130_fd_sc_hd__or3_1
XFILLER_73_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12510_ _12510_/A _17964_/A vssd1 vssd1 vccd1 vccd1 _12511_/A sky130_fd_sc_hd__nor2_2
XFILLER_73_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21708_ _21616_/X _21617_/X _21705_/X vssd1 vssd1 vccd1 vccd1 _21721_/B sky130_fd_sc_hd__o21a_1
X_13490_ _13490_/A _13490_/B vssd1 vssd1 vccd1 vccd1 _13494_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22688_ _21854_/A _21854_/B _22630_/X _22687_/Y vssd1 vssd1 vccd1 vccd1 _22690_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_60_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ _12441_/A _12441_/B vssd1 vssd1 vccd1 vccd1 _12443_/B sky130_fd_sc_hd__nand2_1
X_21639_ _21635_/X _21695_/A _21638_/X vssd1 vssd1 vccd1 vccd1 _21641_/C sky130_fd_sc_hd__a21boi_1
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18646__A1_N _19196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12372_ _12372_/A _12372_/B _12372_/C _12372_/D vssd1 vssd1 vccd1 vccd1 _12384_/B
+ sky130_fd_sc_hd__nand4_1
X_15160_ _15085_/X _15082_/Y _15083_/X vssd1 vssd1 vccd1 vccd1 _15228_/B sky130_fd_sc_hd__a21boi_2
XFILLER_153_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14111_ _23496_/Q vssd1 vssd1 vccd1 vccd1 _14276_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_23309_ _23309_/CLK _23309_/D vssd1 vssd1 vccd1 vccd1 _23309_/Q sky130_fd_sc_hd__dfxtp_1
X_15091_ _14979_/X _15089_/X _15090_/Y vssd1 vssd1 vccd1 vccd1 _15092_/B sky130_fd_sc_hd__o21ai_1
XFILLER_126_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14042_ _23496_/Q vssd1 vssd1 vccd1 vccd1 _14183_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18850_ _19123_/C _18958_/B _18856_/A _19334_/A vssd1 vssd1 vccd1 vccd1 _18852_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_192_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17801_ _17709_/Y _17801_/B _17801_/C vssd1 vssd1 vccd1 vccd1 _17805_/A sky130_fd_sc_hd__nand3b_2
XFILLER_67_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18781_ _19073_/A _18781_/B _18882_/A vssd1 vssd1 vccd1 vccd1 _18889_/B sky130_fd_sc_hd__and3_2
X_15993_ _15993_/A _17235_/A _17450_/C vssd1 vssd1 vccd1 vccd1 _15993_/X sky130_fd_sc_hd__and3_1
X_17732_ _17781_/B vssd1 vssd1 vccd1 vccd1 _17838_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14944_ _14944_/A _14944_/B vssd1 vssd1 vccd1 vccd1 _14945_/C sky130_fd_sc_hd__xor2_1
XFILLER_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12855__B1 _21035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_84 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17663_ _17663_/A _17663_/B vssd1 vssd1 vccd1 vccd1 _17663_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16924__A2_N _16930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22119__B1 _21995_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14875_ _14058_/X _14904_/A _15120_/B _14872_/Y _15155_/A vssd1 vssd1 vccd1 vccd1
+ _14899_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__17794__B1 _17792_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19402_ _19402_/A _19402_/B vssd1 vssd1 vccd1 vccd1 _19402_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16614_ _16614_/A _16828_/A vssd1 vssd1 vccd1 vccd1 _16614_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13826_ _13456_/A _13456_/B _13642_/A vssd1 vssd1 vccd1 vccd1 _13826_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17594_ _17594_/A vssd1 vssd1 vccd1 vccd1 _17595_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__19535__A1 _18435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19333_ _11926_/X _19803_/A _19196_/C _19482_/A _19328_/Y vssd1 vssd1 vccd1 vccd1
+ _19333_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16545_ _16531_/A _16543_/X _16544_/Y vssd1 vssd1 vccd1 vccd1 _16545_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ _13755_/Y _13698_/A _13525_/C _13756_/Y vssd1 vssd1 vccd1 vccd1 _13757_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16119__A _16119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19264_ _19297_/A _19297_/B _19261_/X _19263_/X vssd1 vssd1 vccd1 vccd1 _19275_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_12708_ _13138_/A _13138_/B vssd1 vssd1 vccd1 vccd1 _12923_/C sky130_fd_sc_hd__nand2_1
X_16476_ _16517_/B _16476_/B _16476_/C _16476_/D vssd1 vssd1 vccd1 vccd1 _16477_/C
+ sky130_fd_sc_hd__nand4_1
X_13688_ _22220_/C vssd1 vssd1 vccd1 vccd1 _22508_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__15021__A1 _15019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18215_ _19967_/C vssd1 vssd1 vccd1 vccd1 _20212_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_148_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15427_ _15427_/A _15451_/B vssd1 vssd1 vccd1 vccd1 _15463_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__23095__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19195_ _19195_/A vssd1 vssd1 vccd1 vccd1 _19196_/C sky130_fd_sc_hd__buf_2
X_12639_ _12683_/B _12712_/A vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__nand2_2
XFILLER_157_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14375__A3 _15195_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20583__B _21387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18146_ _23530_/Q vssd1 vssd1 vccd1 vccd1 _18146_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17849__A1 _17742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15358_ _15358_/A _15416_/A vssd1 vssd1 vccd1 vccd1 _15358_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14309_ _14310_/A _14842_/A _14309_/C vssd1 vssd1 vccd1 vccd1 _14846_/B sky130_fd_sc_hd__nand3b_1
X_18077_ _18077_/A vssd1 vssd1 vccd1 vccd1 _20217_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15289_ _15402_/A _15402_/B _15289_/C vssd1 vssd1 vccd1 vccd1 _15291_/A sky130_fd_sc_hd__and3_1
XFILLER_85_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17028_ _16964_/A _16964_/B _16964_/C _16969_/C vssd1 vssd1 vccd1 vccd1 _17028_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18274__A1 _18330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19165__A _19502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18274__B2 _18276_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _18813_/A _18996_/B _18818_/A vssd1 vssd1 vccd1 vccd1 _18980_/A sky130_fd_sc_hd__o21ai_2
XFILLER_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21990_ _22236_/A vssd1 vssd1 vccd1 vccd1 _22090_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20941_ _20941_/A _20941_/B vssd1 vssd1 vccd1 vccd1 _20941_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16588__A1 _12222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13941__A _23499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20872_ _20872_/A _20872_/B _20872_/C vssd1 vssd1 vccd1 vccd1 _21157_/D sky130_fd_sc_hd__nand3_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22611_ _22611_/A _22611_/B vssd1 vssd1 vccd1 vccd1 _22611_/X sky130_fd_sc_hd__or2_1
X_23591_ _23598_/CLK _23591_/D vssd1 vssd1 vccd1 vccd1 _23591_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__16674__D _17098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17001__A2 _17218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22542_ _22513_/A _22513_/C _22541_/X vssd1 vssd1 vccd1 vccd1 _22594_/A sky130_fd_sc_hd__a21oi_1
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22473_ _22473_/A _22473_/B vssd1 vssd1 vccd1 vccd1 _22501_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21424_ _21424_/A _21424_/B vssd1 vssd1 vccd1 vccd1 _21424_/X sky130_fd_sc_hd__or2_1
XANTENNA__12377__A2 _11931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22833__A1 _22830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18501__A2 _11760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21355_ _21330_/A _21330_/B _21330_/C _21331_/B _21266_/X vssd1 vssd1 vccd1 vccd1
+ _21476_/A sky130_fd_sc_hd__a32o_2
XFILLER_108_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20306_ _20306_/A vssd1 vssd1 vccd1 vccd1 _20452_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21286_ _21278_/X _21280_/Y _21285_/Y vssd1 vssd1 vccd1 vccd1 _21380_/A sky130_fd_sc_hd__o21ai_2
XFILLER_162_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23025_ _23025_/A vssd1 vssd1 vccd1 vccd1 _23034_/S sky130_fd_sc_hd__clkbuf_2
X_20237_ _20176_/C _20179_/X _20234_/Y _20235_/X vssd1 vssd1 vccd1 vccd1 _20237_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_103_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11888__A1 _11760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20168_ _20229_/A _20229_/B _20229_/C vssd1 vssd1 vccd1 vccd1 _20171_/B sky130_fd_sc_hd__nand3_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23010__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15108__A _15120_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19803__A _19803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20099_ _20097_/Y _20099_/B _20177_/A vssd1 vssd1 vccd1 vccd1 _20177_/B sky130_fd_sc_hd__nand3b_2
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _12904_/A _12991_/B _12991_/C vssd1 vssd1 vccd1 vccd1 _20584_/A sky130_fd_sc_hd__a21o_1
XFILLER_188_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _16591_/B vssd1 vssd1 vccd1 vccd1 _18503_/B sky130_fd_sc_hd__buf_4
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17323__A _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _18434_/A _14640_/X _14647_/X _16780_/B _14659_/X vssd1 vssd1 vccd1 vccd1
+ _14660_/X sky130_fd_sc_hd__a221o_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11887_/C vssd1 vssd1 vccd1 vccd1 _18503_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_189_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _13616_/A _13615_/A _13609_/X _13610_/Y vssd1 vssd1 vccd1 vccd1 _13627_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_26_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22809_ _22810_/A _22810_/B _22808_/Y vssd1 vssd1 vccd1 vccd1 _22812_/A sky130_fd_sc_hd__o21ai_4
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13262__B1 _23322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14591_ _12113_/X _14544_/X _14585_/X _14590_/X vssd1 vssd1 vccd1 vccd1 _14591_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12467__A _16122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ _16396_/B _16397_/B _16324_/Y vssd1 vssd1 vccd1 vccd1 _16330_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_198_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13542_ _13477_/X _13598_/A _13538_/X vssd1 vssd1 vccd1 vccd1 _13542_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11812__A1 _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15003__A1 _14181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16261_ _16248_/A _16248_/B _16248_/C _16248_/D vssd1 vssd1 vccd1 vccd1 _16261_/Y
+ sky130_fd_sc_hd__a22oi_2
X_13473_ _13468_/X _13472_/X _13460_/D _13460_/A vssd1 vssd1 vccd1 vccd1 _13476_/B
+ sky130_fd_sc_hd__o211ai_1
X_18000_ _18000_/A vssd1 vssd1 vccd1 vccd1 _20081_/B sky130_fd_sc_hd__buf_2
X_15212_ _15212_/A _15211_/Y vssd1 vssd1 vccd1 vccd1 _15214_/A sky130_fd_sc_hd__nor2b_2
X_12424_ _12424_/A vssd1 vssd1 vccd1 vccd1 _19190_/A sky130_fd_sc_hd__buf_4
X_16192_ _16671_/A _16671_/B _16225_/A vssd1 vssd1 vccd1 vccd1 _16192_/X sky130_fd_sc_hd__a21o_1
XANTENNA__19296__A3 _19261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15928__D _17753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15143_ _15144_/B _15144_/A vssd1 vssd1 vccd1 vccd1 _15286_/A sky130_fd_sc_hd__nand2_2
XANTENNA__16503__A1 _15855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ _12355_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12355_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19951_ _20371_/C _19951_/B _19951_/C _19951_/D vssd1 vssd1 vccd1 vccd1 _19952_/A
+ sky130_fd_sc_hd__nand4_1
X_12286_ _12297_/B _12297_/C _12280_/Y _12285_/X vssd1 vssd1 vccd1 vccd1 _12288_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15074_ _15050_/A _15050_/C _15050_/B vssd1 vssd1 vccd1 vccd1 _15074_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_135_990 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18902_ _18902_/A _18902_/B vssd1 vssd1 vccd1 vccd1 _18903_/B sky130_fd_sc_hd__nand2_1
X_14025_ _14075_/A _14262_/A _14035_/A vssd1 vssd1 vccd1 vccd1 _14054_/A sky130_fd_sc_hd__nand3_1
XFILLER_49_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19882_ _19831_/A _19831_/B _19831_/C _19723_/B _19723_/C vssd1 vssd1 vccd1 vccd1
+ _19882_/X sky130_fd_sc_hd__a32o_1
XFILLER_136_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18833_ _18669_/A _18669_/B _18831_/Y _18832_/X vssd1 vssd1 vccd1 vccd1 _18833_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_67_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18008__A1 _18016_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18764_ _12378_/A _12378_/B _17761_/A _17761_/B vssd1 vssd1 vccd1 vccd1 _18765_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__23001__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15976_ _11935_/A _15972_/X _15843_/B _16123_/A _16172_/A vssd1 vssd1 vccd1 vccd1
+ _15976_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_83_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17715_ _17628_/Y _17712_/Y _17899_/A _19957_/D _17899_/B vssd1 vssd1 vccd1 vccd1
+ _17715_/Y sky130_fd_sc_hd__o2111ai_4
X_14927_ _14966_/A _14927_/B _14927_/C _14927_/D vssd1 vssd1 vccd1 vccd1 _14966_/B
+ sky130_fd_sc_hd__nand4_2
X_18695_ _18673_/X _17643_/A _18674_/X _18675_/X vssd1 vssd1 vccd1 vccd1 _18753_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17646_ _17643_/X _17644_/X _17752_/A _20081_/A vssd1 vssd1 vccd1 vccd1 _17646_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17231__A2 _12237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17233__A _17233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16034__A3 _18434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14858_ _14858_/A vssd1 vssd1 vccd1 vccd1 _15155_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13809_ _13809_/A _13809_/B vssd1 vssd1 vccd1 vccd1 _22014_/A sky130_fd_sc_hd__nand2_2
XFILLER_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17577_ _17566_/X _17575_/X _20133_/D _17571_/Y _17845_/D vssd1 vssd1 vccd1 vccd1
+ _17578_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_91_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789_ _14789_/A _14857_/B _14789_/C vssd1 vssd1 vccd1 vccd1 _14814_/B sky130_fd_sc_hd__nand3_2
XFILLER_56_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19316_ _19320_/A _19321_/A _19517_/B vssd1 vssd1 vccd1 vccd1 _19316_/Y sky130_fd_sc_hd__a21oi_1
X_16528_ _16528_/A _16528_/B _16536_/B _16544_/A vssd1 vssd1 vccd1 vccd1 _16544_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_50_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21866__A2 _21971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19247_ _18968_/A _19246_/Y _18969_/D vssd1 vssd1 vccd1 vccd1 _19254_/A sky130_fd_sc_hd__o21a_1
XFILLER_177_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16459_ _16457_/A _16457_/B _16356_/A _16458_/X vssd1 vssd1 vccd1 vccd1 _16459_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_177_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12359__A2 _19534_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_838 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19178_ _19325_/A _19183_/B _19178_/C vssd1 vssd1 vccd1 vccd1 _19178_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__12213__D1 _18952_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18129_ _18129_/A _18129_/B vssd1 vssd1 vccd1 vccd1 _18129_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21140_ _21241_/A _21243_/B _21140_/C vssd1 vssd1 vccd1 vccd1 _21344_/B sky130_fd_sc_hd__nand3_1
XFILLER_117_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12262__D _18531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17408__A _17642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21071_ _21365_/A _21276_/A vssd1 vssd1 vccd1 vccd1 _21071_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20022_ _20184_/A _20184_/B _20185_/A vssd1 vssd1 vccd1 vccd1 _20113_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22968__B input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21973_ _22107_/B _22107_/C _21973_/C _21980_/A vssd1 vssd1 vccd1 vccd1 _21976_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20924_ _21036_/B vssd1 vssd1 vccd1 vccd1 _21282_/A sky130_fd_sc_hd__clkbuf_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _20772_/X _20770_/X _20776_/A _20847_/B _20847_/A vssd1 vssd1 vccd1 vccd1
+ _20856_/C sky130_fd_sc_hd__o2111ai_1
XANTENNA__11903__B _11912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12287__A _12297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22503__B1 _21829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23574_ _23575_/CLK _23574_/D vssd1 vssd1 vccd1 vccd1 _23574_/Q sky130_fd_sc_hd__dfxtp_1
X_20786_ _20921_/A _20921_/B vssd1 vssd1 vccd1 vccd1 _20786_/Y sky130_fd_sc_hd__nand2_2
XFILLER_70_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20935__C _21050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22525_ _22523_/Y _22525_/B vssd1 vssd1 vccd1 vccd1 _22729_/B sky130_fd_sc_hd__nand2b_1
XFILLER_167_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14744__B1 _14738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22456_ _22443_/A _22443_/B _22445_/Y vssd1 vssd1 vccd1 vccd1 _22629_/A sky130_fd_sc_hd__a21oi_2
XFILLER_183_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21407_ _21407_/A _21407_/B vssd1 vssd1 vccd1 vccd1 _21411_/B sky130_fd_sc_hd__nor2_1
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22387_ _22283_/X _22567_/A _13527_/X _22641_/B _22386_/Y vssd1 vssd1 vccd1 vccd1
+ _22463_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_135_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20951__B _20984_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20293__A1 _20290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ _12491_/A _12491_/B _12139_/Y vssd1 vssd1 vccd1 vccd1 _12157_/A sky130_fd_sc_hd__o21ai_1
XFILLER_159_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21338_ _21012_/A _21251_/Y _21154_/Y vssd1 vssd1 vccd1 vccd1 _21404_/A sky130_fd_sc_hd__o21ai_2
XFILLER_135_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12071_ _12071_/A vssd1 vssd1 vccd1 vccd1 _15957_/C sky130_fd_sc_hd__buf_2
XANTENNA__19435__B1 _19431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21269_ _21270_/A _21270_/B _21270_/C vssd1 vssd1 vccd1 vccd1 _21273_/A sky130_fd_sc_hd__a21o_1
XFILLER_104_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23231__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23008_ _23335_/Q input15/X _23012_/S vssd1 vssd1 vccd1 vccd1 _23009_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22990__A0 _13603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22878__B _22878_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _12147_/X _12146_/X _18481_/B _12149_/X _18481_/C vssd1 vssd1 vccd1 vccd1
+ _15830_/X sky130_fd_sc_hd__o2111a_1
XANTENNA__17461__A2 _17465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13284__C _22280_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22337__A3 _22226_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15761_ _15761_/A vssd1 vssd1 vccd1 vccd1 _15761_/X sky130_fd_sc_hd__buf_2
X_12973_ _12962_/A _12962_/B _12962_/C vssd1 vssd1 vccd1 vccd1 _12973_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14677__A _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _17327_/B _17327_/C _17327_/A _17330_/A _17499_/X vssd1 vssd1 vccd1 vccd1
+ _17502_/C sky130_fd_sc_hd__a32o_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _23347_/Q _14531_/A _14546_/A _23315_/Q _14699_/X vssd1 vssd1 vccd1 vccd1
+ _14712_/X sky130_fd_sc_hd__a221o_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _18474_/X _20320_/B _19846_/A _19180_/C vssd1 vssd1 vccd1 vccd1 _18480_/Y
+ sky130_fd_sc_hd__nand4b_2
X_11924_ _11924_/A vssd1 vssd1 vccd1 vccd1 _17626_/A sky130_fd_sc_hd__buf_2
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15692_ _23419_/Q vssd1 vssd1 vccd1 vccd1 _15692_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22894__A _22895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17431_ _17431_/A vssd1 vssd1 vccd1 vccd1 _17733_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _22142_/B _14636_/X _14642_/X _23300_/Q _14587_/X vssd1 vssd1 vccd1 vccd1
+ _14643_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _16365_/A vssd1 vssd1 vccd1 vccd1 _18481_/C sky130_fd_sc_hd__buf_2
XFILLER_82_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16972__A1 _16724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17362_ _17362_/A _17362_/B _17362_/C vssd1 vssd1 vccd1 vccd1 _17362_/Y sky130_fd_sc_hd__nand3_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14574_ _23184_/D vssd1 vssd1 vccd1 vccd1 _14647_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11786_ _18812_/A _12100_/C _11977_/B vssd1 vssd1 vccd1 vccd1 _12145_/B sky130_fd_sc_hd__a21o_2
X_19101_ _23543_/Q _19101_/B _19101_/C vssd1 vssd1 vccd1 vccd1 _19289_/B sky130_fd_sc_hd__nand3b_1
XFILLER_198_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16313_ _16313_/A _16313_/B _16313_/C vssd1 vssd1 vccd1 vccd1 _16396_/B sky130_fd_sc_hd__nand3_2
X_13525_ _13547_/A _21815_/B _13525_/C _21815_/C vssd1 vssd1 vccd1 vccd1 _13544_/A
+ sky130_fd_sc_hd__or4_2
X_17293_ _17221_/X _17222_/Y _17289_/Y _17292_/Y vssd1 vssd1 vccd1 vccd1 _17337_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_41_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15442__A_N _15439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12925__A _21050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20520__A2 _20509_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15939__C _16281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19032_ _18854_/X _19031_/X _18958_/C vssd1 vssd1 vccd1 vccd1 _19138_/B sky130_fd_sc_hd__o21ai_2
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15301__A _15301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16244_ _16254_/A _16254_/B _16239_/Y _16243_/Y vssd1 vssd1 vccd1 vccd1 _16248_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_13456_ _13456_/A _13456_/B vssd1 vssd1 vccd1 vccd1 _21877_/A sky130_fd_sc_hd__nand2_2
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18477__A1 _12410_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12407_ _18470_/C _18810_/A vssd1 vssd1 vccd1 vccd1 _18440_/A sky130_fd_sc_hd__nand2_2
XFILLER_173_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16175_ _16175_/A _16175_/B _16175_/C vssd1 vssd1 vccd1 vccd1 _16179_/B sky130_fd_sc_hd__nand3_2
X_13387_ _13433_/A _13433_/B _13434_/B vssd1 vssd1 vccd1 vccd1 _13414_/A sky130_fd_sc_hd__a21o_1
XFILLER_126_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15126_ _15127_/C _15188_/B _15127_/A vssd1 vssd1 vccd1 vccd1 _15130_/B sky130_fd_sc_hd__a21o_1
XFILLER_154_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338_ _12360_/A _12360_/B _12381_/C _12381_/B _12330_/X vssd1 vssd1 vccd1 vccd1
+ _12338_/Y sky130_fd_sc_hd__a41oi_1
XFILLER_126_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22134__A _22521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19934_ _19909_/B _19909_/C _19909_/A vssd1 vssd1 vccd1 vccd1 _19934_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__23222__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15057_ _15064_/A _15064_/B vssd1 vssd1 vccd1 vccd1 _15067_/B sky130_fd_sc_hd__nand2_1
X_12269_ _12281_/A _16523_/A _16523_/B _12093_/X vssd1 vssd1 vccd1 vccd1 _12271_/D
+ sky130_fd_sc_hd__o31ai_1
XANTENNA__15674__C _15674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__A _20966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14008_ _23496_/Q vssd1 vssd1 vccd1 vccd1 _14135_/A sky130_fd_sc_hd__inv_2
XFILLER_141_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19865_ _19873_/B _19873_/C vssd1 vssd1 vccd1 vccd1 _19867_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18816_ _23395_/Q vssd1 vssd1 vccd1 vccd1 _18998_/D sky130_fd_sc_hd__inv_2
XFILLER_96_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19796_ _19796_/A _19796_/B vssd1 vssd1 vccd1 vccd1 _19796_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16660__B1 _17722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18747_ _18747_/A _18747_/B vssd1 vssd1 vccd1 vccd1 _19288_/B sky130_fd_sc_hd__nand2_1
X_15959_ _23594_/Q vssd1 vssd1 vccd1 vccd1 _16141_/D sky130_fd_sc_hd__inv_2
XFILLER_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_955 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18678_ _18859_/A _18859_/B _18859_/C _18859_/D vssd1 vssd1 vccd1 vccd1 _18678_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_52_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17629_ _18000_/A _17230_/A _17628_/Y vssd1 vssd1 vccd1 vccd1 _17629_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_24_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20640_ _20479_/X _20639_/Y _20495_/C vssd1 vssd1 vccd1 vccd1 _20660_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__19901__A1 _19903_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21213__A _21217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20571_ _20769_/A _13176_/C _13176_/A _20562_/B vssd1 vssd1 vccd1 vccd1 _20571_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22028__B _22028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22310_ _22025_/Y _22309_/Y _22166_/C _22166_/A vssd1 vssd1 vccd1 vccd1 _22310_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_23290_ _23295_/CLK _23290_/D vssd1 vssd1 vccd1 vccd1 _23290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19114__C1 _17567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22241_ _22242_/B _22242_/C _22242_/A vssd1 vssd1 vccd1 vccd1 _22439_/C sky130_fd_sc_hd__a21o_1
XFILLER_180_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22172_ _22391_/A _22392_/B _22172_/C vssd1 vssd1 vccd1 vccd1 _22279_/A sky130_fd_sc_hd__nand3_4
XFILLER_160_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21123_ _21236_/A _21134_/B _21123_/C vssd1 vssd1 vccd1 vccd1 _21123_/X sky130_fd_sc_hd__and3_1
XANTENNA__23213__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21054_ _21169_/A _21054_/B _21054_/C _21054_/D vssd1 vssd1 vccd1 vccd1 _21202_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_154_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20005_ _20011_/A _20011_/B vssd1 vssd1 vccd1 vccd1 _20007_/A sky130_fd_sc_hd__nand2_1
XFILLER_115_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18928__C1 _19082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21956_ _21956_/A _21982_/A vssd1 vssd1 vccd1 vccd1 _21957_/C sky130_fd_sc_hd__nand2_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18943__A2 _18604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _20907_/A vssd1 vssd1 vccd1 vccd1 _20907_/X sky130_fd_sc_hd__buf_2
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21887_ _21791_/Y _21881_/Y _22365_/C _21884_/Y _13650_/A vssd1 vssd1 vccd1 vccd1
+ _21984_/D sky130_fd_sc_hd__o2111ai_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _16604_/A vssd1 vssd1 vccd1 vccd1 _19196_/A sky130_fd_sc_hd__buf_2
XANTENNA__17601__A _17761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ _20843_/B _20842_/A _20842_/B vssd1 vssd1 vccd1 vccd1 _20839_/C sky130_fd_sc_hd__nand3_1
XFILLER_74_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23557_ _23578_/CLK _23557_/D vssd1 vssd1 vccd1 vccd1 _23557_/Q sky130_fd_sc_hd__dfxtp_1
X_11571_ _23587_/Q _23588_/Q vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__nor2_1
XFILLER_74_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20769_ _20769_/A _21124_/B vssd1 vssd1 vccd1 vccd1 _20769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20502__A2 _20481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18171__A3 _17959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _13318_/A vssd1 vssd1 vccd1 vccd1 _21882_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22508_ _22508_/A _22508_/B _22508_/C vssd1 vssd1 vccd1 vccd1 _22509_/C sky130_fd_sc_hd__and3_1
XFILLER_182_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14290_ _14290_/A _14290_/B _14290_/C vssd1 vssd1 vccd1 vccd1 _14358_/B sky130_fd_sc_hd__nand3_2
XFILLER_167_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23488_ _23492_/CLK _23500_/Q vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13241_ _13241_/A vssd1 vssd1 vccd1 vccd1 _13520_/A sky130_fd_sc_hd__clkbuf_2
X_22439_ _22439_/A _22439_/B _22439_/C _22439_/D vssd1 vssd1 vccd1 vccd1 _22439_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18459__B2 _12441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20681__B _21431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19120__A2 _12509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12183__C _19539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20266__B2 _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13172_ _13172_/A _13172_/B _13172_/C vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__and3_1
XFILLER_184_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12123_ _12117_/Y _12119_/Y _12122_/Y vssd1 vssd1 vccd1 vccd1 _12123_/Y sky130_fd_sc_hd__a21boi_1
X_17980_ _17980_/A vssd1 vssd1 vccd1 vccd1 _20210_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__22007__A2 _21892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23204__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22889__A _22895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_800 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16931_ _16066_/C _16377_/X _16605_/X _16647_/C _16121_/Y vssd1 vssd1 vccd1 vccd1
+ _16931_/X sky130_fd_sc_hd__o311a_1
X_12054_ _12311_/A _12053_/X _12029_/A vssd1 vssd1 vccd1 vccd1 _12054_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19263__A _19263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19650_ _12323_/A _20080_/A _19656_/B _19649_/Y vssd1 vssd1 vccd1 vccd1 _19650_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_133_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16862_ _16858_/A _16860_/Y _16861_/X vssd1 vssd1 vccd1 vccd1 _16879_/C sky130_fd_sc_hd__a21o_1
XFILLER_78_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18601_ _18601_/A vssd1 vssd1 vccd1 vccd1 _18932_/A sky130_fd_sc_hd__clkbuf_2
X_15813_ _15813_/A _15813_/B vssd1 vssd1 vccd1 vccd1 _15834_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19581_ _19345_/A _19345_/B _19339_/C vssd1 vssd1 vccd1 vccd1 _19581_/X sky130_fd_sc_hd__a21o_1
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16793_ _14736_/X _16796_/A _16807_/B vssd1 vssd1 vccd1 vccd1 _16794_/B sky130_fd_sc_hd__a21oi_4
XFILLER_19_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18532_ _19543_/B _19123_/B _19262_/A _18945_/C vssd1 vssd1 vccd1 vccd1 _18532_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15744_ _15766_/A vssd1 vssd1 vccd1 vccd1 _16447_/B sky130_fd_sc_hd__clkbuf_4
X_12956_ _21054_/B vssd1 vssd1 vccd1 vccd1 _21276_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18934__A2 _12247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _11969_/B _11907_/B vssd1 vssd1 vccd1 vccd1 _11908_/B sky130_fd_sc_hd__or2_1
X_18463_ _12052_/A _18443_/A _18453_/X _18452_/A _18634_/A vssd1 vssd1 vccd1 vccd1
+ _18464_/C sky130_fd_sc_hd__o221ai_4
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _15674_/C _15648_/A _15814_/A _15599_/X vssd1 vssd1 vccd1 vccd1 _16030_/A
+ sky130_fd_sc_hd__o211ai_2
X_12887_ _12899_/B _12899_/C _12887_/C vssd1 vssd1 vccd1 vccd1 _12887_/X sky130_fd_sc_hd__and3_1
XANTENNA__18607__A _18607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17414_ _17414_/A _17414_/B _17414_/C _17414_/D vssd1 vssd1 vccd1 vccd1 _17414_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__12358__C _16549_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14621_/X _14545_/X _14640_/A _14625_/X vssd1 vssd1 vccd1 vccd1 _14626_/X
+ sky130_fd_sc_hd__a211o_1
X_18394_ _18394_/A _18394_/B _18417_/D vssd1 vssd1 vccd1 vccd1 _18395_/B sky130_fd_sc_hd__nand3_1
X_11838_ _11838_/A vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17345_/A vssd1 vssd1 vccd1 vccd1 _17346_/B sky130_fd_sc_hd__inv_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _13977_/B _14545_/X _14547_/X _12667_/B vssd1 vssd1 vccd1 vccd1 _14557_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12431__A1 _12052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ _15928_/C vssd1 vssd1 vccd1 vccd1 _16049_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_140_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16127__A _17712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15669__C _17766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18162__A3 _17723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ _13732_/A _13553_/A _13490_/A vssd1 vssd1 vccd1 vccd1 _13511_/B sky130_fd_sc_hd__o21ai_1
XFILLER_159_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17276_ _17276_/A _17276_/B vssd1 vssd1 vccd1 vccd1 _17276_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14488_ _14474_/Y _14478_/X _14483_/Y _14487_/Y vssd1 vssd1 vccd1 vccd1 _14488_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19015_ _19043_/A _19044_/A _19045_/A _19045_/B vssd1 vssd1 vccd1 vccd1 _19148_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_146_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16227_ _16225_/X _17142_/A _16183_/X _16194_/Y vssd1 vssd1 vccd1 vccd1 _16227_/X
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_3_7_0_bq_clk_i clkbuf_3_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_bq_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_162_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13439_ _21882_/A _13600_/C _21882_/C vssd1 vssd1 vccd1 vccd1 _13440_/B sky130_fd_sc_hd__nand3_1
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16158_ _16066_/A _17565_/A _16154_/Y _16157_/Y vssd1 vssd1 vccd1 vccd1 _16170_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_138_1012 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19157__B _20369_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17122__B2 _17112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__B1 _18503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15109_ _15253_/C vssd1 vssd1 vccd1 vccd1 _15109_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16089_ _16089_/A _16089_/B _16089_/C vssd1 vssd1 vccd1 vccd1 _16089_/X sky130_fd_sc_hd__and3_2
XFILLER_170_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19917_ _19925_/A _19925_/B _20032_/B _19793_/A vssd1 vssd1 vccd1 vccd1 _19919_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22014__D _22381_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17108__D _17259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19848_ _19848_/A _19848_/B vssd1 vssd1 vccd1 vccd1 _19848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19779_ _19768_/Y _19640_/Y _19775_/Y vssd1 vssd1 vccd1 vccd1 _19916_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__15987__A2 _15969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1022 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21810_ _21803_/Y _21806_/X _21809_/Y vssd1 vssd1 vccd1 vccd1 _21810_/Y sky130_fd_sc_hd__a21oi_1
X_22790_ _22790_/A vssd1 vssd1 vccd1 vccd1 _22861_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__22182__A1 _22560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21741_ _22033_/A _22034_/A _21905_/B vssd1 vssd1 vccd1 vccd1 _21896_/A sky130_fd_sc_hd__nand3_2
XFILLER_149_1163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15739__A2 _15862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21672_ _21672_/A _21695_/B vssd1 vssd1 vccd1 vccd1 _21673_/A sky130_fd_sc_hd__or2_1
XFILLER_40_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23411_ _23443_/CLK _23411_/D vssd1 vssd1 vccd1 vccd1 _23411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18689__A1 _18673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17140__B _17140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20623_ _20619_/Y _20793_/A _20632_/B vssd1 vssd1 vccd1 vccd1 _20624_/A sky130_fd_sc_hd__a21oi_1
XFILLER_177_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20554_ _20516_/A _20524_/A _20552_/Y _20553_/X vssd1 vssd1 vccd1 vccd1 _20578_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_23342_ _23345_/CLK _23342_/D vssd1 vssd1 vccd1 vccd1 _23342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15876__A _19700_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20485_ _20628_/A _20628_/B _23448_/Q vssd1 vssd1 vccd1 vccd1 _20485_/Y sky130_fd_sc_hd__nand3_1
X_23273_ _23492_/CLK _23273_/D vssd1 vssd1 vccd1 vccd1 _23273_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12186__B1 _16674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22224_ _21988_/A _22226_/B _21988_/B _22670_/D _22223_/X vssd1 vssd1 vccd1 vccd1
+ _22225_/C sky130_fd_sc_hd__a41oi_4
XFILLER_156_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22155_ _22388_/C _22160_/B vssd1 vssd1 vccd1 vccd1 _22155_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__23198__A0 _15674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15675__A1 _15674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21106_ _21106_/A _21106_/B vssd1 vssd1 vccd1 vccd1 _21115_/B sky130_fd_sc_hd__nand2_1
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22086_ _22086_/A _22086_/B vssd1 vssd1 vccd1 vccd1 _22086_/Y sky130_fd_sc_hd__nor2_1
XFILLER_154_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18613__A1 _12260_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21037_ _21037_/A _21279_/C vssd1 vssd1 vccd1 vccd1 _21184_/A sky130_fd_sc_hd__nand2_2
XFILLER_102_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18613__B2 _12475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16500__A _16526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19169__A2 _19838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11644__A _23586_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ _12810_/A _12810_/B vssd1 vssd1 vccd1 vccd1 _12810_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__19811__A _19811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13790_ _22064_/A _22064_/B _22024_/C vssd1 vssd1 vccd1 vccd1 _13791_/A sky130_fd_sc_hd__nand3_2
X_22988_ _13802_/B input37/X _22990_/S vssd1 vssd1 vccd1 vccd1 _22989_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20957__A _20957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _23293_/Q vssd1 vssd1 vccd1 vccd1 _20639_/C sky130_fd_sc_hd__clkinv_2
XANTENNA__19530__B _19694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21939_ _21939_/A _21939_/B vssd1 vssd1 vccd1 vccd1 _21940_/A sky130_fd_sc_hd__nand2_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21920__A1 _13465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17969__C _20146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _15460_/A _15460_/B vssd1 vssd1 vccd1 vccd1 _15462_/C sky130_fd_sc_hd__xnor2_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12672_ _13116_/C vssd1 vssd1 vccd1 vccd1 _13184_/A sky130_fd_sc_hd__buf_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19326__C1 _19805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14411_ _14380_/Y _14405_/Y _14410_/Y vssd1 vssd1 vccd1 vccd1 _14418_/A sky130_fd_sc_hd__a21boi_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11623_ _11918_/B vssd1 vssd1 vccd1 vccd1 _11711_/B sky130_fd_sc_hd__buf_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15391_ _15391_/A _15391_/B _15435_/A _15435_/B vssd1 vssd1 vccd1 vccd1 _15391_/Y
+ sky130_fd_sc_hd__nor4_4
XANTENNA__12475__A _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_985 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17130_ _16873_/C _16879_/X _16893_/B vssd1 vssd1 vccd1 vccd1 _17220_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__14393__C _14433_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20487__A1 _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11767__A3 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14342_ _14430_/A _14777_/B vssd1 vssd1 vccd1 vccd1 _14355_/A sky130_fd_sc_hd__nand2_1
XFILLER_168_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17061_ _17061_/A vssd1 vssd1 vccd1 vccd1 _17761_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14273_ _14290_/A _14290_/B _14290_/C vssd1 vssd1 vccd1 vccd1 _14273_/X sky130_fd_sc_hd__and3_1
XFILLER_7_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16012_ _16010_/X _15996_/Y _16011_/Y vssd1 vssd1 vccd1 vccd1 _16012_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_143_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13224_ _13259_/A _13224_/B _13264_/B vssd1 vssd1 vccd1 vccd1 _13732_/C sky130_fd_sc_hd__and3_2
XFILLER_170_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13155_ _13168_/C _13168_/D vssd1 vssd1 vccd1 vccd1 _13162_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23189__A0 _14553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12106_ _11654_/A _11875_/A _12105_/Y vssd1 vssd1 vccd1 vccd1 _12107_/A sky130_fd_sc_hd__o21ai_2
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17963_ _17963_/A _18434_/B _17963_/C vssd1 vssd1 vccd1 vccd1 _17966_/A sky130_fd_sc_hd__nand3_2
XFILLER_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13086_ _13072_/Y _13075_/Y _20595_/C _20595_/B vssd1 vssd1 vccd1 vccd1 _13087_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19702_ _19708_/A vssd1 vssd1 vccd1 vccd1 _19819_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17407__A2 _16683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16914_ _16934_/A _16934_/B _16934_/C vssd1 vssd1 vccd1 vccd1 _16930_/B sky130_fd_sc_hd__nand3_4
X_12037_ _15707_/A vssd1 vssd1 vccd1 vccd1 _15706_/A sky130_fd_sc_hd__buf_2
XANTENNA__19801__B1 _19040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17894_ _17896_/C _17896_/B _17893_/X _17764_/X vssd1 vssd1 vccd1 vccd1 _18030_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__16410__A _18503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15418__A1 _15446_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19633_ _23546_/Q _19633_/B _19633_/C vssd1 vssd1 vccd1 vccd1 _19788_/A sky130_fd_sc_hd__nand3b_1
XFILLER_19_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16845_ _16845_/A _16845_/B _16845_/C vssd1 vssd1 vccd1 vccd1 _16885_/A sky130_fd_sc_hd__nand3_1
XFILLER_20_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19564_ _19533_/X _19534_/X _19559_/Y _19560_/Y vssd1 vssd1 vccd1 vccd1 _19567_/A
+ sky130_fd_sc_hd__o22ai_1
X_16776_ _16776_/A _17008_/A _17008_/C vssd1 vssd1 vccd1 vccd1 _16776_/Y sky130_fd_sc_hd__nand3_1
XFILLER_19_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21970__B _21981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13988_ _14790_/B vssd1 vssd1 vccd1 vccd1 _14911_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_53_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18515_ _18518_/A _18518_/B vssd1 vssd1 vccd1 vccd1 _18520_/A sky130_fd_sc_hd__nand2_1
X_15727_ _15662_/B _15727_/B _16798_/B vssd1 vssd1 vccd1 vccd1 _15731_/A sky130_fd_sc_hd__nand3b_2
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12939_ _20669_/A vssd1 vssd1 vccd1 vccd1 _20955_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_19495_ _19951_/D _20061_/A _19328_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19577_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17241__A _19840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15658_ _15920_/D _15918_/B vssd1 vssd1 vccd1 vccd1 _15659_/A sky130_fd_sc_hd__nand2_1
X_18446_ _18446_/A vssd1 vssd1 vccd1 vccd1 _18453_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_179_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15197__A3 _14777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14609_ _15605_/A _14575_/X _14606_/X _14608_/X vssd1 vssd1 vccd1 vccd1 _14609_/X
+ sky130_fd_sc_hd__a211o_1
X_18377_ _18377_/A _18376_/X vssd1 vssd1 vccd1 vccd1 _18378_/A sky130_fd_sc_hd__or2b_1
XFILLER_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15589_ _23514_/Q _15586_/A _15586_/C vssd1 vssd1 vccd1 vccd1 _15590_/B sky130_fd_sc_hd__o21ai_1
XFILLER_187_771 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17328_ _17161_/B _17152_/B _17155_/X _17154_/X vssd1 vssd1 vccd1 vccd1 _17330_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19168__A _19168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17259_ _17259_/A _18607_/C _18607_/A vssd1 vssd1 vccd1 vccd1 _17260_/B sky130_fd_sc_hd__nand3_2
XANTENNA__22219__A2 _22263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20270_ _18211_/B _20365_/A _18211_/A _20263_/A vssd1 vssd1 vccd1 vccd1 _20270_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17646__A2 _17644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11729__A _19161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22927__A0 _23299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19334__C _19539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16606__B1 _16124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22911_ _22911_/A vssd1 vssd1 vccd1 vccd1 _23291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22842_ _22842_/A vssd1 vssd1 vccd1 vccd1 _22843_/B sky130_fd_sc_hd__inv_2
XFILLER_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19020__A1 _16604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_744 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22773_ _22772_/B _22772_/C _22772_/A vssd1 vssd1 vccd1 vccd1 _22808_/A sky130_fd_sc_hd__o21a_1
XANTENNA__17031__B1 _16780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_524 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21724_ _21709_/B _21712_/Y _21705_/X _21679_/X vssd1 vssd1 vccd1 vccd1 _21728_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22992__A _23038_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21655_ _21660_/B _21660_/D vssd1 vssd1 vccd1 vccd1 _21659_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20606_ _20606_/A _20606_/B vssd1 vssd1 vccd1 vccd1 _20607_/C sky130_fd_sc_hd__nand2_1
XFILLER_177_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21586_ _21627_/B _21540_/X _21627_/C _21627_/D vssd1 vssd1 vccd1 vccd1 _21586_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23325_ _23325_/CLK _23325_/D vssd1 vssd1 vccd1 vccd1 _23325_/Q sky130_fd_sc_hd__dfxtp_2
X_20537_ _13053_/X _20676_/A _20533_/B _20670_/A vssd1 vssd1 vccd1 vccd1 _20542_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15896__A1 _15985_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20468_ _13029_/A _13003_/B _21070_/A _13001_/A vssd1 vssd1 vccd1 vccd1 _20484_/A
+ sky130_fd_sc_hd__a31o_1
X_23256_ _23256_/A _23256_/B vssd1 vssd1 vccd1 vccd1 _23257_/A sky130_fd_sc_hd__and2_1
XFILLER_146_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11639__A _11936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13371__A2 _22186_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22207_ _22207_/A _22207_/B _22207_/C vssd1 vssd1 vccd1 vccd1 _22225_/A sky130_fd_sc_hd__nand3_1
XFILLER_134_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18834__A1 _11822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20399_ _20371_/B _20269_/B _20369_/X _20428_/A vssd1 vssd1 vccd1 vccd1 _20403_/A
+ sky130_fd_sc_hd__a31oi_2
X_23187_ _16510_/C input7/X _23195_/S vssd1 vssd1 vccd1 vccd1 _23188_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22138_ _22139_/A _22139_/B _22139_/C vssd1 vssd1 vccd1 vccd1 _22215_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__22918__A0 _12875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14960_ _14960_/A _14960_/B vssd1 vssd1 vccd1 vccd1 _14965_/B sky130_fd_sc_hd__nor2_1
X_22069_ _22208_/A _22208_/B _22208_/C vssd1 vssd1 vccd1 vccd1 _22069_/Y sky130_fd_sc_hd__nand3_1
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13911_ _13940_/B _13946_/A _13911_/C vssd1 vssd1 vccd1 vccd1 _14069_/A sky130_fd_sc_hd__nand3_1
XANTENNA__13573__B _22553_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input29_A wb_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ _14893_/B _15305_/A _15175_/C vssd1 vssd1 vccd1 vccd1 _14891_/Y sky130_fd_sc_hd__nand3_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12882__A1 _20894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16630_ _16837_/A _16837_/B _16837_/C vssd1 vssd1 vccd1 vccd1 _16649_/A sky130_fd_sc_hd__nand3_1
XFILLER_75_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13842_ _13842_/A _13842_/B vssd1 vssd1 vccd1 vccd1 _13843_/C sky130_fd_sc_hd__nand2_1
XFILLER_90_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16561_ _16564_/B _16542_/Y _16560_/Y vssd1 vssd1 vccd1 vccd1 _16562_/B sky130_fd_sc_hd__a21oi_1
X_13773_ _13243_/Y _13658_/Y _13666_/A vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__o21ai_1
XFILLER_16_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18157__A _18163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18300_ _18305_/A _18305_/B vssd1 vssd1 vccd1 vccd1 _18301_/B sky130_fd_sc_hd__nor2_1
X_15512_ _15513_/C _15536_/B _15513_/B _15513_/D vssd1 vssd1 vccd1 vccd1 _15517_/A
+ sky130_fd_sc_hd__o22ai_2
X_19280_ _19280_/A vssd1 vssd1 vccd1 vccd1 _19924_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12724_ _12724_/A _20966_/B _20781_/C vssd1 vssd1 vccd1 vccd1 _12725_/A sky130_fd_sc_hd__nand3_4
X_16492_ _16492_/A _16492_/B vssd1 vssd1 vccd1 vccd1 _16492_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17573__A1 _16356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18231_ _18269_/A _18231_/B vssd1 vssd1 vccd1 vccd1 _18236_/C sky130_fd_sc_hd__and2_1
XFILLER_176_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15443_ _15434_/B _15438_/B _15432_/Y vssd1 vssd1 vccd1 vccd1 _15476_/A sky130_fd_sc_hd__a21oi_4
XFILLER_176_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12655_ _12634_/X _12648_/X _12651_/X _12652_/X _12654_/Y vssd1 vssd1 vccd1 vccd1
+ _12662_/B sky130_fd_sc_hd__o221ai_1
XFILLER_169_760 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18162_ _20217_/A _17723_/A _17723_/B _20215_/A _18161_/B vssd1 vssd1 vccd1 vccd1
+ _18163_/D sky130_fd_sc_hd__a32o_1
XFILLER_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11606_ _11656_/B vssd1 vssd1 vccd1 vccd1 _11606_/X sky130_fd_sc_hd__buf_2
X_15374_ _15422_/A _15427_/A _15373_/X vssd1 vssd1 vccd1 vccd1 _15377_/A sky130_fd_sc_hd__o21ai_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17325__A1 _16549_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12586_ _12683_/B vssd1 vssd1 vccd1 vccd1 _12875_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_129_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17113_ _17302_/A _17301_/A _17123_/C vssd1 vssd1 vccd1 vccd1 _17113_/X sky130_fd_sc_hd__and3_1
X_14325_ _14367_/C _14325_/B _14367_/B vssd1 vssd1 vccd1 vccd1 _14365_/A sky130_fd_sc_hd__nand3_1
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18093_ _18093_/A _19967_/C _18172_/C _18172_/D vssd1 vssd1 vccd1 vccd1 _18101_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_156_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17044_ _15742_/X _16447_/B _17434_/A _17435_/A _18947_/A vssd1 vssd1 vccd1 vccd1
+ _17252_/A sky130_fd_sc_hd__o221ai_4
XFILLER_143_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output97_A _23580_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14256_ _14256_/A _14324_/B vssd1 vssd1 vccd1 vccd1 _14367_/A sky130_fd_sc_hd__xor2_1
XFILLER_171_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13207_ _12987_/Y _13099_/Y _13100_/X _13208_/B _13208_/A vssd1 vssd1 vccd1 vccd1
+ _13210_/A sky130_fd_sc_hd__o32a_1
XANTENNA__17628__A2 _15933_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14187_ _14187_/A _14187_/B _14187_/C vssd1 vssd1 vccd1 vccd1 _14220_/B sky130_fd_sc_hd__nand3_4
XANTENNA__18620__A _18620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1162 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13467__C _13660_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _13138_/A _13138_/B _13138_/C _13138_/D vssd1 vssd1 vccd1 vccd1 _13140_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _23396_/Q vssd1 vssd1 vccd1 vccd1 _18996_/C sky130_fd_sc_hd__inv_2
XFILLER_86_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13764__A _13766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17236__A _17420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _18154_/A _17944_/Y _23527_/Q _17945_/Y vssd1 vssd1 vccd1 vccd1 _17946_/X
+ sky130_fd_sc_hd__o211a_1
X_13069_ _13055_/X _13060_/X _13061_/Y vssd1 vssd1 vccd1 vccd1 _20565_/D sky130_fd_sc_hd__o21ai_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16140__A _16140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15682__C _15974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17877_ _17610_/X _17752_/A _17710_/X _17760_/B _17754_/Y vssd1 vssd1 vccd1 vccd1
+ _17878_/B sky130_fd_sc_hd__o221ai_1
XFILLER_94_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19616_ _19616_/A _19616_/B vssd1 vssd1 vccd1 vccd1 _19638_/C sky130_fd_sc_hd__nand2_1
XANTENNA__14298__C _14298_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16828_ _16828_/A _17064_/A vssd1 vssd1 vccd1 vccd1 _16828_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19002__A1 _18439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19547_ _19547_/A vssd1 vssd1 vccd1 vccd1 _19547_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16759_ _16768_/A _16759_/B _16759_/C vssd1 vssd1 vccd1 vccd1 _16759_/Y sky130_fd_sc_hd__nand3_1
XFILLER_179_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19478_ _19478_/A vssd1 vssd1 vccd1 vccd1 _19670_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_94_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18429_ _18429_/A _18429_/B vssd1 vssd1 vccd1 vccd1 _18433_/A sky130_fd_sc_hd__nand2_1
XFILLER_181_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19305__A2 _11801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21440_ _21500_/A _21440_/B _21440_/C _21448_/B vssd1 vssd1 vccd1 vccd1 _21442_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__17316__A1 _16464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17316__B2 _17305_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18513__B1 _17712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12265__D _17134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21371_ _21546_/A _21371_/B _21371_/C _21440_/B vssd1 vssd1 vccd1 vccd1 _21371_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_119_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16315__A _16315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15878__A1 _20142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20322_ _20322_/A _20322_/B vssd1 vssd1 vccd1 vccd1 _20323_/C sky130_fd_sc_hd__xnor2_1
X_23110_ _23381_/Q input31/X _23110_/S vssd1 vssd1 vccd1 vccd1 _23111_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20253_ _20252_/A _20252_/B _20252_/C vssd1 vssd1 vccd1 vccd1 _20253_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__17619__A2 _16478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23041_ _23097_/A vssd1 vssd1 vccd1 vccd1 _23110_/S sky130_fd_sc_hd__buf_2
XFILLER_115_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20184_ _20184_/A _20184_/B vssd1 vssd1 vccd1 vccd1 _20186_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21891__A _21891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19361__A _19361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22128__A1 _13547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20139__B1 _17414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22825_ _22856_/A _22856_/D _22856_/C vssd1 vssd1 vccd1 vccd1 _22854_/B sky130_fd_sc_hd__nand3_1
XFILLER_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21887__B1 _22365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22756_ _22756_/A _22756_/B _22756_/C _22756_/D vssd1 vssd1 vccd1 vccd1 _22764_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_73_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21707_ _21705_/X _21679_/X _21709_/B vssd1 vssd1 vccd1 vccd1 _21723_/B sky130_fd_sc_hd__a21o_1
XFILLER_158_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22687_ _22749_/A _22749_/B vssd1 vssd1 vccd1 vccd1 _22687_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12440_ _16661_/C _19010_/A _19193_/C vssd1 vssd1 vccd1 vccd1 _12441_/B sky130_fd_sc_hd__and3_1
XFILLER_139_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21638_ _21668_/B _21432_/A _21432_/B _21637_/A _21635_/X vssd1 vssd1 vccd1 vccd1
+ _21638_/X sky130_fd_sc_hd__a32o_1
XFILLER_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12371_ _12363_/A _12363_/B _12363_/C _12363_/D vssd1 vssd1 vccd1 vccd1 _12372_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21569_ _21611_/A _21577_/C vssd1 vssd1 vccd1 vccd1 _21569_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15767__C _16619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ _14108_/Y _15085_/B _15085_/C _14039_/A vssd1 vssd1 vccd1 vccd1 _14110_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_10_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23308_ _23309_/CLK _23308_/D vssd1 vssd1 vccd1 vccd1 _23308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15090_ _15090_/A _15090_/B vssd1 vssd1 vccd1 vccd1 _15090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14541__A1 _21832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041_ _14009_/X _14020_/Y _14063_/A vssd1 vssd1 vccd1 vccd1 _14056_/A sky130_fd_sc_hd__o21ai_1
XFILLER_181_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23239_ _23438_/Q input23/X _23239_/S vssd1 vssd1 vccd1 vccd1 _23240_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18807__A1 _12130_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22603__A2 _22756_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18283__A2 _18335_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17800_ _17798_/X _17799_/Y _17779_/Y _17786_/Y vssd1 vssd1 vccd1 vccd1 _17801_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18780_ _19073_/A _18781_/B _18882_/A vssd1 vssd1 vccd1 vccd1 _18889_/A sky130_fd_sc_hd__a21oi_4
X_15992_ _16443_/C vssd1 vssd1 vccd1 vccd1 _17450_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_94_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17731_ _17634_/B _17728_/X _17838_/B _17725_/Y _17629_/Y vssd1 vssd1 vccd1 vccd1
+ _17781_/B sky130_fd_sc_hd__o2111ai_1
X_14943_ _14943_/A _14943_/B _14966_/B vssd1 vssd1 vccd1 vccd1 _14945_/B sky130_fd_sc_hd__nand3_1
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16046__A1 _16194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23551__CLK _23558_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17662_ _17662_/A vssd1 vssd1 vccd1 vccd1 _17662_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14874_ _14874_/A _14903_/A vssd1 vssd1 vccd1 vccd1 _14899_/A sky130_fd_sc_hd__nand2_1
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22119__A1 _21936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19401_ _19401_/A vssd1 vssd1 vccd1 vccd1 _19401_/Y sky130_fd_sc_hd__inv_2
X_16613_ _12513_/A _12511_/A _16612_/A _17594_/A vssd1 vssd1 vccd1 vccd1 _16828_/A
+ sky130_fd_sc_hd__o211ai_4
X_13825_ _21923_/A _22064_/C _21924_/A vssd1 vssd1 vccd1 vccd1 _13825_/Y sky130_fd_sc_hd__nand3_1
XFILLER_63_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17593_ _17593_/A vssd1 vssd1 vccd1 vccd1 _17593_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__20210__A _20210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19332_ _19332_/A _19332_/B _19332_/C vssd1 vssd1 vccd1 vccd1 _19340_/A sky130_fd_sc_hd__nand3_2
XANTENNA__19535__A2 _11841_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16544_ _16544_/A _16544_/B vssd1 vssd1 vccd1 vccd1 _16544_/Y sky130_fd_sc_hd__nand2_1
X_13756_ _13756_/A _13756_/B vssd1 vssd1 vccd1 vccd1 _13756_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16119__B _16153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _12703_/X _12706_/Y _13041_/B _13184_/A _12812_/A vssd1 vssd1 vccd1 vccd1
+ _13138_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_188_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19263_ _19263_/A _19614_/A _19900_/A vssd1 vssd1 vccd1 vccd1 _19263_/X sky130_fd_sc_hd__and3_1
X_16475_ _16474_/B _16475_/B _16475_/C vssd1 vssd1 vccd1 vccd1 _16476_/C sky130_fd_sc_hd__nand3b_1
X_13687_ _13864_/A _22663_/D _13743_/A vssd1 vssd1 vccd1 vccd1 _21839_/B sky130_fd_sc_hd__and3_1
XANTENNA__15021__A2 _15195_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18214_ _18286_/A _18214_/B vssd1 vssd1 vccd1 vccd1 _18226_/A sky130_fd_sc_hd__nand2_1
XFILLER_176_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15426_ _15426_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15451_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19194_ _11936_/X _19196_/B _19195_/A vssd1 vssd1 vccd1 vccd1 _19194_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14765__D1 _15301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12638_ _23292_/Q vssd1 vssd1 vccd1 vccd1 _12712_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18145_ _18054_/Y _18057_/Y _18060_/Y vssd1 vssd1 vccd1 vccd1 _18145_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17849__A2 _17741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15357_ _15459_/B _15488_/B _15459_/A vssd1 vssd1 vccd1 vccd1 _15357_/X sky130_fd_sc_hd__or3_1
XANTENNA__14780__A1 _14245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12569_ _23450_/Q vssd1 vssd1 vccd1 vccd1 _20628_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_184_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14308_ _14842_/A _14309_/C _14310_/A vssd1 vssd1 vccd1 vccd1 _14846_/A sky130_fd_sc_hd__a21bo_1
X_18076_ _18161_/C _17406_/B _17406_/A _18001_/X _18211_/D vssd1 vssd1 vccd1 vccd1
+ _18084_/A sky130_fd_sc_hd__a311o_1
XFILLER_172_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21976__A _21976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15288_ _15288_/A _15288_/B vssd1 vssd1 vccd1 vccd1 _15402_/B sky130_fd_sc_hd__xnor2_4
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17027_ _17025_/Y _17026_/Y _17369_/A vssd1 vssd1 vccd1 vccd1 _17027_/Y sky130_fd_sc_hd__a21boi_1
X_14239_ _15254_/B vssd1 vssd1 vccd1 vccd1 _15082_/D sky130_fd_sc_hd__buf_2
XFILLER_171_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17394__A1_N _17140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19165__B _19308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18978_ _18978_/A _18978_/B vssd1 vssd1 vccd1 vccd1 _18983_/B sky130_fd_sc_hd__nand2_1
XFILLER_105_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _17540_/X _17686_/X _17832_/D _17835_/X vssd1 vssd1 vccd1 vccd1 _17929_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20940_ _20940_/A _20940_/B _20940_/C vssd1 vssd1 vccd1 vccd1 _20940_/X sky130_fd_sc_hd__and3_1
XFILLER_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16588__A2 _12223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20871_ _21157_/B _20754_/A _20865_/Y _20870_/X vssd1 vssd1 vccd1 vccd1 _21017_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22610_ _22610_/A _22633_/B vssd1 vssd1 vccd1 vccd1 _22611_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23590_ _23598_/CLK _23590_/D vssd1 vssd1 vccd1 vccd1 _23590_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13271__A1 _13226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13660__C _13660_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22541_ _22541_/A _22541_/B _22541_/C _22541_/D vssd1 vssd1 vccd1 vccd1 _22541_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_50_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22472_ _22475_/C _22475_/D vssd1 vssd1 vccd1 vccd1 _22473_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13940__A_N _13911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21423_ _21342_/Y _21343_/Y _21411_/A _21411_/B vssd1 vssd1 vccd1 vccd1 _21423_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__18498__C1 _18465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13574__A2 _13527_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18501__A3 _15882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21354_ _21354_/A _21402_/B vssd1 vssd1 vccd1 vccd1 _21354_/X sky130_fd_sc_hd__and2_1
XFILLER_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20305_ _20359_/A _20359_/B vssd1 vssd1 vccd1 vccd1 _20313_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15884__A _15884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22046__B1 _21913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21285_ _21279_/Y _21285_/B _21285_/C vssd1 vssd1 vccd1 vccd1 _21285_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23024_ _23024_/A vssd1 vssd1 vccd1 vccd1 _23342_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13731__C1 _13415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20236_ _20234_/Y _20235_/X _20176_/C _20179_/X vssd1 vssd1 vccd1 vccd1 _20236_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11888__A2 _11885_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11917__A _23589_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20167_ _20167_/A _20167_/B _20232_/A vssd1 vssd1 vccd1 vccd1 _20229_/B sky130_fd_sc_hd__nand3_1
XFILLER_104_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20098_ _20099_/B _20177_/A _20097_/Y vssd1 vssd1 vccd1 vccd1 _20103_/C sky130_fd_sc_hd__a21bo_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _16591_/A vssd1 vssd1 vccd1 vccd1 _18503_/A sky130_fd_sc_hd__buf_4
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11871_ _11871_/A vssd1 vssd1 vccd1 vccd1 _12373_/A sky130_fd_sc_hd__buf_4
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _21766_/A _21767_/A _22039_/C vssd1 vssd1 vccd1 vccd1 _13610_/Y sky130_fd_sc_hd__nand3_4
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22808_ _22808_/A _22808_/B _22808_/C vssd1 vssd1 vccd1 vccd1 _22808_/Y sky130_fd_sc_hd__nor3_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _13349_/X _14550_/X _14647_/A _15713_/C _14589_/X vssd1 vssd1 vccd1 vccd1
+ _14590_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12467__B _16122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ _13538_/A _13538_/B _13598_/A _13477_/X vssd1 vssd1 vccd1 vccd1 _13541_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22739_ _22736_/X _22738_/Y _23280_/Q vssd1 vssd1 vccd1 vccd1 _22821_/B sky130_fd_sc_hd__o21ai_2
XFILLER_186_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11812__A2 _11807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18435__A _18435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16260_ _16258_/C _16258_/B _16258_/A vssd1 vssd1 vccd1 vccd1 _16260_/Y sky130_fd_sc_hd__a21oi_2
X_13472_ _13341_/X _13320_/X _13470_/X _22096_/B vssd1 vssd1 vccd1 vccd1 _13472_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_186_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22371__A1_N _13527_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15211_ _15282_/A _15211_/B _15282_/B vssd1 vssd1 vccd1 vccd1 _15211_/Y sky130_fd_sc_hd__nand3_1
X_12423_ _12423_/A _12423_/B vssd1 vssd1 vccd1 vccd1 _12445_/A sky130_fd_sc_hd__nand2_1
X_16191_ _16191_/A _16195_/A vssd1 vssd1 vccd1 vccd1 _16671_/B sky130_fd_sc_hd__nand2_1
XFILLER_166_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15142_ _15053_/A _15064_/B _15053_/B vssd1 vssd1 vccd1 vccd1 _15144_/A sky130_fd_sc_hd__a21bo_1
X_12354_ _12353_/X _12379_/A _12314_/Y _12310_/A vssd1 vssd1 vccd1 vccd1 _12355_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_138_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16503__A2 _15856_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19950_ _16408_/A _19838_/A _20079_/A vssd1 vssd1 vccd1 vccd1 _19951_/C sky130_fd_sc_hd__o21ai_1
X_15073_ _14962_/A _14965_/B _15220_/B _15439_/C vssd1 vssd1 vccd1 vccd1 _15148_/A
+ sky130_fd_sc_hd__o31a_1
X_12285_ _12374_/A _12238_/X _12284_/Y _11682_/Y _11717_/C vssd1 vssd1 vccd1 vccd1
+ _12285_/X sky130_fd_sc_hd__o221a_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18901_ _18751_/X _18752_/X _18878_/Y _18886_/Y vssd1 vssd1 vccd1 vccd1 _18901_/X
+ sky130_fd_sc_hd__o211a_1
X_14024_ _14086_/B _14024_/B _23355_/Q vssd1 vssd1 vccd1 vccd1 _14035_/A sky130_fd_sc_hd__nand3_1
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19881_ _19796_/A _19796_/B _19880_/Y vssd1 vssd1 vccd1 vccd1 _19889_/A sky130_fd_sc_hd__o21ai_2
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20063__A2 _20210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18832_ _18635_/Y _18796_/X _18804_/B vssd1 vssd1 vccd1 vccd1 _18832_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16121__C _16840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18008__A2 _17323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19205__A1 _19203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18763_ _18763_/A _18763_/B vssd1 vssd1 vccd1 vccd1 _18767_/A sky130_fd_sc_hd__nand2_1
X_15975_ _15975_/A _15975_/B vssd1 vssd1 vccd1 vccd1 _16172_/A sky130_fd_sc_hd__nand2_4
XFILLER_110_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22420__A _22420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_430 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17714_ _17714_/A vssd1 vssd1 vccd1 vccd1 _17899_/A sky130_fd_sc_hd__clkbuf_2
X_14926_ _14926_/A _14926_/B _14926_/C vssd1 vssd1 vccd1 vccd1 _14927_/D sky130_fd_sc_hd__nand3_1
XFILLER_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18694_ _18529_/A _18522_/A _18522_/B _18528_/Y vssd1 vssd1 vccd1 vccd1 _18751_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17645_ _19670_/A vssd1 vssd1 vccd1 vccd1 _20081_/A sky130_fd_sc_hd__buf_2
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14857_ _14857_/A _14857_/B vssd1 vssd1 vccd1 vccd1 _14900_/A sky130_fd_sc_hd__nand2_1
XFILLER_90_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19508__A2 _19307_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13808_ _13366_/B _13602_/Y _13603_/X vssd1 vssd1 vccd1 vccd1 _13809_/B sky130_fd_sc_hd__o21ai_1
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17576_ _19694_/A vssd1 vssd1 vccd1 vccd1 _20133_/D sky130_fd_sc_hd__buf_2
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14788_ _14788_/A _14857_/A _14788_/C vssd1 vssd1 vccd1 vccd1 _14857_/B sky130_fd_sc_hd__nand3_1
XFILLER_56_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19315_ _16437_/X _19858_/A _19491_/A _19314_/Y vssd1 vssd1 vccd1 vccd1 _19517_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_177_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16527_ _12346_/A _16536_/B _16528_/A _16544_/A vssd1 vssd1 vccd1 vccd1 _16529_/A
+ sky130_fd_sc_hd__a22o_1
X_13739_ _13739_/A _13739_/B _13739_/C vssd1 vssd1 vccd1 vccd1 _13739_/Y sky130_fd_sc_hd__nor3_1
XFILLER_91_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19246_ _19246_/A vssd1 vssd1 vccd1 vccd1 _19246_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16458_ _16458_/A vssd1 vssd1 vccd1 vccd1 _16458_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13005__B2 _20781_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23447__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12213__C1 _19648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15409_ _15409_/A _15511_/C vssd1 vssd1 vccd1 vccd1 _15413_/A sky130_fd_sc_hd__nand2_1
XFILLER_129_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16389_ _16389_/A vssd1 vssd1 vccd1 vccd1 _16389_/X sky130_fd_sc_hd__buf_2
X_19177_ _19186_/A _18992_/B _19186_/B vssd1 vssd1 vccd1 vccd1 _19177_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_118_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18999__B _23396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18128_ _17924_/A _17924_/B _17924_/C _18045_/A vssd1 vssd1 vccd1 vccd1 _18132_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_118_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18059_ _18059_/A _18059_/B _18072_/B vssd1 vssd1 vccd1 vccd1 _18060_/B sky130_fd_sc_hd__and3_1
XANTENNA__23597__CLK _23598_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18080__A _18080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21070_ _21070_/A vssd1 vssd1 vccd1 vccd1 _21365_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20021_ _20021_/A _20113_/A vssd1 vssd1 vccd1 vccd1 _20185_/A sky130_fd_sc_hd__or2b_1
XFILLER_141_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11737__A _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22968__C input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20769__B _21124_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13952__A _14246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17424__A _17959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21972_ _21972_/A vssd1 vssd1 vccd1 vccd1 _21980_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18955__B1 _18944_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20923_ _21036_/A vssd1 vssd1 vccd1 vccd1 _21281_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20854_ _20854_/A _20854_/B vssd1 vssd1 vccd1 vccd1 _20856_/B sky130_fd_sc_hd__nand2_1
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12287__B _12297_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23573_ _23578_/CLK _23573_/D vssd1 vssd1 vccd1 vccd1 _23573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20785_ _20778_/X _20920_/A _20783_/Y _20790_/B vssd1 vssd1 vccd1 vccd1 _20789_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__19380__B1 _17431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22524_ _22524_/A _22524_/B _22524_/C _22524_/D vssd1 vssd1 vccd1 vccd1 _22525_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_194_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20935__D _21177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22208__C _22208_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22455_ _22455_/A vssd1 vssd1 vccd1 vccd1 _22529_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21406_ _21335_/A _21354_/X _21404_/B _21404_/A vssd1 vssd1 vccd1 vccd1 _21407_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_109_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22386_ _22386_/A _22386_/B vssd1 vssd1 vccd1 vccd1 _22386_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20293__A2 _20243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21337_ _21264_/Y _21240_/A _21342_/C vssd1 vssd1 vccd1 vccd1 _21340_/A sky130_fd_sc_hd__o21ai_1
XFILLER_190_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12070_ _23258_/B vssd1 vssd1 vccd1 vccd1 _12070_/Y sky130_fd_sc_hd__inv_2
X_21268_ _21268_/A _21387_/B vssd1 vssd1 vccd1 vccd1 _21270_/C sky130_fd_sc_hd__nand2_1
XFILLER_104_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23007_ _23007_/A vssd1 vssd1 vccd1 vccd1 _23334_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11647__A _11960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20219_ _20048_/Y _20139_/Y _20216_/X _20218_/Y _20148_/A vssd1 vssd1 vccd1 vccd1
+ _20219_/X sky130_fd_sc_hd__o221a_1
XFILLER_173_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21199_ _20509_/B _21190_/X _21195_/X _21198_/Y vssd1 vssd1 vccd1 vccd1 _21267_/C
+ sky130_fd_sc_hd__o22ai_2
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22990__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13862__A _22713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_bq_clk_i clkbuf_4_9_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _23582_/CLK
+ sky130_fd_sc_hd__clkbuf_8
X_15760_ _15750_/Y _15754_/X _15759_/X vssd1 vssd1 vccd1 vccd1 _15760_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12972_ _12972_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _13141_/C sky130_fd_sc_hd__xor2_2
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17749__A1 _17285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18946__B1 _12353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input11_A wb_dat_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11923_ _11916_/X _11921_/Y _15841_/B vssd1 vssd1 vccd1 vccd1 _11924_/A sky130_fd_sc_hd__o21ai_1
X_14711_ _23410_/Q _14693_/X _14698_/X _23442_/Q _14710_/X vssd1 vssd1 vccd1 vccd1
+ _14711_/X sky130_fd_sc_hd__a221o_2
XFILLER_46_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _15691_/A vssd1 vssd1 vccd1 vccd1 _16315_/A sky130_fd_sc_hd__buf_2
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22894__B _22895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _17430_/A vssd1 vssd1 vccd1 vccd1 _17487_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _22896_/D vssd1 vssd1 vccd1 vccd1 _14642_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11854_ _15707_/B vssd1 vssd1 vccd1 vccd1 _16365_/A sky130_fd_sc_hd__buf_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15775__A3 _17409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17361_ _17359_/B _17361_/B _17514_/A vssd1 vssd1 vccd1 vccd1 _17362_/C sky130_fd_sc_hd__nand3b_1
X_14573_ _23419_/Q vssd1 vssd1 vccd1 vccd1 _15674_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_198_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14693__A _14693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11785_ _12145_/A vssd1 vssd1 vccd1 vccd1 _18755_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19100_ _19100_/A vssd1 vssd1 vccd1 vccd1 _19104_/A sky130_fd_sc_hd__inv_2
XFILLER_159_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11797__A1 _16049_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16312_ _16464_/A _16311_/X _16309_/A _16309_/B vssd1 vssd1 vccd1 vccd1 _16313_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_14_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13524_ _13732_/C vssd1 vssd1 vccd1 vccd1 _21815_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_159_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17292_ _17292_/A _17292_/B vssd1 vssd1 vccd1 vccd1 _17292_/Y sky130_fd_sc_hd__nand2_1
XFILLER_198_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16724__A2 _16723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19031_ _18675_/A _19218_/A _19203_/A _19196_/A vssd1 vssd1 vccd1 vccd1 _19031_/X
+ sky130_fd_sc_hd__o22a_1
X_16243_ _16243_/A _16253_/A vssd1 vssd1 vccd1 vccd1 _16243_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13455_ _22035_/C vssd1 vssd1 vccd1 vccd1 _22269_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_3_0_bq_clk_i_A clkbuf_4_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ _23392_/Q vssd1 vssd1 vccd1 vccd1 _18810_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16174_ _16168_/C _16174_/B _16174_/C vssd1 vssd1 vccd1 vccd1 _16175_/C sky130_fd_sc_hd__nand3b_1
XANTENNA__18477__A2 _18434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13386_ _21883_/A _13804_/B _22521_/C vssd1 vssd1 vccd1 vccd1 _13434_/B sky130_fd_sc_hd__and3_2
XFILLER_182_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19708__B _19708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15125_ _15124_/Y _15013_/D _15013_/C vssd1 vssd1 vccd1 vccd1 _15127_/A sky130_fd_sc_hd__a21bo_1
X_12337_ _12360_/A _12360_/B _12381_/C _12381_/B vssd1 vssd1 vccd1 vccd1 _12337_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22134__B _22476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19933_ _19909_/A _19909_/B _19909_/C _19769_/Y _19932_/Y vssd1 vssd1 vccd1 vccd1
+ _19933_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15056_ _15408_/A _14944_/B _14933_/A _14939_/B vssd1 vssd1 vccd1 vccd1 _15064_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18229__A2 _18157_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19426__A1 _12508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12268_ _19323_/A vssd1 vssd1 vccd1 vccd1 _19675_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12660__B _20966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14007_ _14007_/A _14007_/B vssd1 vssd1 vccd1 vccd1 _14236_/B sky130_fd_sc_hd__xnor2_1
X_19864_ _19864_/A _19864_/B _19864_/C vssd1 vssd1 vccd1 vccd1 _19873_/C sky130_fd_sc_hd__nand3_1
X_12199_ _12199_/A _12199_/B _12199_/C _12199_/D vssd1 vssd1 vccd1 vccd1 _12203_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput90 _23264_/Q vssd1 vssd1 vccd1 vccd1 y[2] sky130_fd_sc_hd__buf_2
XFILLER_150_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18815_ _18996_/B vssd1 vssd1 vccd1 vccd1 _19504_/A sky130_fd_sc_hd__clkbuf_4
X_19795_ _19744_/X _19743_/X _19750_/Y _19749_/Y vssd1 vssd1 vccd1 vccd1 _19894_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18746_ _18746_/A vssd1 vssd1 vccd1 vccd1 _23521_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15958_ _16612_/B vssd1 vssd1 vccd1 vccd1 _17061_/A sky130_fd_sc_hd__buf_2
XANTENNA__18059__B _18059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14909_ _14909_/A _14909_/B _14909_/C vssd1 vssd1 vccd1 vccd1 _14927_/B sky130_fd_sc_hd__nand3_1
X_18677_ _19203_/A _15882_/A _18503_/Y vssd1 vssd1 vccd1 vccd1 _18677_/Y sky130_fd_sc_hd__o21ai_2
X_15889_ _12222_/X _12223_/X _15864_/A vssd1 vssd1 vccd1 vccd1 _15889_/X sky130_fd_sc_hd__a21o_2
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17628_ _16781_/B _15933_/Y _17625_/C _19840_/A vssd1 vssd1 vccd1 vccd1 _17628_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17898__B _19957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15699__A _15699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17559_ _17558_/X _17555_/A _17806_/A vssd1 vssd1 vccd1 vccd1 _17559_/Y sky130_fd_sc_hd__o21ai_1
X_20570_ _20570_/A vssd1 vssd1 vccd1 vccd1 _20736_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19229_ _19206_/X _19202_/Y _19213_/Y _19189_/X _19228_/X vssd1 vssd1 vccd1 vccd1
+ _19232_/A sky130_fd_sc_hd__o2111ai_1
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14108__A _23497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18803__A _18803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22240_ _22240_/A _22240_/B vssd1 vssd1 vccd1 vccd1 _22242_/A sky130_fd_sc_hd__nand2_1
XFILLER_192_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22171_ _22057_/X _22168_/X _22381_/C _22391_/A vssd1 vssd1 vccd1 vccd1 _22171_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_132_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21122_ _20773_/A _20773_/C _21124_/A _21514_/A _21125_/A vssd1 vssd1 vccd1 vccd1
+ _21123_/C sky130_fd_sc_hd__a41o_1
XFILLER_133_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21053_ _21053_/A _21053_/B _21053_/C vssd1 vssd1 vccd1 vccd1 _21212_/A sky130_fd_sc_hd__nand3_4
XFILLER_143_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20004_ _19939_/Y _19940_/X _20011_/B _20011_/A vssd1 vssd1 vccd1 vccd1 _20004_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_100_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input3_A wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1159 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21955_ _22089_/A _21982_/B vssd1 vssd1 vccd1 vccd1 _21956_/A sky130_fd_sc_hd__nand2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20906_ _20906_/A vssd1 vssd1 vccd1 vccd1 _20906_/X sky130_fd_sc_hd__buf_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19800__C _19800_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21886_ _22121_/A _13492_/A _21885_/Y vssd1 vssd1 vccd1 vccd1 _21984_/C sky130_fd_sc_hd__o21ai_2
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20837_ _20837_/A vssd1 vssd1 vccd1 vccd1 _20842_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__22488__B1 _22647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_650 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23556_ _23558_/CLK _23556_/D vssd1 vssd1 vccd1 vccd1 _23556_/Q sky130_fd_sc_hd__dfxtp_1
X_11570_ _23586_/Q _23585_/Q vssd1 vssd1 vccd1 vccd1 _11918_/B sky130_fd_sc_hd__nor2_2
X_20768_ _21030_/A _21030_/C vssd1 vssd1 vccd1 vccd1 _20880_/A sky130_fd_sc_hd__nand2_1
XFILLER_196_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22507_ _22090_/A _13599_/X _22505_/B _22506_/X vssd1 vssd1 vccd1 vccd1 _22507_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_196_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23487_ _23499_/CLK _23499_/Q vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
X_20699_ _20699_/A _20699_/B _20699_/C vssd1 vssd1 vccd1 vccd1 _20718_/A sky130_fd_sc_hd__nand3_2
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _13247_/D vssd1 vssd1 vccd1 vccd1 _13680_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22438_ _22242_/A _22242_/B _22242_/C _22342_/B vssd1 vssd1 vccd1 vccd1 _22438_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_182_146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17974__D _17974_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12183__D _16674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13171_ _13171_/A _13171_/B vssd1 vssd1 vccd1 vccd1 _13171_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22369_ _22297_/B _22368_/Y _22647_/A _22362_/Y _22548_/A vssd1 vssd1 vccd1 vccd1
+ _22496_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_123_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12122_ _18836_/A _18836_/B _12130_/A vssd1 vssd1 vccd1 vccd1 _12122_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13153__B1 _12634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18616__C1 _18615_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16930_ _16935_/A _16930_/B _16936_/B _16936_/C vssd1 vssd1 vccd1 vccd1 _17166_/B
+ sky130_fd_sc_hd__nand4_4
X_12053_ _12053_/A vssd1 vssd1 vccd1 vccd1 _12053_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_120_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18092__B1 _18093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16861_ _15644_/X _15791_/X _11971_/X _11972_/X _15647_/B vssd1 vssd1 vccd1 vccd1
+ _16861_/X sky130_fd_sc_hd__a221o_1
XANTENNA__14688__A _14688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18600_ _18600_/A _18600_/B _18600_/C vssd1 vssd1 vccd1 vccd1 _18601_/A sky130_fd_sc_hd__nand3_2
XFILLER_19_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15812_ _15761_/X _15762_/Y _15763_/Y _15706_/A _16365_/A vssd1 vssd1 vccd1 vccd1
+ _15813_/B sky130_fd_sc_hd__o2111ai_2
X_19580_ _19207_/X _19196_/Y _19345_/A _19345_/B _19201_/C vssd1 vssd1 vccd1 vccd1
+ _19580_/Y sky130_fd_sc_hd__o2111ai_1
X_16792_ _16792_/A _16792_/B vssd1 vssd1 vccd1 vccd1 _17365_/C sky130_fd_sc_hd__nor2_1
XFILLER_133_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18531_ _18531_/A vssd1 vssd1 vccd1 vccd1 _19262_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15743_ _15729_/X _16187_/A _15662_/C vssd1 vssd1 vccd1 vccd1 _15766_/A sky130_fd_sc_hd__o21a_1
X_12955_ _12950_/X _12952_/X _12954_/Y vssd1 vssd1 vccd1 vccd1 _12955_/Y sky130_fd_sc_hd__a21oi_2
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _12254_/A vssd1 vssd1 vccd1 vccd1 _11906_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18462_ _18462_/A _18462_/B vssd1 vssd1 vccd1 vccd1 _18464_/B sky130_fd_sc_hd__nand2_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _12929_/A _23452_/Q _12930_/A vssd1 vssd1 vccd1 vccd1 _12887_/C sky130_fd_sc_hd__and3_1
X_15674_ _15674_/A _15727_/B _15674_/C vssd1 vssd1 vccd1 vccd1 _15814_/A sky130_fd_sc_hd__nand3_4
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17413_ _16408_/A _16741_/A _17425_/A vssd1 vssd1 vccd1 vccd1 _17557_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__18607__B _18947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12358__D _18778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ _11849_/A _16921_/C _11849_/C _19180_/C _12475_/B vssd1 vssd1 vccd1 vccd1
+ _11837_/Y sky130_fd_sc_hd__a32oi_4
X_14625_ _21902_/B _14550_/A _14547_/A _20894_/B vssd1 vssd1 vccd1 vccd1 _14625_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18393_ _18393_/A _18393_/B vssd1 vssd1 vccd1 vccd1 _18414_/C sky130_fd_sc_hd__nand2_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16408__A _16408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17344_ _17179_/A _17170_/B _17220_/X vssd1 vssd1 vccd1 vccd1 _17345_/A sky130_fd_sc_hd__a21o_1
X_14556_ _11604_/X _14544_/X _14548_/X _14555_/X vssd1 vssd1 vccd1 vccd1 _14556_/X
+ sky130_fd_sc_hd__a211o_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11768_ _18805_/A vssd1 vssd1 vccd1 vccd1 _15928_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__12431__A2 _19190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13507_ _13507_/A _13507_/B vssd1 vssd1 vccd1 vccd1 _13507_/Y sky130_fd_sc_hd__nor2_1
X_17275_ _17275_/A _17275_/B vssd1 vssd1 vccd1 vccd1 _17276_/B sky130_fd_sc_hd__nand2_1
X_14487_ _14487_/A _14487_/B _14487_/C vssd1 vssd1 vccd1 vccd1 _14487_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__21968__B _21981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11699_ _11830_/A vssd1 vssd1 vccd1 vccd1 _15699_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19014_ _16437_/A _12103_/X _19210_/A _19191_/A _19013_/X vssd1 vssd1 vccd1 vccd1
+ _19045_/B sky130_fd_sc_hd__o221ai_4
X_13438_ _21883_/A _13810_/B _21883_/C vssd1 vssd1 vccd1 vccd1 _13440_/A sky130_fd_sc_hd__nand3_1
X_16226_ _16661_/A _17148_/A vssd1 vssd1 vccd1 vccd1 _17142_/A sky130_fd_sc_hd__nand2_2
XANTENNA__19647__A1 _19656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19647__B2 _19675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16157_ _16157_/A _16157_/B vssd1 vssd1 vccd1 vccd1 _16157_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__21454__A1 _21455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13369_ _23471_/Q vssd1 vssd1 vccd1 vccd1 _21905_/B sky130_fd_sc_hd__buf_2
XFILLER_182_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11942__A1 _12167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_1024 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15108_ _15120_/B vssd1 vssd1 vccd1 vccd1 _15319_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16088_ _16423_/A _16423_/B vssd1 vssd1 vccd1 vccd1 _16425_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13486__B _13486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18870__A2 _18665_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19916_ _19916_/A _19916_/B _19916_/C _19916_/D vssd1 vssd1 vccd1 vccd1 _20032_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_138_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_728 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15039_ _15208_/A _15075_/B vssd1 vssd1 vccd1 vccd1 _15041_/A sky130_fd_sc_hd__nand2_1
XFILLER_170_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16618__D1 _16027_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22954__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21757__A2 _21906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19847_ _20320_/B _20320_/C _19847_/C vssd1 vssd1 vccd1 vccd1 _19847_/X sky130_fd_sc_hd__and3_1
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16633__A1 _17431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19778_ _19295_/X _19916_/B _19916_/C _19778_/D vssd1 vssd1 vccd1 vccd1 _19783_/A
+ sky130_fd_sc_hd__nand4b_1
XFILLER_3_1034 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22706__B2 _22754_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18729_ _18726_/Y _18727_/X _18728_/Y vssd1 vssd1 vccd1 vccd1 _18910_/A sky130_fd_sc_hd__o21ai_1
XFILLER_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22182__A2 _22560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21740_ _22047_/B _21740_/B vssd1 vssd1 vccd1 vccd1 _22034_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1055 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21671_ _21671_/A _21671_/B vssd1 vssd1 vccd1 vccd1 _21695_/B sky130_fd_sc_hd__nor2_1
XFILLER_178_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23410_ _23442_/CLK _23410_/D vssd1 vssd1 vccd1 vccd1 _23410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20622_ _14615_/X _20504_/A _13014_/Y _20496_/X _20784_/C vssd1 vssd1 vccd1 vccd1
+ _20632_/B sky130_fd_sc_hd__o311a_1
XFILLER_149_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18689__A2 _17643_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23341_ _23343_/CLK _23341_/D vssd1 vssd1 vccd1 vccd1 _23341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20553_ _20553_/A _20553_/B _20553_/C vssd1 vssd1 vccd1 vccd1 _20553_/X sky130_fd_sc_hd__and3_1
XANTENNA__21878__B _22263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23272_ _23559_/CLK _23272_/D vssd1 vssd1 vccd1 vccd1 _23272_/Q sky130_fd_sc_hd__dfxtp_1
X_20484_ _20484_/A _20484_/B _20484_/C vssd1 vssd1 vccd1 vccd1 _20518_/A sky130_fd_sc_hd__nand3_1
XFILLER_193_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12186__A1 _12184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1072 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22223_ _22090_/A _13553_/X _22221_/A _22221_/B vssd1 vssd1 vccd1 vccd1 _22223_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17149__A _17149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22154_ _13415_/X _22164_/A _22388_/C _22051_/X _22032_/Y vssd1 vssd1 vccd1 vccd1
+ _22154_/Y sky130_fd_sc_hd__o32ai_2
XFILLER_172_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16988__A _16988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23198__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16872__A1 _15882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21105_ _21268_/A _12981_/C _20978_/A _21101_/Y _21102_/Y vssd1 vssd1 vccd1 vccd1
+ _21106_/B sky130_fd_sc_hd__a221o_1
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19364__A _19364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22085_ _22086_/A _22086_/B _22093_/C _22093_/D vssd1 vssd1 vccd1 vccd1 _22088_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_99_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22945__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21036_ _21036_/A _21036_/B _21036_/C vssd1 vssd1 vccd1 vccd1 _21279_/C sky130_fd_sc_hd__nand3_2
XFILLER_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11925__A _17626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19811__B _20055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22987_ _22987_/A vssd1 vssd1 vccd1 vccd1 _23325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12740_ _23294_/Q vssd1 vssd1 vccd1 vccd1 _12874_/B sky130_fd_sc_hd__inv_2
XANTENNA__16388__B1 _17450_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21938_ _21938_/A _21938_/B _21939_/A _21939_/B vssd1 vssd1 vccd1 vccd1 _21994_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19530__C _19799_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16927__A2 _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _13177_/B _13177_/C vssd1 vssd1 vccd1 vccd1 _13116_/C sky130_fd_sc_hd__nand2_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21869_ _21824_/A _21824_/C _21813_/X vssd1 vssd1 vccd1 vccd1 _21957_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__19326__B1 _19017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14410_ _14439_/C _14410_/B _14410_/C _14410_/D vssd1 vssd1 vccd1 vccd1 _14410_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11622_ _11918_/A vssd1 vssd1 vccd1 vccd1 _11625_/A sky130_fd_sc_hd__buf_2
XFILLER_169_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15299_/B _15388_/X _15385_/Y _15403_/A vssd1 vssd1 vccd1 vccd1 _15435_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12475__B _12475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ _13933_/A _14263_/Y _14329_/A _14260_/Y vssd1 vssd1 vccd1 vccd1 _14356_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_183_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23539_ _23566_/CLK _23539_/D vssd1 vssd1 vccd1 vccd1 _23539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19539__A _19539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17060_ _17060_/A vssd1 vssd1 vccd1 vccd1 _17761_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14272_ _14269_/Y _14054_/Y _14271_/X vssd1 vssd1 vccd1 vccd1 _14290_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__14166__A2 _14331_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16011_ _15867_/C _15879_/A _15879_/B _16010_/X _16000_/Y vssd1 vssd1 vccd1 vccd1
+ _16011_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_13_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20239__A2 _20237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13223_ _21745_/A vssd1 vssd1 vccd1 vccd1 _13264_/B sky130_fd_sc_hd__buf_2
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13154_ _13114_/X _13116_/Y _13153_/X vssd1 vssd1 vccd1 vccd1 _13168_/D sky130_fd_sc_hd__a21o_1
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23189__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _18445_/A _18447_/B _12105_/C vssd1 vssd1 vccd1 vccd1 _12105_/Y sky130_fd_sc_hd__nand3_4
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17962_ _18211_/A _17752_/X _17959_/Y _17960_/X _18157_/D vssd1 vssd1 vccd1 vccd1
+ _17962_/X sky130_fd_sc_hd__o311a_1
XANTENNA__21379__A1_N _21376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13085_ _13085_/A _13085_/B vssd1 vssd1 vccd1 vccd1 _20595_/C sky130_fd_sc_hd__nor2_1
XFILLER_3_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22936__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19701_ _19701_/A _19701_/B vssd1 vssd1 vccd1 vccd1 _19708_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11816__A1_N _11717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16913_ _16913_/A _16913_/B vssd1 vssd1 vccd1 vccd1 _16934_/C sky130_fd_sc_hd__nand2_1
X_12036_ _12036_/A _12036_/B _16796_/A vssd1 vssd1 vccd1 vccd1 _15707_/A sky130_fd_sc_hd__nand3_1
X_17893_ _17644_/X _17763_/X _17710_/X _17752_/A _17610_/X vssd1 vssd1 vccd1 vccd1
+ _17893_/X sky130_fd_sc_hd__o32a_1
XFILLER_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19632_ _19633_/B _19633_/C _23546_/Q vssd1 vssd1 vccd1 vccd1 _19636_/B sky130_fd_sc_hd__a21boi_1
XFILLER_65_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16844_ _16825_/Y _16823_/Y _16839_/Y _16843_/Y vssd1 vssd1 vccd1 vccd1 _16845_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__13429__A1 _13430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14626__B1 _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19563_ _19588_/A vssd1 vssd1 vccd1 vccd1 _19587_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19014__C1 _19013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16775_ _16435_/C _16755_/Y _17010_/B _17009_/C vssd1 vssd1 vccd1 vccd1 _17008_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13987_ _14396_/A vssd1 vssd1 vccd1 vccd1 _14806_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18514_ _18514_/A _18514_/B _18514_/C vssd1 vssd1 vccd1 vccd1 _18518_/B sky130_fd_sc_hd__nand3_2
XFILLER_20_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ _16593_/A vssd1 vssd1 vccd1 vccd1 _16860_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19494_ _19840_/A _19969_/A _20062_/B _19494_/D vssd1 vssd1 vccd1 vccd1 _19494_/X
+ sky130_fd_sc_hd__and4_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _12709_/X _12936_/X _12945_/A vssd1 vssd1 vccd1 vccd1 _13107_/B sky130_fd_sc_hd__o21ai_2
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18445_ _18445_/A _18445_/B _18972_/A _18447_/B vssd1 vssd1 vccd1 vccd1 _18446_/A
+ sky130_fd_sc_hd__nand4_2
X_15657_ _15656_/X _16658_/B _15713_/B vssd1 vssd1 vccd1 vccd1 _15918_/B sky130_fd_sc_hd__o21ai_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _23295_/Q vssd1 vssd1 vccd1 vccd1 _12875_/B sky130_fd_sc_hd__clkbuf_4
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11570__A _23586_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14608_ _21744_/B _14550_/A _14539_/X _18997_/A _14607_/X vssd1 vssd1 vccd1 vccd1
+ _14608_/X sky130_fd_sc_hd__a221o_1
XFILLER_194_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18376_ _20366_/B _18376_/B _18376_/C _18376_/D vssd1 vssd1 vccd1 vccd1 _18376_/X
+ sky130_fd_sc_hd__or4_1
X_15588_ _15588_/A _15588_/B vssd1 vssd1 vccd1 vccd1 _23502_/D sky130_fd_sc_hd__nor2_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17879__B1 _17747_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17327_ _17327_/A _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17330_/B sky130_fd_sc_hd__nand3_1
XFILLER_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14539_ _23112_/D vssd1 vssd1 vccd1 vccd1 _14539_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17258_ _17267_/A _17267_/B _17267_/C vssd1 vssd1 vccd1 vccd1 _17258_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16209_ _16209_/A _16675_/A vssd1 vssd1 vccd1 vccd1 _16209_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17189_ _17189_/A _17189_/B vssd1 vssd1 vccd1 vccd1 _17189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21978__A2 _21864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16303__B1 _15682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16601__A _17108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22927__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16606__A1 _16604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22910_ _12608_/X input34/X _22918_/S vssd1 vssd1 vccd1 vccd1 _22911_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15217__A _15286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22841_ _22840_/A _22840_/B _22840_/C vssd1 vssd1 vccd1 vccd1 _22842_/A sky130_fd_sc_hd__o21a_1
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14093__A1 _14070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19556__B1 _19554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15290__B1 _15402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19020__A2 _11846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22772_ _22772_/A _22772_/B _22772_/C vssd1 vssd1 vccd1 vccd1 _22774_/B sky130_fd_sc_hd__nor3_1
XFILLER_65_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16909__A2 _16908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17031__A1 _14631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_756 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21723_ _21723_/A _21723_/B _21723_/C _21723_/D vssd1 vssd1 vccd1 vccd1 _21723_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_80_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__23104__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21654_ _21654_/A _21654_/B _23572_/Q vssd1 vssd1 vccd1 vccd1 _21660_/D sky130_fd_sc_hd__nand3_1
XFILLER_184_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20605_ _20605_/A _20605_/B vssd1 vssd1 vccd1 vccd1 _20606_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15887__A _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21585_ _21627_/B _21627_/C _21627_/D vssd1 vssd1 vccd1 vccd1 _21585_/X sky130_fd_sc_hd__and3_1
XFILLER_137_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23324_ _23327_/CLK _23324_/D vssd1 vssd1 vccd1 vccd1 _23324_/Q sky130_fd_sc_hd__dfxtp_2
X_20536_ _20535_/X _20533_/A _20525_/X vssd1 vssd1 vccd1 vccd1 _20542_/A sky130_fd_sc_hd__a21oi_1
XFILLER_137_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15896__A2 _15866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_500 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23255_ _23255_/A vssd1 vssd1 vccd1 vccd1 _23445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20467_ _20907_/A _20906_/A _12876_/A vssd1 vssd1 vccd1 vccd1 _21070_/A sky130_fd_sc_hd__o21a_1
XFILLER_180_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21969__A2 _21981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22206_ _22177_/Y _22195_/Y _22200_/Y _22205_/Y vssd1 vssd1 vccd1 vccd1 _22207_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__12742__C _20639_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18834__A2 _19196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13371__A3 _13802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23186_ _23254_/S vssd1 vssd1 vccd1 vccd1 _23195_/S sky130_fd_sc_hd__clkbuf_2
X_20398_ _18376_/C _20368_/C _20368_/D _20314_/X vssd1 vssd1 vccd1 vccd1 _20428_/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14015__B _14015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22137_ _21884_/B _21996_/Y _21999_/Y vssd1 vssd1 vccd1 vccd1 _22139_/C sky130_fd_sc_hd__o21ai_2
XFILLER_160_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22918__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22068_ _21934_/B _21934_/A _21918_/B _21939_/A _21940_/B vssd1 vssd1 vccd1 vccd1
+ _22208_/C sky130_fd_sc_hd__a32oi_4
XFILLER_102_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_67 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21019_ _21243_/A _21243_/B _21019_/C _21353_/A vssd1 vssd1 vccd1 vccd1 _21029_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_130_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14871__A3 _14621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ _23354_/Q vssd1 vssd1 vccd1 vccd1 _13911_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_58_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14890_ _14890_/A vssd1 vssd1 vccd1 vccd1 _15305_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12882__A2 _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13841_ _13820_/Y _13830_/Y _13834_/Y _13836_/A vssd1 vssd1 vccd1 vccd1 _13843_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_90_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16560_ _16556_/Y _16558_/X _16559_/Y vssd1 vssd1 vccd1 vccd1 _16560_/Y sky130_fd_sc_hd__a21oi_2
X_13772_ _13634_/X _13630_/Y _13768_/Y _13771_/Y _13636_/X vssd1 vssd1 vccd1 vccd1
+ _13772_/X sky130_fd_sc_hd__o2111a_1
XFILLER_74_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15511_ _15508_/X _15509_/Y _15511_/C _15511_/D vssd1 vssd1 vccd1 vccd1 _15513_/D
+ sky130_fd_sc_hd__and4bb_1
XFILLER_128_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12723_ _12723_/A vssd1 vssd1 vccd1 vccd1 _12723_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16491_ _16490_/X _16052_/X _16433_/X _16757_/D vssd1 vssd1 vccd1 vccd1 _16492_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17573__A2 _17565_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18770__A1 _18771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18230_ _18269_/A _18231_/B vssd1 vssd1 vccd1 vccd1 _18236_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15442_ _15439_/B _15442_/B _15442_/C _15442_/D vssd1 vssd1 vccd1 vccd1 _15478_/C
+ sky130_fd_sc_hd__and4b_1
X_12654_ _12654_/A _12723_/A vssd1 vssd1 vccd1 vccd1 _12654_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18507__D1 _19847_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ _11610_/C _11773_/C _11604_/X vssd1 vssd1 vccd1 vccd1 _11611_/A sky130_fd_sc_hd__a21bo_1
XFILLER_88_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18161_ _20271_/A _18161_/B _18161_/C _20217_/A vssd1 vssd1 vccd1 vccd1 _18163_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_156_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17499__A2_N _17155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15373_ _15310_/B _15369_/A _15369_/B _15533_/A _15371_/B vssd1 vssd1 vccd1 vccd1
+ _15373_/X sky130_fd_sc_hd__a32o_1
XFILLER_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12585_ _23301_/Q vssd1 vssd1 vccd1 vccd1 _12683_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__17325__A2 _17323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17112_ _17112_/A _17112_/B vssd1 vssd1 vccd1 vccd1 _17123_/C sky130_fd_sc_hd__nor2_1
XFILLER_12_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14324_ _14324_/A _14324_/B vssd1 vssd1 vccd1 vccd1 _14325_/B sky130_fd_sc_hd__xor2_1
X_18092_ _17974_/C _18947_/C _17567_/X _18093_/A _18172_/C vssd1 vssd1 vccd1 vccd1
+ _18101_/B sky130_fd_sc_hd__a32o_1
XFILLER_117_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23480__CLK _23492_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17043_ _17043_/A vssd1 vssd1 vccd1 vccd1 _18947_/A sky130_fd_sc_hd__clkbuf_4
X_14255_ _14255_/A _14255_/B vssd1 vssd1 vccd1 vccd1 _14324_/B sky130_fd_sc_hd__nand2_1
XFILLER_109_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _20464_/A _20464_/D _20464_/B _20464_/C vssd1 vssd1 vccd1 vccd1 _13208_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_99_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13110__A _21050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14186_ _14133_/B _14121_/Y _14116_/X _14118_/X vssd1 vssd1 vccd1 vccd1 _14187_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_139_1141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _13129_/X _13135_/Y _13136_/Y vssd1 vssd1 vccd1 vccd1 _13143_/A sky130_fd_sc_hd__a21bo_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18994_ _18812_/A _18812_/B _18812_/C _18814_/A vssd1 vssd1 vccd1 vccd1 _18996_/A
+ sky130_fd_sc_hd__o31ai_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22142__B _22142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17945_ _17945_/A _17945_/B vssd1 vssd1 vccd1 vccd1 _17945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13068_ _13131_/A _13179_/A _12833_/B _12836_/B vssd1 vssd1 vccd1 vccd1 _13070_/B
+ sky130_fd_sc_hd__a31oi_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13764__B _13766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21039__A _21174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15682__D _15682_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12019_ _12019_/A vssd1 vssd1 vccd1 vccd1 _15905_/A sky130_fd_sc_hd__buf_2
XANTENNA__21981__B _21981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17876_ _17876_/A _17876_/B vssd1 vssd1 vccd1 vccd1 _17878_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19615_ _19381_/X _19614_/X _19620_/A _19764_/A vssd1 vssd1 vccd1 vccd1 _19615_/X
+ sky130_fd_sc_hd__o211a_1
X_16827_ _15855_/Y _15856_/Y _17061_/A _17060_/A vssd1 vssd1 vccd1 vccd1 _17064_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_94_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18056__B1_N _23530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15811__A2 _16802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19546_ _19560_/B _19560_/C _19560_/A vssd1 vssd1 vccd1 vccd1 _19546_/Y sky130_fd_sc_hd__o21ai_2
X_16758_ _16763_/A _16763_/B _16763_/C vssd1 vssd1 vccd1 vccd1 _16768_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19002__A2 _18440_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1022 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17013__A1 _23520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15709_ _15709_/A _15899_/A vssd1 vssd1 vccd1 vccd1 _15721_/A sky130_fd_sc_hd__nand2_1
XFILLER_181_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19477_ _19477_/A _19477_/B vssd1 vssd1 vccd1 vccd1 _19477_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16689_ _16674_/X _16676_/Y _16682_/Y _16688_/Y vssd1 vssd1 vccd1 vccd1 _16706_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_22_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18428_ _23538_/Q _18431_/B vssd1 vssd1 vccd1 vccd1 _18429_/B sky130_fd_sc_hd__xnor2_1
XFILLER_146_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18359_ _18207_/X _18208_/X _18358_/Y _18320_/Y vssd1 vssd1 vccd1 vccd1 _18403_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_21_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18513__A1 _18435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21370_ _21370_/A vssd1 vssd1 vccd1 vccd1 _21371_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20321_ _20321_/A _20321_/B vssd1 vssd1 vccd1 vccd1 _20322_/B sky130_fd_sc_hd__xnor2_1
XFILLER_162_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15878__A2 _16549_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13658__C _13660_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13020__A _23296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23040_ input40/X _23184_/B input6/X _23040_/D vssd1 vssd1 vccd1 vccd1 _23097_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_66_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20252_ _20252_/A _20252_/B _20252_/C vssd1 vssd1 vccd1 vccd1 _20252_/X sky130_fd_sc_hd__and3_1
Xclkbuf_4_11_0_bq_clk_i clkbuf_3_5_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _23538_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_127_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16827__A1 _15855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13955__A _23502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20183_ _20183_/A _20183_/B vssd1 vssd1 vccd1 vccd1 _20189_/A sky130_fd_sc_hd__xnor2_1
XFILLER_131_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13510__B1 _22388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21891__B _22558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22128__A2 _13599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22824_ _22856_/C _22856_/D _22856_/A vssd1 vssd1 vccd1 vccd1 _22824_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__20139__A1 _19504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22755_ _22716_/D _22392_/A _22392_/B _22756_/D _22756_/A vssd1 vssd1 vccd1 vccd1
+ _22764_/A sky130_fd_sc_hd__a32o_1
XFILLER_53_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16358__A3 _15802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21706_ _23575_/Q vssd1 vssd1 vccd1 vccd1 _21709_/B sky130_fd_sc_hd__inv_2
XFILLER_197_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22686_ _22615_/B _22615_/A _22685_/X vssd1 vssd1 vccd1 vccd1 _22749_/B sky130_fd_sc_hd__o21ai_1
XFILLER_197_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21412__A _23567_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21637_ _21637_/A _21668_/B _21637_/C vssd1 vssd1 vccd1 vccd1 _21695_/A sky130_fd_sc_hd__and3_1
XFILLER_178_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12370_ _12350_/Y _12372_/C _12384_/A _12369_/X vssd1 vssd1 vccd1 vccd1 _12370_/Y
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__15318__A1 _15233_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21568_ _21568_/A _21568_/B vssd1 vssd1 vccd1 vccd1 _21577_/C sky130_fd_sc_hd__nor2_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23307_ _23307_/CLK _23307_/D vssd1 vssd1 vccd1 vccd1 _23307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20519_ _20518_/X _20492_/B _20512_/B vssd1 vssd1 vccd1 vccd1 _20523_/B sky130_fd_sc_hd__a21o_1
XFILLER_197_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21499_ _21548_/B _21548_/D _21595_/C _21546_/A _21434_/X vssd1 vssd1 vccd1 vccd1
+ _21554_/C sky130_fd_sc_hd__a41o_1
XFILLER_5_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_8_0_bq_clk_i_A clkbuf_4_9_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18721__A _18721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14040_ _14026_/X _14121_/A _14039_/Y vssd1 vssd1 vccd1 vccd1 _14063_/A sky130_fd_sc_hd__o21ai_1
XFILLER_107_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23238_ _23238_/A vssd1 vssd1 vccd1 vccd1 _23437_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__22603__A3 _13816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23169_ _23169_/A vssd1 vssd1 vccd1 vccd1 _23178_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_133_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input41_A x[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15991_ _15991_/A vssd1 vssd1 vccd1 vccd1 _17235_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12304__A1 _19082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22367__A2 _13527_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17730_ _17838_/B _17725_/Y _17729_/X vssd1 vssd1 vccd1 vccd1 _17781_/A sky130_fd_sc_hd__a21o_1
XFILLER_121_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14942_ _14943_/B _14966_/B _14943_/A vssd1 vssd1 vccd1 vccd1 _14947_/A sky130_fd_sc_hd__a21o_1
XFILLER_88_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16046__A2 _16315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17661_ _17661_/A _17661_/B _17661_/C vssd1 vssd1 vccd1 vccd1 _17662_/A sky130_fd_sc_hd__nand3_2
XFILLER_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14873_ _14058_/X _14904_/A _14872_/Y vssd1 vssd1 vccd1 vccd1 _14903_/A sky130_fd_sc_hd__o21ai_1
X_19400_ _19390_/X _19393_/Y _19398_/B vssd1 vssd1 vccd1 vccd1 _19400_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_169_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22119__A2 _21994_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16612_ _16612_/A _16612_/B _16612_/C vssd1 vssd1 vccd1 vccd1 _16832_/A sky130_fd_sc_hd__nand3_1
XFILLER_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13824_ _13626_/Y _13627_/Y _13821_/Y _13823_/Y vssd1 vssd1 vccd1 vccd1 _13824_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_29_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17592_ _17592_/A vssd1 vssd1 vccd1 vccd1 _17593_/A sky130_fd_sc_hd__buf_4
XFILLER_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19331_ _19196_/C _19482_/A _19847_/C _19328_/Y _19543_/A vssd1 vssd1 vccd1 vccd1
+ _19332_/C sky130_fd_sc_hd__o2111ai_1
X_16543_ _16530_/A _16530_/B _16530_/C vssd1 vssd1 vccd1 vccd1 _16543_/X sky130_fd_sc_hd__a21o_1
XFILLER_188_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13755_ _13755_/A _13755_/B _13755_/C vssd1 vssd1 vccd1 vccd1 _13755_/Y sky130_fd_sc_hd__nand3_1
XFILLER_189_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19262_ _19262_/A vssd1 vssd1 vccd1 vccd1 _19614_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12706_ _12677_/X _12704_/X _20645_/C _12705_/X vssd1 vssd1 vccd1 vccd1 _12706_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_149_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16474_ _16474_/A _16474_/B vssd1 vssd1 vccd1 vccd1 _16476_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16754__B1 _16778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13686_ _13686_/A vssd1 vssd1 vccd1 vccd1 _13743_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18213_ _20269_/D _17323_/X _17324_/X _18212_/X vssd1 vssd1 vccd1 vccd1 _18214_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__15021__A3 _15195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13568__B1 _21892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15425_ _15424_/B _15424_/C _15424_/A vssd1 vssd1 vccd1 vccd1 _15426_/B sky130_fd_sc_hd__a21oi_1
X_19193_ _19327_/B _19700_/A _19193_/C vssd1 vssd1 vccd1 vccd1 _19195_/A sky130_fd_sc_hd__nand3_1
X_12637_ _13019_/C _20639_/A _13019_/B vssd1 vssd1 vccd1 vccd1 _12637_/X sky130_fd_sc_hd__and3_4
XFILLER_15_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18144_ _18149_/D _18144_/B _18144_/C _18149_/B vssd1 vssd1 vccd1 vccd1 _18144_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_89_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12568_ _12568_/A vssd1 vssd1 vccd1 vccd1 _23519_/D sky130_fd_sc_hd__clkbuf_1
X_15356_ _15356_/A vssd1 vssd1 vccd1 vccd1 _15488_/B sky130_fd_sc_hd__inv_2
XANTENNA__18797__A_N _18799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14307_ _14307_/A vssd1 vssd1 vccd1 vccd1 _14310_/A sky130_fd_sc_hd__clkbuf_1
X_18075_ _18075_/A _18075_/B _18014_/B vssd1 vssd1 vccd1 vccd1 _18114_/B sky130_fd_sc_hd__or3b_1
XFILLER_176_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12499_ _16141_/A _16795_/A vssd1 vssd1 vccd1 vccd1 _17964_/A sky130_fd_sc_hd__nand2_4
X_15287_ _15214_/A _15214_/B _15286_/Y vssd1 vssd1 vccd1 vccd1 _15288_/B sky130_fd_sc_hd__o21ai_4
XFILLER_172_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18631__A _18788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17026_ _16792_/B _17026_/B _17026_/C _17026_/D vssd1 vssd1 vccd1 vccd1 _17026_/Y
+ sky130_fd_sc_hd__nand4b_1
XFILLER_176_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14238_ _14302_/B _14302_/C vssd1 vssd1 vccd1 vccd1 _14294_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16809__A1 _15736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ _14818_/A _14818_/B _14821_/A vssd1 vssd1 vccd1 vccd1 _14227_/A sky130_fd_sc_hd__and3_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19165__C _19165_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23004__A0 _21852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21992__A _21992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _11864_/X _11865_/X _19505_/A _19504_/A _19157_/A vssd1 vssd1 vccd1 vccd1
+ _18978_/B sky130_fd_sc_hd__o221a_2
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _17928_/A _17928_/B vssd1 vssd1 vccd1 vccd1 _17928_/Y sky130_fd_sc_hd__nand2_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19223__A2 _19179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17234__A1 _19494_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17859_ _16684_/X _16683_/X _20055_/C _17766_/C _20055_/D vssd1 vssd1 vccd1 vccd1
+ _17859_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18982__A1 _12130_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20870_ _20872_/A _20872_/B _20872_/C vssd1 vssd1 vccd1 vccd1 _20870_/X sky130_fd_sc_hd__and3_1
XFILLER_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19529_ _19528_/Y _19333_/Y _19340_/A _19345_/C vssd1 vssd1 vccd1 vccd1 _19562_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18734__A1 _19279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22540_ _22730_/B _22540_/B vssd1 vssd1 vccd1 vccd1 _22540_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_718 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22471_ _13470_/X _22754_/B _22465_/Y _22468_/X vssd1 vssd1 vccd1 vccd1 _22475_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_148_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16326__A _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21422_ _21422_/A _21422_/B vssd1 vssd1 vccd1 vccd1 _23547_/D sky130_fd_sc_hd__xor2_1
XFILLER_182_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18498__B1 _18458_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21353_ _21353_/A vssd1 vssd1 vccd1 vccd1 _21576_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18541__A _18541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20304_ _20303_/C _20303_/A _23553_/Q vssd1 vssd1 vccd1 vccd1 _20359_/B sky130_fd_sc_hd__a21o_1
XANTENNA__22046__A1 _21906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_918 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21284_ _21048_/A _21048_/B _20957_/X _20645_/Y vssd1 vssd1 vccd1 vccd1 _21285_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23023_ _23342_/Q input23/X _23023_/S vssd1 vssd1 vccd1 vccd1 _23024_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13685__A _22220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20235_ _20232_/Y _20162_/X _20228_/Y _20231_/Y vssd1 vssd1 vccd1 vccd1 _20235_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_131_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20166_ _20167_/B _20232_/A _20167_/A vssd1 vssd1 vccd1 vccd1 _20229_/A sky130_fd_sc_hd__a21o_1
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11917__B _23590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20097_ _19991_/B _19991_/C _19991_/A _19998_/X vssd1 vssd1 vccd1 vccd1 _20097_/Y
+ sky130_fd_sc_hd__a31oi_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11933__A _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11870_ _16044_/A vssd1 vssd1 vccd1 vccd1 _11871_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22807_ _22803_/X _22802_/Y _22840_/B _22789_/X _22788_/X vssd1 vssd1 vccd1 vccd1
+ _22808_/C sky130_fd_sc_hd__a2111oi_1
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20999_ _20884_/X _20885_/X _20996_/X _20998_/Y vssd1 vssd1 vccd1 vccd1 _20999_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12467__C _18755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13540_ _13540_/A _13540_/B _13540_/C vssd1 vssd1 vccd1 vccd1 _13540_/Y sky130_fd_sc_hd__nand3_1
XFILLER_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22738_ _22738_/A _22738_/B vssd1 vssd1 vccd1 vccd1 _22738_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18435__B _18435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _13471_/A vssd1 vssd1 vccd1 vccd1 _22096_/B sky130_fd_sc_hd__clkbuf_2
X_22669_ _22667_/D _22476_/A _22476_/B _22725_/A _22670_/C vssd1 vssd1 vccd1 vccd1
+ _22671_/C sky130_fd_sc_hd__a32o_1
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16080__A1_N _15889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15210_ _15282_/A _15211_/B _15282_/B vssd1 vssd1 vccd1 vccd1 _15212_/A sky130_fd_sc_hd__a21oi_1
X_12422_ _19512_/C _19530_/D _18511_/A _12422_/D vssd1 vssd1 vccd1 vccd1 _12423_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_173_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16190_ _15604_/X _16658_/C _15921_/B vssd1 vssd1 vccd1 vccd1 _16195_/A sky130_fd_sc_hd__o21ai_1
XFILLER_127_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12353_ _12353_/A vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__buf_2
X_15141_ _15141_/A _15141_/B vssd1 vssd1 vccd1 vccd1 _15144_/B sky130_fd_sc_hd__nand2_2
XANTENNA__19547__A _19547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15072_ _15072_/A _15072_/B vssd1 vssd1 vccd1 vccd1 _23273_/D sky130_fd_sc_hd__nor2_1
XFILLER_181_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12284_ _12282_/X _12283_/Y _15699_/A vssd1 vssd1 vccd1 vccd1 _12284_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_153_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18900_ _18893_/A _18893_/B _18893_/C _18895_/X vssd1 vssd1 vccd1 vccd1 _18900_/X
+ sky130_fd_sc_hd__a31o_1
X_14023_ _14078_/A _14191_/A _14023_/C vssd1 vssd1 vccd1 vccd1 _14086_/B sky130_fd_sc_hd__nand3_2
XFILLER_136_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19880_ _19880_/A _19880_/B _19893_/B vssd1 vssd1 vccd1 vccd1 _19880_/Y sky130_fd_sc_hd__nand3_1
XFILLER_107_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18831_ _18634_/A _18634_/B _18639_/A _18639_/B vssd1 vssd1 vccd1 vccd1 _18831_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_122_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18661__B1 _19011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22123__D _22510_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14203__B _14203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18762_ _18599_/A _18599_/B _18602_/Y vssd1 vssd1 vccd1 vccd1 _18763_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__16121__D _16634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18008__A3 _17324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19205__A2 _17408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15974_ _16856_/A _16856_/B _15974_/C _15974_/D vssd1 vssd1 vccd1 vccd1 _15975_/B
+ sky130_fd_sc_hd__nand4_4
X_17713_ _19670_/A _17635_/A _17625_/Y vssd1 vssd1 vccd1 vccd1 _17714_/A sky130_fd_sc_hd__o21ai_1
XFILLER_48_442 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14925_ _14926_/B _14923_/C _14923_/A vssd1 vssd1 vccd1 vccd1 _14927_/C sky130_fd_sc_hd__a21o_1
X_18693_ _18667_/Y _18672_/Y _18689_/X _18692_/X vssd1 vssd1 vccd1 vccd1 _18751_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_36_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12939__A _20669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17767__A2 _17763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11843__A _11846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17644_ _17644_/A vssd1 vssd1 vccd1 vccd1 _17644_/X sky130_fd_sc_hd__clkbuf_2
X_14856_ _14809_/Y _14810_/X _14811_/X vssd1 vssd1 vccd1 vccd1 _14856_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15242__A3 _15310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13789__B1 _21744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13807_ _21744_/C _13602_/A _13783_/A _13483_/C vssd1 vssd1 vccd1 vccd1 _13809_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_63_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17575_ _17575_/A vssd1 vssd1 vccd1 vccd1 _17575_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14787_ _14788_/A _14857_/A _14788_/C vssd1 vssd1 vccd1 vccd1 _14789_/A sky130_fd_sc_hd__a21o_1
X_11999_ _11999_/A _11999_/B _18814_/A vssd1 vssd1 vccd1 vccd1 _12184_/A sky130_fd_sc_hd__and3_2
XFILLER_189_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19314_ _11822_/X _19499_/A _18656_/Y vssd1 vssd1 vccd1 vccd1 _19314_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16526_ _16526_/A _16526_/B _16526_/C _16526_/D vssd1 vssd1 vccd1 vccd1 _16544_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12461__B1 _12460_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ _13739_/A _13739_/B _13739_/C vssd1 vssd1 vccd1 vccd1 _13738_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19245_ _19245_/A vssd1 vssd1 vccd1 vccd1 _19245_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16457_ _16457_/A _16457_/B _17845_/D _16457_/D vssd1 vssd1 vccd1 vccd1 _16457_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_32_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13005__A2 _20782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13669_ _13680_/C _13673_/A vssd1 vssd1 vccd1 vccd1 _13672_/C sky130_fd_sc_hd__nand2_1
XFILLER_143_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15408_ _15408_/A vssd1 vssd1 vccd1 vccd1 _15511_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_19176_ _19325_/A _19183_/B _19178_/C vssd1 vssd1 vccd1 vccd1 _19176_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__21987__A _21987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16388_ _16054_/X _16055_/X _17450_/C _16309_/A _16309_/B vssd1 vssd1 vccd1 vccd1
+ _16395_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18127_ _18124_/Y _18134_/C _18132_/B vssd1 vssd1 vccd1 vccd1 _18127_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15339_ _15339_/A vssd1 vssd1 vccd1 vccd1 _15528_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18058_ _18058_/A _18139_/B _18139_/C _18058_/D vssd1 vssd1 vccd1 vccd1 _18060_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17009_ _17009_/A _17009_/B _17009_/C vssd1 vssd1 vccd1 vccd1 _17012_/A sky130_fd_sc_hd__nand3_1
XFILLER_132_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20020_ _20017_/X _19904_/X _20015_/X _20016_/Y vssd1 vssd1 vccd1 vccd1 _20113_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_141_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14269__A1 _14068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_995 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14269__B2 _15195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17424__B _19949_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21971_ _22107_/A _21971_/B vssd1 vssd1 vccd1 vccd1 _21973_/C sky130_fd_sc_hd__nand2_1
XFILLER_67_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20922_ _20929_/B vssd1 vssd1 vccd1 vccd1 _20934_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15769__A1 _16447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13229__C1 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20853_ _20853_/A _20853_/B vssd1 vssd1 vccd1 vccd1 _20854_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1059 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13244__A2 _13732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23572_ _23578_/CLK _23572_/D vssd1 vssd1 vccd1 vccd1 _23572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20784_ _20921_/A _20921_/B _20784_/C vssd1 vssd1 vccd1 vccd1 _20790_/B sky130_fd_sc_hd__and3_1
XFILLER_195_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_331 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19380__A1 _18673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19380__B2 _12324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22523_ _22524_/A _22524_/B _22524_/C _22524_/D vssd1 vssd1 vccd1 vccd1 _22523_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_195_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16056__A _17062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22454_ _22454_/A _22454_/B vssd1 vssd1 vccd1 vccd1 _23565_/D sky130_fd_sc_hd__xor2_4
XFILLER_136_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21405_ _21335_/A _21354_/X _21407_/A _21404_/Y vssd1 vssd1 vccd1 vccd1 _21411_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22385_ _22479_/B vssd1 vssd1 vccd1 vccd1 _22641_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__15402__C_N _15442_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22505__B _22505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21336_ _21402_/B _21336_/B vssd1 vssd1 vccd1 vccd1 _21342_/C sky130_fd_sc_hd__nand2_1
XANTENNA__20293__A3 _20242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_884 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21267_ _21207_/C _21270_/A _21267_/C vssd1 vssd1 vccd1 vccd1 _21270_/B sky130_fd_sc_hd__nand3b_1
XFILLER_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23006_ _23334_/Q input14/X _23012_/S vssd1 vssd1 vccd1 vccd1 _23007_/A sky130_fd_sc_hd__mux2_1
X_20218_ _20271_/C _20271_/D _20215_/X vssd1 vssd1 vccd1 vccd1 _20218_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19814__B _20055_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21198_ _21431_/C _21387_/B _21194_/Y _21307_/A vssd1 vssd1 vccd1 vccd1 _21198_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__22521__A _22521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20149_ _20156_/B vssd1 vssd1 vccd1 vccd1 _20158_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _12979_/A _12981_/B _12980_/A _12955_/Y vssd1 vssd1 vccd1 vccd1 _12972_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12759__A _23451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17749__A2 _17980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18946__B2 _17431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_892 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14710_ _23378_/Q _14635_/A _14709_/X vssd1 vssd1 vccd1 vccd1 _14710_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11959_/A _11634_/B _23591_/Q vssd1 vssd1 vccd1 vccd1 _15841_/B sky130_fd_sc_hd__a21o_2
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15690_ _15686_/X _15716_/C _16591_/D vssd1 vssd1 vccd1 vccd1 _15691_/A sky130_fd_sc_hd__o21ai_2
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14396__D _14760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14641_ _23332_/Q vssd1 vssd1 vccd1 vccd1 _22142_/B sky130_fd_sc_hd__buf_2
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _11853_/A vssd1 vssd1 vccd1 vccd1 _14729_/A sky130_fd_sc_hd__buf_2
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17360_ _17036_/X _17200_/A _17200_/C vssd1 vssd1 vccd1 vccd1 _17362_/B sky130_fd_sc_hd__a21boi_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14572_ _23266_/Q _14520_/X _14568_/X _14571_/X vssd1 vssd1 vccd1 vccd1 _14572_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11784_ _11999_/B _18814_/A _11784_/C vssd1 vssd1 vccd1 vccd1 _12145_/A sky130_fd_sc_hd__nand3_2
XANTENNA__20505__A1 _20502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16311_ _16311_/A vssd1 vssd1 vccd1 vccd1 _16311_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11797__A2 _18859_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _13523_/A _22637_/C vssd1 vssd1 vccd1 vccd1 _13525_/C sky130_fd_sc_hd__nand2_1
X_17291_ _17291_/A _17291_/B vssd1 vssd1 vccd1 vccd1 _17292_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15917__D1 _17233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19030_ _19138_/A _19139_/A vssd1 vssd1 vccd1 vccd1 _19033_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16242_ _16242_/A _16242_/B vssd1 vssd1 vccd1 vccd1 _16253_/A sky130_fd_sc_hd__nand2_1
X_13454_ _13552_/A _13313_/X _13446_/A vssd1 vssd1 vccd1 vccd1 _13458_/A sky130_fd_sc_hd__o21ai_1
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12405_ _18811_/B vssd1 vssd1 vccd1 vccd1 _12410_/C sky130_fd_sc_hd__clkbuf_4
X_16173_ _16174_/C _16174_/B _16172_/X _16137_/X vssd1 vssd1 vccd1 vccd1 _16175_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_13385_ _13417_/A vssd1 vssd1 vccd1 vccd1 _22521_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17685__A1 _17535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ _15124_/A _15124_/B vssd1 vssd1 vccd1 vccd1 _15124_/Y sky130_fd_sc_hd__nand2_1
X_12336_ _12336_/A _12336_/B _12336_/C _12336_/D vssd1 vssd1 vccd1 vccd1 _12366_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_154_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15955__D _23592_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22134__C _22521_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19932_ _19932_/A _19932_/B vssd1 vssd1 vccd1 vccd1 _19932_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12267_ _18947_/B vssd1 vssd1 vccd1 vccd1 _12508_/D sky130_fd_sc_hd__clkbuf_2
X_15055_ _15353_/C vssd1 vssd1 vccd1 vccd1 _15408_/A sky130_fd_sc_hd__buf_2
XANTENNA__19426__A2 _19116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__C _21039_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output72_A _14705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14006_ _14006_/A _14835_/A vssd1 vssd1 vccd1 vccd1 _14007_/B sky130_fd_sc_hd__xnor2_1
X_19863_ _19943_/A _19943_/B _19863_/C vssd1 vssd1 vccd1 vccd1 _19864_/C sky130_fd_sc_hd__nand3_1
X_12198_ _12198_/A _12198_/B vssd1 vssd1 vccd1 vccd1 _12203_/A sky130_fd_sc_hd__nand2_2
XFILLER_123_984 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput80 _14572_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[4] sky130_fd_sc_hd__buf_2
Xoutput91 _23265_/Q vssd1 vssd1 vccd1 vccd1 y[3] sky130_fd_sc_hd__buf_2
XFILLER_150_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18814_ _18814_/A _23395_/Q vssd1 vssd1 vccd1 vccd1 _18996_/B sky130_fd_sc_hd__nand2_2
X_19794_ _19625_/B _19772_/Y _19768_/Y vssd1 vssd1 vccd1 vccd1 _19794_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18745_ _18745_/A _18745_/B vssd1 vssd1 vccd1 vccd1 _18746_/A sky130_fd_sc_hd__and2_1
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16660__A2 _16665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15957_ _17963_/A _16800_/D _15957_/C vssd1 vssd1 vccd1 vccd1 _16612_/B sky130_fd_sc_hd__nand3_1
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14908_ _14968_/A _14968_/B _14908_/C _14968_/C vssd1 vssd1 vccd1 vccd1 _14909_/C
+ sky130_fd_sc_hd__nand4_1
X_18676_ _18481_/X _18473_/A _18486_/A _18474_/X vssd1 vssd1 vccd1 vccd1 _18681_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15888_ _15878_/X _15879_/Y _16423_/A vssd1 vssd1 vccd1 vccd1 _15888_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17627_ _17627_/A vssd1 vssd1 vccd1 vccd1 _18000_/A sky130_fd_sc_hd__clkbuf_4
X_14839_ _14236_/B _14826_/X _14824_/X _14830_/A _14235_/A vssd1 vssd1 vccd1 vccd1
+ _14840_/C sky130_fd_sc_hd__o2111ai_1
XANTENNA__17898__C _20164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17260__A _17260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17558_ _17426_/A _17557_/Y _17430_/A _17553_/Y vssd1 vssd1 vccd1 vccd1 _17558_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16509_ _17723_/C vssd1 vssd1 vccd1 vccd1 _18017_/D sky130_fd_sc_hd__buf_2
X_17489_ _17478_/X _17477_/Y _17290_/A _17486_/Y _17488_/X vssd1 vssd1 vccd1 vccd1
+ _17497_/D sky130_fd_sc_hd__o2111ai_4
XANTENNA__21213__C _21218_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19228_ _19188_/A _19188_/B _19188_/C vssd1 vssd1 vccd1 vccd1 _19228_/X sky130_fd_sc_hd__a21o_1
XFILLER_165_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19114__A1 _12167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1019 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19159_ _18984_/B _19309_/A _19158_/Y vssd1 vssd1 vccd1 vccd1 _19162_/A sky130_fd_sc_hd__o21ai_2
XFILLER_11_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18091__A _20133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16604__A _16604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22170_ _13642_/X _22484_/A _22167_/C _22169_/X vssd1 vssd1 vccd1 vccd1 _22170_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_173_884 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21121_ _21121_/A _21121_/B _21121_/C _21554_/D vssd1 vssd1 vccd1 vccd1 _21125_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_133_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21052_ _20934_/B _21176_/C _21184_/A _21040_/B vssd1 vssd1 vccd1 vccd1 _21053_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_119_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20003_ _20003_/A _20003_/B _20003_/C _20003_/D vssd1 vssd1 vccd1 vccd1 _20011_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_99_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11712__A2 _11721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22185__B1 _22142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21954_ _21982_/A _22089_/A _21982_/B vssd1 vssd1 vccd1 vccd1 _21957_/A sky130_fd_sc_hd__nand3b_1
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20905_ _21072_/A _21172_/A _20905_/C _21299_/A vssd1 vssd1 vccd1 vccd1 _20905_/Y
+ sky130_fd_sc_hd__nand4_1
X_21885_ _21791_/Y _21881_/Y _21884_/Y vssd1 vssd1 vccd1 vccd1 _21885_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18266__A _23534_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15611__B1 _15605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _20836_/A vssd1 vssd1 vccd1 vccd1 _20842_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23555_ _23578_/CLK _23555_/D vssd1 vssd1 vccd1 vccd1 _23555_/Q sky130_fd_sc_hd__dfxtp_1
X_20767_ _20765_/A _20765_/B _20763_/A vssd1 vssd1 vccd1 vccd1 _21030_/C sky130_fd_sc_hd__o21ai_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15402__B _15402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22506_ _22281_/X _22371_/X _22372_/X _22366_/Y _22509_/B vssd1 vssd1 vccd1 vccd1
+ _22506_/X sky130_fd_sc_hd__o41a_1
XANTENNA__14717__A2 _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23486_ _23499_/CLK _23498_/Q vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_1
X_20698_ _20624_/X _20631_/X _20636_/X _20653_/Y vssd1 vssd1 vccd1 vccd1 _20699_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_183_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22437_ _22357_/B _22341_/C _22436_/B vssd1 vssd1 vccd1 vccd1 _22538_/B sky130_fd_sc_hd__a21o_1
XFILLER_148_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17116__B1 _17112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21999__B1 _22476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13170_ _13172_/A _13172_/C _13172_/B _13191_/A _13169_/B vssd1 vssd1 vccd1 vccd1
+ _13171_/B sky130_fd_sc_hd__a32o_1
X_22368_ _22564_/A _22564_/B _22569_/B vssd1 vssd1 vccd1 vccd1 _22368_/Y sky130_fd_sc_hd__nand3_2
XFILLER_191_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12121_ _12121_/A _12121_/B vssd1 vssd1 vccd1 vccd1 _18836_/B sky130_fd_sc_hd__nand2_1
XFILLER_151_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21319_ _21319_/A _21319_/B vssd1 vssd1 vccd1 vccd1 _21319_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14034__A _23498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22299_ _22510_/A _22476_/C _22510_/C vssd1 vssd1 vccd1 vccd1 _22300_/B sky130_fd_sc_hd__and3_1
XFILLER_151_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ _12052_/A vssd1 vssd1 vccd1 vccd1 _12311_/A sky130_fd_sc_hd__buf_4
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_835 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13873__A _21971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16860_ _16860_/A _16860_/B _16860_/C _17066_/C vssd1 vssd1 vccd1 vccd1 _16860_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_42_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19263__C _19900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15811_ _12147_/A _16802_/A _15974_/C _12149_/A _15974_/D vssd1 vssd1 vccd1 vccd1
+ _15813_/A sky130_fd_sc_hd__o2111ai_4
XANTENNA__17064__B _17260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16791_ _16988_/A _16983_/B _16983_/C vssd1 vssd1 vccd1 vccd1 _16792_/B sky130_fd_sc_hd__nand3_1
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18530_ _18528_/Y _18529_/Y _18526_/Y _18519_/Y vssd1 vssd1 vccd1 vccd1 _18554_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__22715__A2 _22564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15742_ _15765_/A vssd1 vssd1 vccd1 vccd1 _15742_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12954_ _13041_/B _13181_/B vssd1 vssd1 vccd1 vccd1 _12954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _11913_/A _11905_/B _11905_/C vssd1 vssd1 vccd1 vccd1 _12254_/A sky130_fd_sc_hd__nand3b_2
XFILLER_34_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18461_ _18461_/A _18461_/B _18461_/C vssd1 vssd1 vccd1 vccd1 _18462_/B sky130_fd_sc_hd__nor3_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15673_ _15735_/B vssd1 vssd1 vccd1 vccd1 _15727_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ _12894_/C vssd1 vssd1 vccd1 vccd1 _12899_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23587__CLK _23588_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17412_ _17406_/Y _17407_/Y _17411_/Y vssd1 vssd1 vccd1 vccd1 _17425_/A sky130_fd_sc_hd__o21ai_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18607__C _18607_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14624_ _23298_/Q vssd1 vssd1 vccd1 vccd1 _20894_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_92_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18392_ _18392_/A _18392_/B vssd1 vssd1 vccd1 vccd1 _18393_/B sky130_fd_sc_hd__and2_1
X_11836_ _18600_/C vssd1 vssd1 vccd1 vccd1 _12475_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12416__B1 _18997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18147__A2 _23529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19344__A1 _19218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17350_/C _17350_/D vssd1 vssd1 vccd1 vccd1 _17346_/A sky130_fd_sc_hd__nand2_1
XFILLER_14_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16158__A1 _16066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14555_ input44/X _14549_/X _14550_/X _13226_/X _14554_/X vssd1 vssd1 vccd1 vccd1
+ _14555_/X sky130_fd_sc_hd__a221o_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _16497_/A _12265_/B _12343_/A _11766_/Y vssd1 vssd1 vccd1 vccd1 _11805_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_53_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16127__C _16314_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13506_ _22553_/C _13712_/D _13505_/X _13502_/X vssd1 vssd1 vccd1 vccd1 _13507_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_187_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17274_ _17270_/Y _17273_/Y _17268_/C vssd1 vssd1 vccd1 vccd1 _17276_/A sky130_fd_sc_hd__o21ai_1
X_14486_ _14486_/A _14486_/B _14486_/C vssd1 vssd1 vccd1 vccd1 _14487_/C sky130_fd_sc_hd__nand3_1
X_11698_ _12239_/A _12240_/A vssd1 vssd1 vccd1 vccd1 _11830_/A sky130_fd_sc_hd__nor2_2
XFILLER_174_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21220__B1_N _21215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19013_ _19013_/A vssd1 vssd1 vccd1 vccd1 _19013_/X sky130_fd_sc_hd__clkbuf_4
X_16225_ _16225_/A vssd1 vssd1 vccd1 vccd1 _16225_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13483__A_N _13264_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13437_ _13634_/A _13634_/B _13804_/B vssd1 vssd1 vccd1 vccd1 _13490_/B sky130_fd_sc_hd__and3_1
XANTENNA__12195__A2 _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18855__B1 _18854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16156_ _19363_/C _19363_/D _17057_/A vssd1 vssd1 vccd1 vccd1 _16157_/B sky130_fd_sc_hd__and3_1
XFILLER_115_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13368_ _13349_/X _13365_/Y _13367_/Y vssd1 vssd1 vccd1 vccd1 _13376_/A sky130_fd_sc_hd__o21a_1
XFILLER_6_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11942__A2 _12168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ _15107_/A _15107_/B _15107_/C vssd1 vssd1 vccd1 vccd1 _15188_/A sky130_fd_sc_hd__nand3_2
XFILLER_6_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12319_ _18941_/B vssd1 vssd1 vccd1 vccd1 _19534_/C sky130_fd_sc_hd__buf_2
XFILLER_114_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16087_ _16167_/C _17414_/A _17414_/B _15890_/A _15890_/B vssd1 vssd1 vccd1 vccd1
+ _16423_/B sky130_fd_sc_hd__a32o_1
XFILLER_114_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13299_ _13299_/A vssd1 vssd1 vccd1 vccd1 _13497_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18870__A3 _18666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19915_ _19776_/X _19783_/X _20306_/A _20196_/B vssd1 vssd1 vccd1 vccd1 _19919_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__16881__A2 _16592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ _15208_/A _15075_/B _14926_/C _14926_/A _15037_/Y vssd1 vssd1 vccd1 vccd1
+ _15038_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16618__C1 _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17255__A _19381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19846_ _19846_/A vssd1 vssd1 vccd1 vccd1 _20320_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_95_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19777_ _19916_/A _19916_/B _19916_/C _20031_/A _19776_/X vssd1 vssd1 vccd1 vccd1
+ _19781_/A sky130_fd_sc_hd__a311o_1
X_16989_ _16989_/A _16989_/B vssd1 vssd1 vccd1 vccd1 _16989_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_570 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14644__A1 _23364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18728_ _18728_/A _18728_/B vssd1 vssd1 vccd1 vccd1 _18728_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_743 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18659_ _12187_/Y _18656_/Y _18959_/A vssd1 vssd1 vccd1 vccd1 _18662_/A sky130_fd_sc_hd__o21ai_1
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21670_ _21671_/B _21671_/A vssd1 vssd1 vccd1 vccd1 _21672_/A sky130_fd_sc_hd__and2_1
XFILLER_197_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16318__B _17845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20621_ _20621_/A _20778_/A vssd1 vssd1 vccd1 vccd1 _20793_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17223__A1_N _17077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16149__A1 _16447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21142__A1 _21542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18543__C1 _18524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23340_ _23401_/CLK _23340_/D vssd1 vssd1 vccd1 vccd1 _23340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20552_ _20552_/A vssd1 vssd1 vccd1 vccd1 _20552_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20290__A_N _20237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21878__C _22226_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20782__C _20782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23271_ _23584_/CLK _23271_/D vssd1 vssd1 vccd1 vccd1 _23271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20483_ _20625_/A _20625_/B _13003_/B _20634_/A _21054_/D vssd1 vssd1 vccd1 vccd1
+ _20484_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_121_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12186__A2 _12185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22222_ _22510_/B vssd1 vssd1 vccd1 vccd1 _22670_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17149__B _17631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22153_ _22153_/A vssd1 vssd1 vccd1 vccd1 _22388_/C sky130_fd_sc_hd__buf_2
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21104_ _12640_/X _12637_/X _21490_/B _20966_/A _21103_/X vssd1 vssd1 vccd1 vccd1
+ _21106_/A sky130_fd_sc_hd__o2111ai_4
XANTENNA__16872__A2 _16382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22084_ _22084_/A vssd1 vssd1 vccd1 vccd1 _22093_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_160_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21035_ _21358_/A _21358_/B _21035_/C vssd1 vssd1 vccd1 vccd1 _21037_/A sky130_fd_sc_hd__nand3_1
XFILLER_101_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18613__A3 _17595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16500__C _16536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19811__C _20055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22986_ _13349_/X input36/X _22990_/S vssd1 vssd1 vccd1 vccd1 _22987_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16388__A1 _16054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21937_ _21783_/X _21755_/X _21760_/X vssd1 vssd1 vccd1 vccd1 _21941_/A sky130_fd_sc_hd__a21boi_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19530__D _19530_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16509__A _17723_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18782__C1 _18666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16927__A3 _17391_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11941__A _16591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12618_/A _12915_/A _12668_/X _12794_/A vssd1 vssd1 vccd1 vccd1 _13177_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_151_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21868_ _21826_/X _21834_/Y _21844_/X vssd1 vssd1 vccd1 vccd1 _21965_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__19326__A1 _18440_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12756__B _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11648_/A vssd1 vssd1 vccd1 vccd1 _11918_/A sky130_fd_sc_hd__buf_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20819_ _20819_/A _20819_/B _20819_/C _20819_/D vssd1 vssd1 vccd1 vccd1 _20820_/C
+ sky130_fd_sc_hd__nand4_1
X_21799_ _13466_/A _13765_/X _22564_/C _21792_/Y _13663_/A vssd1 vssd1 vccd1 vccd1
+ _21799_/X sky130_fd_sc_hd__o2111a_1
XFILLER_196_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12475__C _19659_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14340_ _14340_/A _14340_/B vssd1 vssd1 vccd1 vccd1 _14356_/B sky130_fd_sc_hd__nand2_1
XFILLER_196_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23538_ _23538_/CLK _23538_/D vssd1 vssd1 vccd1 vccd1 _23538_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_196_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19539__B _19539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14271_ _14777_/A _14760_/B _14777_/C vssd1 vssd1 vccd1 vccd1 _14271_/X sky130_fd_sc_hd__and3_1
XANTENNA__14166__A3 _14331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23469_ _23571_/CLK _23481_/Q vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__dfxtp_1
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ _16010_/A vssd1 vssd1 vccd1 vccd1 _16010_/X sky130_fd_sc_hd__buf_2
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13222_ _23333_/Q vssd1 vssd1 vccd1 vccd1 _21745_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14571__B1 _14693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16312__A1 _16464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13153_ _12622_/X _12624_/X _12634_/X vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12104_ _18756_/B _16365_/A _15682_/A vssd1 vssd1 vccd1 vccd1 _12104_/X sky130_fd_sc_hd__and3_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ _17958_/A _16742_/A _17859_/Y vssd1 vssd1 vccd1 vccd1 _18157_/D sky130_fd_sc_hd__o21ai_2
XFILLER_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13084_ _13088_/B _13083_/Y _13101_/C vssd1 vssd1 vccd1 vccd1 _20594_/B sky130_fd_sc_hd__o21ai_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19705__D _19966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19700_ _19700_/A _19700_/B _19700_/C _19700_/D vssd1 vssd1 vccd1 vccd1 _19701_/B
+ sky130_fd_sc_hd__nand4_4
X_12035_ _11998_/Y _12008_/X _12049_/B vssd1 vssd1 vccd1 vccd1 _12035_/Y sky130_fd_sc_hd__o21ai_1
X_16912_ _16911_/Y _16900_/B _16900_/A vssd1 vssd1 vccd1 vccd1 _16934_/B sky130_fd_sc_hd__o21ai_2
XFILLER_78_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17892_ _18017_/B _18017_/C _16408_/X _17303_/A vssd1 vssd1 vccd1 vccd1 _17896_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__16076__B1 _16335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19631_ _20120_/A _19924_/A _19295_/X _19448_/Y _19630_/Y vssd1 vssd1 vccd1 vccd1
+ _19633_/C sky130_fd_sc_hd__o221ai_2
X_16843_ _16843_/A _16843_/B vssd1 vssd1 vccd1 vccd1 _16843_/Y sky130_fd_sc_hd__nand2_2
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14626__A1 _14621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15823__B1 _16451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19562_ _19562_/A _19562_/B _19562_/C vssd1 vssd1 vccd1 vccd1 _19588_/A sky130_fd_sc_hd__nand3_1
XFILLER_168_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19014__B1 _19210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16774_ _17010_/C _16774_/B vssd1 vssd1 vccd1 vccd1 _17009_/C sky130_fd_sc_hd__nand2_1
XFILLER_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13986_ _14386_/A vssd1 vssd1 vccd1 vccd1 _14360_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18513_ _18435_/B _11921_/Y _17712_/B _19534_/C _18508_/Y vssd1 vssd1 vccd1 vccd1
+ _18514_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_19_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15725_ _15723_/B _15723_/C _15723_/A vssd1 vssd1 vccd1 vccd1 _15725_/Y sky130_fd_sc_hd__a21oi_4
X_19493_ _19543_/A vssd1 vssd1 vccd1 vccd1 _20061_/A sky130_fd_sc_hd__clkbuf_2
X_12937_ _12627_/X _12654_/A _12604_/Y vssd1 vssd1 vccd1 vccd1 _12945_/A sky130_fd_sc_hd__o21ai_1
XFILLER_74_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11851__A _11851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18444_ _18444_/A vssd1 vssd1 vccd1 vccd1 _18452_/A sky130_fd_sc_hd__clkbuf_4
X_15656_ _15715_/A vssd1 vssd1 vccd1 vccd1 _15656_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12868_ _20528_/A _20528_/B vssd1 vssd1 vccd1 vccd1 _12935_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14607_ input42/X _14549_/A _14547_/A _20481_/B vssd1 vssd1 vccd1 vccd1 _14607_/X
+ sky130_fd_sc_hd__a22o_1
X_18375_ _18376_/B _18376_/C _18376_/D _20366_/B vssd1 vssd1 vccd1 vccd1 _18377_/A
+ sky130_fd_sc_hd__o22a_1
X_11819_ _12297_/B _12287_/C _11818_/Y vssd1 vssd1 vccd1 vccd1 _11913_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__17328__B1 _17155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13062__B1 _13061_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15587_ _15586_/A _15569_/B _23514_/Q vssd1 vssd1 vccd1 vccd1 _15588_/B sky130_fd_sc_hd__a21oi_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _13056_/A vssd1 vssd1 vccd1 vccd1 _20969_/A sky130_fd_sc_hd__buf_2
XFILLER_105_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17326_ _17891_/A _17326_/B _17326_/C _17326_/D vssd1 vssd1 vccd1 vccd1 _17327_/C
+ sky130_fd_sc_hd__nand4_1
X_14538_ _14538_/A _14538_/B _14538_/C _14535_/A vssd1 vssd1 vccd1 vccd1 _23112_/D
+ sky130_fd_sc_hd__nor4b_2
XFILLER_186_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1046 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17257_ _17058_/B _17039_/Y _17252_/A _16625_/X vssd1 vssd1 vccd1 vccd1 _17267_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_105_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14469_ _14835_/C _14472_/D _14469_/C _14469_/D vssd1 vssd1 vccd1 vccd1 _14474_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_146_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16208_ _16032_/A _16033_/A _16865_/A _16866_/A vssd1 vssd1 vccd1 vccd1 _16675_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17188_ _16948_/A _16948_/B _16946_/X vssd1 vssd1 vccd1 vccd1 _17189_/B sky130_fd_sc_hd__a21oi_1
XFILLER_155_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16139_ _16174_/C _16174_/B _16168_/C vssd1 vssd1 vccd1 vccd1 _16139_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16303__A1 _15862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14314__B1 _14207_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16606__A2 _16311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19829_ _19835_/A _19836_/A _19836_/B vssd1 vssd1 vccd1 vccd1 _19830_/A sky130_fd_sc_hd__nand3_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14617__A1 _23582_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14617__B2 _14879_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22840_ _22840_/A _22840_/B _22840_/C vssd1 vssd1 vccd1 vccd1 _22843_/A sky130_fd_sc_hd__or3_1
XFILLER_186_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19556__A1 _19040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13960__B _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22771_ _22789_/A _22789_/B _22770_/C vssd1 vssd1 vccd1 vccd1 _22772_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__18764__C1 _17761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17031__A2 _16668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__A _18756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21722_ _21728_/C _21722_/B vssd1 vssd1 vccd1 vccd1 _21726_/A sky130_fd_sc_hd__and2b_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_768 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21653_ _21654_/A _21654_/B _23572_/Q vssd1 vssd1 vccd1 vccd1 _21660_/B sky130_fd_sc_hd__a21o_1
XFILLER_36_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20604_ _13202_/A _13208_/A _20465_/C vssd1 vssd1 vccd1 vccd1 _20606_/A sky130_fd_sc_hd__o21ai_1
XFILLER_162_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21584_ _21625_/A _21625_/B _21625_/C vssd1 vssd1 vccd1 vccd1 _21627_/D sky130_fd_sc_hd__nand3_1
XFILLER_138_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15887__B _15890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23323_ _23325_/CLK _23323_/D vssd1 vssd1 vccd1 vccd1 _23323_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13688__A _22220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20535_ _12622_/X _12624_/X _13056_/A vssd1 vssd1 vccd1 vccd1 _20535_/X sky130_fd_sc_hd__a21o_1
XFILLER_193_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16064__A _16064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20466_ _13079_/B _13078_/B _13078_/A vssd1 vssd1 vccd1 vccd1 _20551_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__18819__B1 _19505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23254_ _23445_/Q input31/X _23254_/S vssd1 vssd1 vccd1 vccd1 _23255_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22205_ _22215_/A _22215_/B vssd1 vssd1 vccd1 vccd1 _22205_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__19375__A _19568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23185_ _23241_/A vssd1 vssd1 vccd1 vccd1 _23254_/S sky130_fd_sc_hd__buf_2
XANTENNA__22091__A2 _21987_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20397_ _20384_/A _20339_/A _20384_/C vssd1 vssd1 vccd1 vccd1 _20397_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_134_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22136_ _22136_/A _22136_/B _22136_/C _22136_/D vssd1 vssd1 vccd1 vccd1 _22139_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20314__A _20366_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19525__D _19525_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11936__A _11936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22067_ _22061_/Y _22054_/A _22211_/A _22211_/B vssd1 vssd1 vccd1 vccd1 _22208_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__15408__A _15408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21018_ _21018_/A vssd1 vssd1 vccd1 vccd1 _21353_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__21051__B1 _12634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14608__A1 _21744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14608__B2 _18997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13840_ _13646_/B _13646_/C _13646_/A _13655_/A _13671_/C vssd1 vssd1 vccd1 vccd1
+ _13843_/A sky130_fd_sc_hd__a32o_1
XFILLER_63_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13771_ _21880_/A _13659_/Y _13770_/Y vssd1 vssd1 vccd1 vccd1 _13771_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_90_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22969_ _23025_/A vssd1 vssd1 vccd1 vccd1 _23038_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15510_ _15511_/C _15511_/D _15508_/X _15509_/Y vssd1 vssd1 vccd1 vccd1 _15513_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__18157__C _18157_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12722_ _12722_/A vssd1 vssd1 vccd1 vccd1 _12722_/X sky130_fd_sc_hd__buf_2
X_16490_ _16490_/A _17974_/D _17035_/C vssd1 vssd1 vccd1 vccd1 _16490_/X sky130_fd_sc_hd__and3_1
XFILLER_16_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18770__A2 _18966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15441_ _15441_/A _15441_/B vssd1 vssd1 vccd1 vccd1 _23279_/D sky130_fd_sc_hd__nor2_1
X_12653_ _20528_/A _20528_/B _20782_/C vssd1 vssd1 vccd1 vccd1 _12723_/A sky130_fd_sc_hd__nand3_1
XFILLER_169_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18507__C1 _19381_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18160_ _20269_/D _18272_/A _18324_/A _18279_/B _18090_/A vssd1 vssd1 vccd1 vccd1
+ _18182_/B sky130_fd_sc_hd__a41o_1
X_11604_ _11656_/B vssd1 vssd1 vccd1 vccd1 _11604_/X sky130_fd_sc_hd__buf_2
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15372_ _15446_/B vssd1 vssd1 vccd1 vccd1 _15533_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12584_ _23289_/Q vssd1 vssd1 vccd1 vccd1 _12678_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_156_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23510__D input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17325__A3 _17324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17111_ _17118_/B vssd1 vssd1 vccd1 vccd1 _17301_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_157_957 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14323_ _14344_/B _14318_/Y _14319_/Y _14324_/A vssd1 vssd1 vccd1 vccd1 _14420_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_184_743 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18091_ _20133_/B vssd1 vssd1 vccd1 vccd1 _18172_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_144_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17042_ _17039_/Y _17041_/Y _15884_/A _16147_/A vssd1 vssd1 vccd1 vccd1 _17047_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14254_ _14347_/C _14251_/Y _14361_/A _14253_/Y vssd1 vssd1 vccd1 vccd1 _14255_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_143_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13205_ _13205_/A _13205_/B _13205_/C vssd1 vssd1 vccd1 vccd1 _20464_/C sky130_fd_sc_hd__nand3_2
XFILLER_136_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14185_ _14121_/B _14756_/A _15175_/C _14174_/Y _14984_/A vssd1 vssd1 vccd1 vccd1
+ _14187_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_180_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13136_ _13136_/A _13136_/B _13136_/C vssd1 vssd1 vccd1 vccd1 _13136_/Y sky130_fd_sc_hd__nand3_1
XFILLER_180_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18993_ _16032_/X _16033_/X _18439_/X _18440_/X _19805_/A vssd1 vssd1 vccd1 vccd1
+ _18993_/Y sky130_fd_sc_hd__o221ai_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22142__C _22186_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__A _11846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17944_ _17538_/X _17527_/C _17935_/D vssd1 vssd1 vccd1 vccd1 _17944_/Y sky130_fd_sc_hd__o21ai_1
X_13067_ _13062_/X _13065_/Y _13066_/X vssd1 vssd1 vccd1 vccd1 _13077_/A sky130_fd_sc_hd__o21ai_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21039__B _21039_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13764__C _23477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12018_ _15904_/A vssd1 vssd1 vccd1 vccd1 _12018_/X sky130_fd_sc_hd__buf_2
X_17875_ _17874_/Y _17869_/Y _17867_/Y vssd1 vssd1 vccd1 vccd1 _17881_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__21981__C _21981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19614_ _19614_/A _19614_/B _19903_/B vssd1 vssd1 vccd1 vccd1 _19614_/X sky130_fd_sc_hd__and3_1
XFILLER_94_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16826_ _17073_/A _17073_/B _16823_/Y _16825_/Y vssd1 vssd1 vccd1 vccd1 _16836_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19538__A1 _12282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14876__B _14876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19545_ _19363_/Y _19540_/A _19371_/B _19365_/Y vssd1 vssd1 vccd1 vccd1 _19560_/A
+ sky130_fd_sc_hd__a2bb2oi_2
X_16757_ _16757_/A _16757_/B _16757_/C _16757_/D vssd1 vssd1 vccd1 vccd1 _16763_/C
+ sky130_fd_sc_hd__nand4_1
X_13969_ _13965_/X _13966_/X _14797_/A vssd1 vssd1 vccd1 vccd1 _13969_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15708_ _12147_/A _16802_/A _16591_/C _15704_/B _16591_/D vssd1 vssd1 vccd1 vccd1
+ _15899_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_94_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19476_ _19325_/A _19183_/C _19183_/B vssd1 vssd1 vccd1 vccd1 _19476_/Y sky130_fd_sc_hd__a21boi_2
X_16688_ _11766_/B _17230_/A _16693_/A vssd1 vssd1 vccd1 vccd1 _16688_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__20894__A _20894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18427_ _18207_/X _18208_/X _18420_/C vssd1 vssd1 vccd1 vccd1 _18431_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__23098__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _15639_/A _15648_/A _15639_/C vssd1 vssd1 vccd1 vccd1 _16677_/C sky130_fd_sc_hd__nand3_4
XFILLER_179_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18358_ _18394_/A _18394_/B vssd1 vssd1 vccd1 vccd1 _18358_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18513__A2 _11921_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17309_ _16464_/X _17506_/A _17318_/A vssd1 vssd1 vccd1 vccd1 _17313_/A sky130_fd_sc_hd__o21ai_1
XFILLER_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18289_ _18345_/A _18289_/B vssd1 vssd1 vccd1 vccd1 _18349_/B sky130_fd_sc_hd__and2_1
XFILLER_175_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17721__B1 _17029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20320_ _20320_/A _20320_/B _20320_/C vssd1 vssd1 vccd1 vccd1 _20321_/B sky130_fd_sc_hd__and3_1
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15878__A3 _15887_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_832 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20251_ _20120_/X _20205_/X _20307_/A _20250_/Y vssd1 vssd1 vccd1 vccd1 _20255_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_143_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16612__A _16612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20084__A1 _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16827__A2 _15856_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20182_ _20182_/A _20182_/B vssd1 vssd1 vccd1 vccd1 _20183_/B sky130_fd_sc_hd__xnor2_4
XFILLER_131_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17443__A _17443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22823_ _22818_/Y _22819_/Y _22822_/Y vssd1 vssd1 vccd1 vccd1 _22856_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__20139__A2 _19505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13274__B1 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22754_ _22754_/A _22754_/B _22754_/C _22754_/D vssd1 vssd1 vccd1 vccd1 _22756_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_71_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21705_ _21705_/A vssd1 vssd1 vccd1 vccd1 _21705_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__23089__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22685_ _22631_/A _22631_/B _22683_/A _22683_/B vssd1 vssd1 vccd1 vccd1 _22685_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21636_ _21428_/X _21668_/A _21545_/X vssd1 vssd1 vccd1 vccd1 _21637_/A sky130_fd_sc_hd__a21bo_1
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21567_ _21566_/A _21566_/B _21566_/C vssd1 vssd1 vccd1 vccd1 _21568_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__16515__B2 _16370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23306_ _23307_/CLK _23306_/D vssd1 vssd1 vccd1 vccd1 _23306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20518_ _20518_/A vssd1 vssd1 vccd1 vccd1 _20518_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21498_ _21502_/A vssd1 vssd1 vccd1 vccd1 _21595_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20449_ _20449_/A _20449_/B vssd1 vssd1 vccd1 vccd1 _20449_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23237_ _23437_/Q input22/X _23239_/S vssd1 vssd1 vccd1 vccd1 _23238_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23168_ _23168_/A vssd1 vssd1 vccd1 vccd1 _23406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_194 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22119_ _21936_/B _21994_/Y _21995_/Y _22075_/Y _22078_/Y vssd1 vssd1 vccd1 vccd1
+ _22119_/X sky130_fd_sc_hd__o2111a_1
XFILLER_0_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15990_ _15999_/C _15999_/A vssd1 vssd1 vccd1 vccd1 _15990_/Y sky130_fd_sc_hd__nand2_1
X_23099_ _23099_/A vssd1 vssd1 vccd1 vccd1 _23375_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14042__A _23496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12304__A2 _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A wb_dat_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ _14931_/Y _14932_/X _14947_/B vssd1 vssd1 vccd1 vccd1 _14941_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17660_ _17666_/A _17666_/B _17667_/A vssd1 vssd1 vccd1 vccd1 _17661_/C sky130_fd_sc_hd__a21o_1
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14872_ _14097_/X _14115_/Y _14870_/Y _14871_/X vssd1 vssd1 vccd1 vccd1 _14872_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_36_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16611_ _16655_/B _16655_/C vssd1 vssd1 vccd1 vccd1 _16645_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13823_ _13632_/X _13641_/Y _13643_/Y vssd1 vssd1 vccd1 vccd1 _13823_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17591_ _17591_/A vssd1 vssd1 vccd1 vccd1 _17591_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19330_ _17408_/X _19803_/A _19335_/A vssd1 vssd1 vccd1 vccd1 _19332_/A sky130_fd_sc_hd__o21ai_1
X_16542_ _16564_/A _16565_/B vssd1 vssd1 vccd1 vccd1 _16542_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13754_ _13754_/A _13754_/B vssd1 vssd1 vccd1 vccd1 _13754_/Y sky130_fd_sc_hd__nand2_1
XFILLER_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16203__B1 _15932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19261_ _19261_/A _19903_/B _19261_/C vssd1 vssd1 vccd1 vccd1 _19261_/X sky130_fd_sc_hd__and3_1
XFILLER_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12705_ _12851_/C vssd1 vssd1 vccd1 vccd1 _12705_/X sky130_fd_sc_hd__buf_2
X_16473_ _16475_/B _16475_/C vssd1 vssd1 vccd1 vccd1 _16474_/A sky130_fd_sc_hd__nand2_1
X_13685_ _22220_/C vssd1 vssd1 vccd1 vccd1 _22663_/D sky130_fd_sc_hd__buf_2
XANTENNA__16754__B2 _16792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18212_ _18277_/D _20138_/B _20138_/A vssd1 vssd1 vccd1 vccd1 _18212_/X sky130_fd_sc_hd__and3_1
X_15424_ _15424_/A _15424_/B _15424_/C vssd1 vssd1 vccd1 vccd1 _15426_/A sky130_fd_sc_hd__and3_1
XANTENNA__13568__A1 _22474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19192_ _16437_/X _19668_/A _19210_/A _19649_/A vssd1 vssd1 vccd1 vccd1 _19192_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12636_ _12742_/A vssd1 vssd1 vccd1 vccd1 _20639_/A sky130_fd_sc_hd__buf_2
XFILLER_15_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18143_ _18263_/B _18143_/B vssd1 vssd1 vccd1 vccd1 _18262_/C sky130_fd_sc_hd__nor2_2
XFILLER_12_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15355_ _15350_/X _15352_/Y _15354_/Y vssd1 vssd1 vccd1 vccd1 _15383_/A sky130_fd_sc_hd__a21oi_1
X_12567_ _12567_/A _12566_/Y vssd1 vssd1 vccd1 vccd1 _12568_/A sky130_fd_sc_hd__or2b_1
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14306_ _14306_/A _14306_/B _14306_/C vssd1 vssd1 vccd1 vccd1 _14309_/C sky130_fd_sc_hd__nand3_1
XANTENNA__13121__A _13121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18074_ _17838_/B _17838_/C _18036_/A _18036_/B _17838_/A vssd1 vssd1 vccd1 vccd1
+ _18123_/B sky130_fd_sc_hd__a221o_1
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15286_ _15286_/A _15286_/B _15286_/C vssd1 vssd1 vccd1 vccd1 _15286_/Y sky130_fd_sc_hd__nand3_2
XFILLER_184_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ _23591_/Q _23592_/Q vssd1 vssd1 vccd1 vccd1 _16795_/A sky130_fd_sc_hd__nor2_2
XANTENNA__21976__C _21976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17025_ _17025_/A vssd1 vssd1 vccd1 vccd1 _17025_/Y sky130_fd_sc_hd__inv_2
X_14237_ _14230_/A _14156_/B _14156_/C vssd1 vssd1 vccd1 vccd1 _14302_/C sky130_fd_sc_hd__a21o_1
XFILLER_50_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__23252__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15974__C _15974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21799__D1 _13663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16809__A2 _15738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14168_ _14164_/A _14164_/B _14166_/X _14167_/Y vssd1 vssd1 vccd1 vccd1 _14821_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19165__D _20369_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11576__A _23590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19208__B1 _19207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23004__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13119_/A _13119_/B _20663_/C vssd1 vssd1 vccd1 vccd1 _13121_/C sky130_fd_sc_hd__and3_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21992__B _22508_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _14203_/A _14203_/B _13942_/X vssd1 vssd1 vccd1 vccd1 _14099_/X sky130_fd_sc_hd__a21o_1
X_18976_ _18971_/X _18981_/A _18975_/X vssd1 vssd1 vccd1 vccd1 _18978_/A sky130_fd_sc_hd__o21ai_1
XFILLER_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_760 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _17928_/A _17928_/B _17836_/Y _18129_/B vssd1 vssd1 vccd1 vccd1 _17932_/A
+ sky130_fd_sc_hd__a211o_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17234__A2 _17766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17858_ _17591_/X _17593_/X _17766_/B _17595_/X _17766_/C vssd1 vssd1 vccd1 vccd1
+ _17858_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_94_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16442__B1 _11898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18982__A2 _20080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16809_ _15736_/A _15738_/A _17434_/A _17435_/A _17043_/A vssd1 vssd1 vccd1 vccd1
+ _16810_/A sky130_fd_sc_hd__o221ai_4
XFILLER_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17789_ _16523_/A _16523_/B _18211_/C _18163_/B _19862_/A vssd1 vssd1 vccd1 vccd1
+ _17792_/C sky130_fd_sc_hd__o311a_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19528_ _19335_/A _19335_/B _19332_/B vssd1 vssd1 vccd1 vccd1 _19528_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18734__A2 _19280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19459_ _19456_/Y _19459_/B vssd1 vssd1 vccd1 vccd1 _19460_/A sky130_fd_sc_hd__and2b_1
XFILLER_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22470_ _22465_/Y _22468_/X _22469_/X vssd1 vssd1 vccd1 vccd1 _22475_/C sky130_fd_sc_hd__a21bo_1
XFILLER_72_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_888 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16326__B _16326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21421_ _23566_/Q _21349_/B _21420_/Y _21262_/B vssd1 vssd1 vccd1 vccd1 _21422_/B
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_148_743 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__22047__C _22186_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19695__B1 _11670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21352_ _21352_/A _21352_/B vssd1 vssd1 vccd1 vccd1 _23546_/D sky130_fd_sc_hd__xor2_1
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20303_ _20303_/A _23553_/Q _20303_/C vssd1 vssd1 vccd1 vccd1 _20359_/A sky130_fd_sc_hd__nand3_1
XFILLER_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15181__B1 _15301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21283_ _21440_/B _21432_/A _21432_/B _21502_/A _21276_/A vssd1 vssd1 vccd1 vccd1
+ _21285_/B sky130_fd_sc_hd__a32o_1
XFILLER_190_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20234_ _20228_/Y _20231_/Y _20233_/Y vssd1 vssd1 vccd1 vccd1 _20234_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_190_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23022_ _23022_/A vssd1 vssd1 vccd1 vccd1 _23341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_835 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20165_ _20161_/Y _20162_/X _20229_/C vssd1 vssd1 vccd1 vccd1 _20175_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__19653__A _19653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23320__CLK input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20799__A _20799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20096_ _20096_/A _20096_/B _20096_/C vssd1 vssd1 vccd1 vccd1 _20177_/A sky130_fd_sc_hd__nand3_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22510__C _22510_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11933__B _18859_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22806_ _22788_/X _22789_/X _22805_/X vssd1 vssd1 vccd1 vccd1 _22808_/B sky130_fd_sc_hd__o21a_1
XFILLER_77_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ _21000_/A _21000_/B _21132_/A _21131_/B vssd1 vssd1 vccd1 vccd1 _20998_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_129_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12467__D _18755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12470__A1 _18531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22737_ _21854_/A _21854_/B _22813_/A _22687_/Y vssd1 vssd1 vccd1 vccd1 _22738_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_164_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12470__B2 _12463_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ _13470_/A vssd1 vssd1 vccd1 vccd1 _13470_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22668_ _22671_/A _22720_/A _22666_/X _22667_/X vssd1 vssd1 vccd1 vccd1 _22676_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ _12455_/D vssd1 vssd1 vccd1 vccd1 _12422_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_21619_ _23571_/Q vssd1 vssd1 vccd1 vccd1 _21619_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22599_ _22599_/A _22599_/B vssd1 vssd1 vccd1 vccd1 _22599_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__20296__A1 _20183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ _15138_/X _15140_/B _15140_/C vssd1 vssd1 vccd1 vccd1 _15141_/B sky130_fd_sc_hd__nand3b_1
XFILLER_154_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12352_ _11931_/A _11931_/B _12314_/Y _12310_/A _12379_/A vssd1 vssd1 vccd1 vccd1
+ _12355_/A sky130_fd_sc_hd__a221o_1
XFILLER_5_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15071_ _15220_/A _14749_/X _15220_/B vssd1 vssd1 vccd1 vccd1 _15072_/B sky130_fd_sc_hd__a21oi_1
X_12283_ _12282_/B _19156_/C _12282_/A vssd1 vssd1 vccd1 vccd1 _12283_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14022_ _14078_/A _14044_/B _14191_/C _13901_/B vssd1 vssd1 vccd1 vccd1 _14075_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__17067__B _17077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22993__A0 _21744_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18661__A1 _12113_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18830_ _18830_/A _18830_/B _18647_/A vssd1 vssd1 vccd1 vccd1 _18830_/Y sky130_fd_sc_hd__nor3b_4
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_676 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18761_ _18599_/Y _18754_/Y _18758_/Y _18760_/Y vssd1 vssd1 vccd1 vccd1 _18771_/A
+ sky130_fd_sc_hd__o211ai_4
X_15973_ _15855_/Y _15856_/Y _16126_/A _17092_/A vssd1 vssd1 vccd1 vccd1 _16123_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18949__C1 _19261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17712_ _17712_/A _17712_/B _17960_/B _17712_/D vssd1 vssd1 vccd1 vccd1 _17712_/Y
+ sky130_fd_sc_hd__nand4_4
X_14924_ _14966_/A _14927_/B _14922_/Y _14923_/X vssd1 vssd1 vccd1 vccd1 _14943_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18692_ _18880_/A _18773_/A _18784_/C vssd1 vssd1 vccd1 vccd1 _18692_/X sky130_fd_sc_hd__and3_1
XFILLER_76_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17643_ _17643_/A vssd1 vssd1 vccd1 vccd1 _17643_/X sky130_fd_sc_hd__clkbuf_4
X_14855_ _14855_/A _14855_/B vssd1 vssd1 vccd1 vccd1 _14855_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__21036__C _21036_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13806_ _13616_/B _21916_/A _13805_/Y vssd1 vssd1 vccd1 vccd1 _13812_/B sky130_fd_sc_hd__o21ai_1
X_17574_ _17446_/B _17580_/A _17437_/X _17433_/X vssd1 vssd1 vccd1 vccd1 _17578_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_14786_ _14782_/Y _14783_/X _14789_/C vssd1 vssd1 vccd1 vccd1 _14814_/A sky130_fd_sc_hd__o21bai_2
X_11998_ _12166_/A _11996_/Y _11997_/X vssd1 vssd1 vccd1 vccd1 _11998_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16525_ _16526_/B _16526_/D _16526_/A _17248_/C vssd1 vssd1 vccd1 vccd1 _16528_/A
+ sky130_fd_sc_hd__a22o_1
X_19313_ _19304_/X _19307_/Y _19309_/Y _19312_/Y _19158_/Y vssd1 vssd1 vccd1 vccd1
+ _19321_/A sky130_fd_sc_hd__o2111ai_4
X_13737_ _13735_/X _13705_/D _13585_/A _13736_/X vssd1 vssd1 vccd1 vccd1 _13739_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12461__A1 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15969__C _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22148__B _22270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19244_ _19244_/A _19244_/B _19244_/C vssd1 vssd1 vccd1 vccd1 _19245_/A sky130_fd_sc_hd__nand3_1
X_16456_ _17259_/A vssd1 vssd1 vccd1 vccd1 _17845_/D sky130_fd_sc_hd__clkbuf_4
X_13668_ _13668_/A _13668_/B vssd1 vssd1 vccd1 vccd1 _13673_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15935__C1 _16372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19126__C1 _18607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15407_ _15383_/A _15406_/X _15383_/C vssd1 vssd1 vccd1 vccd1 _15430_/A sky130_fd_sc_hd__a21o_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19175_ _18993_/Y _19173_/X _19182_/B vssd1 vssd1 vccd1 vccd1 _19178_/C sky130_fd_sc_hd__o21bai_1
XFILLER_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12213__A1 _12093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ _20493_/D vssd1 vssd1 vccd1 vccd1 _12915_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16387_ _16462_/B _16443_/C _16309_/A _16309_/B vssd1 vssd1 vccd1 vccd1 _16395_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21987__B _21987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ _13599_/A vssd1 vssd1 vccd1 vccd1 _13599_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_185_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18126_ _18126_/A vssd1 vssd1 vccd1 vccd1 _18134_/C sky130_fd_sc_hd__clkbuf_2
X_15338_ _15338_/A _23506_/Q vssd1 vssd1 vccd1 vccd1 _15339_/A sky130_fd_sc_hd__xnor2_1
XFILLER_118_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15985__B _15985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22164__A _22164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18057_ _18058_/D _18072_/D _18072_/C _18058_/A _18154_/A vssd1 vssd1 vccd1 vccd1
+ _18057_/Y sky130_fd_sc_hd__a41oi_2
XANTENNA__19429__B1 _19116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15269_ _15270_/B _15326_/A _15270_/A vssd1 vssd1 vccd1 vccd1 _15271_/A sky130_fd_sc_hd__a21o_1
XFILLER_172_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17008_ _17008_/A _17008_/B _17008_/C _17011_/A vssd1 vssd1 vccd1 vccd1 _17008_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_104_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22984__A0 _13379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14269__A2 _14069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16663__B1 _16194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18959_ _18959_/A _18959_/B _18959_/C vssd1 vssd1 vccd1 vccd1 _18959_/Y sky130_fd_sc_hd__nand3_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21970_ _21970_/A _21981_/B vssd1 vssd1 vccd1 vccd1 _22107_/C sky130_fd_sc_hd__nand2_1
XANTENNA__17424__C _17959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20921_ _20921_/A _20921_/B _21036_/C vssd1 vssd1 vccd1 vccd1 _20929_/B sky130_fd_sc_hd__nand3_1
XANTENNA__15225__B _15225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15769__A2 _15766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20852_ _20840_/A _20845_/A _20849_/B vssd1 vssd1 vccd1 vccd1 _20856_/A sky130_fd_sc_hd__a21o_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13244__A3 _13732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23571_ _23571_/CLK _23571_/D vssd1 vssd1 vccd1 vccd1 _23571_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12865__A _21039_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20783_ _20783_/A _20783_/B vssd1 vssd1 vccd1 vccd1 _20783_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19380__A2 _17846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22522_ _22517_/Y _22521_/X _22609_/A _22607_/A _22419_/Y vssd1 vssd1 vccd1 vccd1
+ _22524_/D sky130_fd_sc_hd__o2111ai_2
XFILLER_195_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19648__A _19648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22453_ _22451_/Y _22452_/Y _22354_/A vssd1 vssd1 vccd1 vccd1 _22454_/B sky130_fd_sc_hd__a21oi_4
XFILLER_157_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21404_ _21404_/A _21404_/B vssd1 vssd1 vccd1 vccd1 _21404_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17143__A1 _16908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22384_ _22384_/A vssd1 vssd1 vccd1 vccd1 _22567_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21335_ _21335_/A vssd1 vssd1 vccd1 vccd1 _21336_/B sky130_fd_sc_hd__inv_2
XANTENNA__15154__B1 _15488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21266_ _21082_/B _21083_/B _21161_/Y _21265_/Y vssd1 vssd1 vccd1 vccd1 _21266_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__22975__A0 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23005_ _23005_/A vssd1 vssd1 vccd1 vccd1 _23333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20217_ _20217_/A _20217_/B _20269_/C _20217_/D vssd1 vssd1 vccd1 vccd1 _20271_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_132_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21197_ _21365_/A _21299_/A _21358_/C _21295_/B vssd1 vssd1 vccd1 vccd1 _21307_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19814__C _20055_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22521__B _22861_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20148_ _20148_/A _20148_/B _20148_/C vssd1 vssd1 vccd1 vccd1 _20156_/B sky130_fd_sc_hd__nand3_1
XFILLER_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20079_ _20079_/A vssd1 vssd1 vccd1 vccd1 _20164_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1080 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12970_ _20663_/D vssd1 vssd1 vccd1 vccd1 _12979_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18946__A2 _17975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _11947_/A _23256_/B vssd1 vssd1 vccd1 vccd1 _11921_/Y sky130_fd_sc_hd__nand2_4
XFILLER_58_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12478__C _12478_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17631__A _17631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14640_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_1127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _11852_/A vssd1 vssd1 vccd1 vccd1 _12378_/B sky130_fd_sc_hd__buf_2
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19356__C1 _17567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14571_ _13264_/C _14550_/X _14693_/A _11784_/C _14570_/X vssd1 vssd1 vccd1 vccd1
+ _14571_/X sky130_fd_sc_hd__a221o_1
XANTENNA__22871__B1_N _22878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _11977_/B vssd1 vssd1 vccd1 vccd1 _11784_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__20505__A2 _20504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16310_ _16310_/A _16310_/B vssd1 vssd1 vccd1 vccd1 _16313_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13522_ _22562_/B vssd1 vssd1 vccd1 vccd1 _22637_/C sky130_fd_sc_hd__buf_2
XFILLER_158_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17290_ _17290_/A _17297_/D vssd1 vssd1 vccd1 vccd1 _17292_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16241_ _16251_/A _16281_/B _16251_/D _16240_/Y vssd1 vssd1 vccd1 vccd1 _16243_/A
+ sky130_fd_sc_hd__a31o_1
X_13453_ _13453_/A vssd1 vssd1 vccd1 vccd1 _13552_/A sky130_fd_sc_hd__buf_2
XFILLER_186_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ _23390_/Q _23391_/Q vssd1 vssd1 vccd1 vccd1 _18811_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16172_ _16172_/A _17445_/A _17235_/A vssd1 vssd1 vccd1 vccd1 _16172_/X sky130_fd_sc_hd__and3_1
X_13384_ _13304_/X _13308_/Y _21902_/C _13379_/X vssd1 vssd1 vccd1 vccd1 _13417_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_166_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15123_ _15163_/A _15188_/A _15164_/A _15164_/B vssd1 vssd1 vccd1 vccd1 _15188_/B
+ sky130_fd_sc_hd__nand4_1
X_12335_ _12339_/A _12339_/B _12335_/C _12335_/D vssd1 vssd1 vccd1 vccd1 _12336_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15145__B1 _15286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19931_ _19625_/A _19625_/D _19626_/X vssd1 vssd1 vccd1 vccd1 _19931_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15054_ _15054_/A vssd1 vssd1 vccd1 vccd1 _15353_/C sky130_fd_sc_hd__clkbuf_2
X_12266_ _12273_/B _12273_/C _12273_/D _12273_/A vssd1 vssd1 vccd1 vccd1 _12266_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__21769__A1 _13465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14005_ _14005_/A _14005_/B vssd1 vssd1 vccd1 vccd1 _14835_/A sky130_fd_sc_hd__nand2_1
X_19862_ _19862_/A _19862_/B _19862_/C vssd1 vssd1 vccd1 vccd1 _19864_/B sky130_fd_sc_hd__and3_1
X_12197_ _12199_/C _12199_/D vssd1 vssd1 vccd1 vccd1 _12198_/B sky130_fd_sc_hd__nand2_2
XFILLER_122_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput70 _14697_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_123_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput81 _14579_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[5] sky130_fd_sc_hd__buf_2
Xoutput92 _23266_/Q vssd1 vssd1 vccd1 vccd1 y[4] sky130_fd_sc_hd__buf_2
XANTENNA_output65_A _14556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18813_ _18813_/A vssd1 vssd1 vccd1 vccd1 _19505_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19793_ _19793_/A vssd1 vssd1 vccd1 vccd1 _20306_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18744_ _19288_/A _18747_/B _18747_/A vssd1 vssd1 vccd1 vccd1 _18745_/B sky130_fd_sc_hd__a21o_1
X_15956_ _15956_/A _16802_/B _15956_/C _16795_/C vssd1 vssd1 vccd1 vccd1 _17963_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_95_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14230__A _14230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17328__A2_N _17152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18937__A2 _18604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ _14788_/A _14788_/C _14857_/A vssd1 vssd1 vccd1 vccd1 _14909_/B sky130_fd_sc_hd__a21boi_1
X_18675_ _18675_/A _18675_/B _18675_/C vssd1 vssd1 vccd1 vccd1 _18675_/X sky130_fd_sc_hd__or3_1
X_15887_ _15890_/A _15890_/B _15887_/C vssd1 vssd1 vccd1 vccd1 _16423_/A sky130_fd_sc_hd__nand3_2
XANTENNA__20886__B _21124_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17626_ _17626_/A vssd1 vssd1 vccd1 vccd1 _17627_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14838_ _14831_/B _14831_/C _14831_/A vssd1 vssd1 vccd1 vccd1 _14840_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23143__A0 _19156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17898__D _17898_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12434__A1 _12121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17557_ _17557_/A _17557_/B vssd1 vssd1 vccd1 vccd1 _17557_/Y sky130_fd_sc_hd__nand2_1
X_14769_ _15112_/C _13948_/X _14879_/A _15112_/D vssd1 vssd1 vccd1 vccd1 _14774_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ _16530_/A _16558_/A vssd1 vssd1 vccd1 vccd1 _16512_/A sky130_fd_sc_hd__nor2_1
X_17488_ _17481_/C _17481_/D _17487_/Y vssd1 vssd1 vccd1 vccd1 _17488_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19227_ _19256_/A _19256_/C vssd1 vssd1 vccd1 vccd1 _19227_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16439_ _11882_/X _11883_/X _16064_/A vssd1 vssd1 vccd1 vccd1 _16523_/D sky130_fd_sc_hd__a21o_2
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18372__A _23536_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19114__A2 _12168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_724 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19158_ _19158_/A _19304_/A vssd1 vssd1 vccd1 vccd1 _19158_/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18109_ _18110_/B _18110_/A vssd1 vssd1 vccd1 vccd1 _18109_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19089_ _19089_/A _19089_/B vssd1 vssd1 vccd1 vccd1 _19090_/D sky130_fd_sc_hd__nand2_1
XFILLER_145_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21120_ _21387_/C vssd1 vssd1 vccd1 vccd1 _21514_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21051_ _21184_/A _21179_/A _12634_/X _21043_/A vssd1 vssd1 vccd1 vccd1 _21053_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_87_803 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20432__A1 _20411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20002_ _19883_/Y _19884_/X _19888_/D vssd1 vssd1 vccd1 vccd1 _20003_/B sky130_fd_sc_hd__o21ai_1
XFILLER_101_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20142__A _20142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11764__A _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22724__A3 _22664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21953_ _21957_/B _21953_/B _21953_/C vssd1 vssd1 vccd1 vccd1 _21964_/A sky130_fd_sc_hd__nand3b_2
XFILLER_27_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ _21054_/D vssd1 vssd1 vccd1 vccd1 _21299_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21884_ _21884_/A _21884_/B vssd1 vssd1 vccd1 vccd1 _21884_/Y sky130_fd_sc_hd__nand2_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23134__A0 _12100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20835_ _20690_/A _20711_/A _20654_/X _20668_/Y vssd1 vssd1 vccd1 vccd1 _20839_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__16067__A _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23554_ _23578_/CLK _23554_/D vssd1 vssd1 vccd1 vccd1 _23554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20766_ _20766_/A _20766_/B vssd1 vssd1 vccd1 vccd1 _23541_/D sky130_fd_sc_hd__xnor2_1
XFILLER_126_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22505_ _22509_/A _22505_/B _22509_/B vssd1 vssd1 vccd1 vccd1 _22505_/X sky130_fd_sc_hd__and3_1
XANTENNA__19378__A _19534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23485_ _23499_/CLK _23497_/Q vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20697_ _20654_/X _20668_/Y _20718_/B _20715_/C vssd1 vssd1 vccd1 vccd1 _20697_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_7_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22436_ _22436_/A _22436_/B vssd1 vssd1 vccd1 vccd1 _22538_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17116__A1 _19494_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11939__A _12207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22367_ _22284_/Y _13527_/X _22479_/A _22279_/Y vssd1 vssd1 vccd1 vccd1 _22370_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ _11999_/B _18812_/B _11773_/C _12099_/D vssd1 vssd1 vccd1 vccd1 _18836_/A
+ sky130_fd_sc_hd__o211ai_2
X_21318_ _21317_/A _21317_/B _21317_/C _21317_/D vssd1 vssd1 vccd1 vccd1 _21318_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22298_ _22122_/Y _22362_/A _22297_/Y vssd1 vssd1 vccd1 vccd1 _22300_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18616__A1 _12090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17626__A _17626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12051_ _12051_/A vssd1 vssd1 vccd1 vccd1 _12052_/A sky130_fd_sc_hd__buf_4
XFILLER_85_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21249_ _21245_/X _21248_/Y _23565_/Q vssd1 vssd1 vccd1 vccd1 _21249_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16530__A _16530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20959__C1 _12692_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_847 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18092__A2 _18947_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11674__A _23397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15810_ _16019_/A _16019_/B vssd1 vssd1 vccd1 vccd1 _15810_/X sky130_fd_sc_hd__and2_1
X_16790_ _16585_/Y _16587_/Y _16744_/Y _16750_/Y vssd1 vssd1 vccd1 vccd1 _16983_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__16995__B1_N _23523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15850__A1 _18675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22715__A3 _22564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15741_ _16798_/B _14553_/X _15727_/B _15677_/Y vssd1 vssd1 vccd1 vccd1 _15765_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19041__A1 _19040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _13157_/B vssd1 vssd1 vccd1 vccd1 _13181_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _11912_/C _11912_/D _11903_/A vssd1 vssd1 vccd1 vccd1 _11905_/C sky130_fd_sc_hd__a21o_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ _15712_/A _16187_/B _15672_/C vssd1 vssd1 vccd1 vccd1 _15674_/A sky130_fd_sc_hd__nand3_1
X_18460_ _18460_/A vssd1 vssd1 vccd1 vccd1 _18461_/C sky130_fd_sc_hd__buf_2
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12884_ _20669_/A _12884_/B _20908_/A _20801_/C vssd1 vssd1 vccd1 vccd1 _12894_/C
+ sky130_fd_sc_hd__nand4_2
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23513__D input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17411_ _17408_/X _17644_/A _17410_/Y vssd1 vssd1 vccd1 vccd1 _17411_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _23330_/Q vssd1 vssd1 vccd1 vccd1 _21902_/B sky130_fd_sc_hd__buf_2
XFILLER_33_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18391_ _18356_/A _18356_/B _18355_/A vssd1 vssd1 vccd1 vccd1 _18393_/A sky130_fd_sc_hd__a21o_1
X_11835_ _18597_/B vssd1 vssd1 vccd1 vccd1 _18600_/C sky130_fd_sc_hd__clkbuf_4
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12416__A1 _12410_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19344__A2 _17643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17342_ _17220_/X _17179_/X _17350_/C _17350_/D vssd1 vssd1 vccd1 vccd1 _17347_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_53_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14554_ _23263_/Q _14551_/X _14698_/A _14553_/X vssd1 vssd1 vccd1 vccd1 _14554_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16158__A2 _17565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11766_ _11766_/A _11766_/B _11766_/C vssd1 vssd1 vccd1 vccd1 _11766_/Y sky130_fd_sc_hd__nor3_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13505_ _13498_/A _13498_/B _13450_/Y _13495_/X vssd1 vssd1 vccd1 vccd1 _13505_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_159_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17273_ _17039_/Y _17048_/Y _17271_/X _17272_/Y vssd1 vssd1 vccd1 vccd1 _17273_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__16127__D _16314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14485_ _14441_/Y _14445_/Y _14468_/A _14453_/Y vssd1 vssd1 vccd1 vccd1 _14487_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_187_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11697_ _11649_/X _11721_/A _11647_/B vssd1 vssd1 vccd1 vccd1 _12240_/A sky130_fd_sc_hd__a21oi_1
XFILLER_186_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19012_ _19012_/A _19012_/B vssd1 vssd1 vccd1 vccd1 _19045_/A sky130_fd_sc_hd__nand2_1
X_16224_ _16242_/A vssd1 vssd1 vccd1 vccd1 _16246_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13436_ _13474_/A _13474_/B _13460_/D _13460_/A vssd1 vssd1 vccd1 vccd1 _13461_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16155_ _15971_/X _16598_/B _16590_/A vssd1 vssd1 vccd1 vccd1 _16157_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11849__A _11849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22145__C _22145_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13367_ _13348_/X _13366_/Y _13416_/A vssd1 vssd1 vccd1 vccd1 _13367_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_170_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _15107_/B _15107_/C _15107_/A vssd1 vssd1 vccd1 vccd1 _15163_/A sky130_fd_sc_hd__a21o_1
XFILLER_170_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12318_ _12318_/A vssd1 vssd1 vccd1 vccd1 _12381_/C sky130_fd_sc_hd__clkbuf_1
X_16086_ _19363_/D vssd1 vssd1 vccd1 vccd1 _17414_/B sky130_fd_sc_hd__buf_4
XFILLER_142_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13298_ _22569_/B vssd1 vssd1 vccd1 vccd1 _22558_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19914_ _19925_/A _19925_/B vssd1 vssd1 vccd1 vccd1 _20196_/B sky130_fd_sc_hd__and2_1
X_15037_ _14918_/C _14918_/B _14918_/A vssd1 vssd1 vccd1 vccd1 _15037_/Y sky130_fd_sc_hd__a21oi_1
X_12249_ _12246_/Y _12247_/Y _16372_/A _18945_/C _19180_/C vssd1 vssd1 vccd1 vccd1
+ _12271_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_142_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18083__A2 _18219_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19845_ _19504_/X _19505_/X _17406_/B _17406_/A _20369_/B vssd1 vssd1 vccd1 vccd1
+ _20079_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_123_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19776_ _19640_/Y _19768_/Y _19775_/Y vssd1 vssd1 vccd1 vccd1 _19776_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_988 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16988_ _16988_/A vssd1 vssd1 vccd1 vccd1 _16988_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18727_ _18722_/Y _18723_/Y _18914_/B _18914_/A vssd1 vssd1 vccd1 vccd1 _18727_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19032__A1 _18854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12655__A1 _12634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15939_ _16251_/A _16237_/A _16281_/B _16251_/D vssd1 vssd1 vccd1 vccd1 _15948_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23531__CLK _23538_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18658_ _11848_/X _18645_/A _18657_/Y vssd1 vssd1 vccd1 vccd1 _18959_/A sky130_fd_sc_hd__o21ai_4
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17609_ _17609_/A _17609_/B _17770_/A _17770_/B vssd1 vssd1 vccd1 vccd1 _17616_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18589_ _18589_/A _18589_/B _23540_/Q vssd1 vssd1 vccd1 vccd1 _18589_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_3_2_0_bq_clk_i_A clkbuf_3_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13304__A _23323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20620_ _20628_/A _20620_/B _20620_/C vssd1 vssd1 vccd1 vccd1 _20778_/A sky130_fd_sc_hd__nand3_2
XANTENNA__12958__A2 _13151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13080__A1 _12906_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16149__A2 _15766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19198__A _19703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20551_ _20551_/A _20551_/B _20551_/C vssd1 vssd1 vccd1 vccd1 _20579_/A sky130_fd_sc_hd__nand3_1
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23270_ _23492_/CLK _23270_/D vssd1 vssd1 vccd1 vccd1 _23270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20482_ _20482_/A _20482_/B vssd1 vssd1 vccd1 vccd1 _21054_/D sky130_fd_sc_hd__nand2_2
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22221_ _22221_/A _22221_/B vssd1 vssd1 vccd1 vccd1 _22226_/B sky130_fd_sc_hd__nor2_2
XFILLER_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14580__A1 _23268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14580__B2 _12712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_811 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17149__C _17712_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22152_ _22562_/C _22562_/A vssd1 vssd1 vccd1 vccd1 _22164_/A sky130_fd_sc_hd__nand2_2
XFILLER_145_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21103_ _20978_/A _21101_/Y _21102_/Y vssd1 vssd1 vccd1 vccd1 _21103_/X sky130_fd_sc_hd__a21o_1
XFILLER_160_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22083_ _22083_/A _22083_/B _22083_/C vssd1 vssd1 vccd1 vccd1 _22084_/A sky130_fd_sc_hd__nand3_1
XFILLER_154_49 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16609__B1 _17235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21034_ _21281_/A _21282_/A _21050_/C vssd1 vssd1 vccd1 vccd1 _21176_/C sky130_fd_sc_hd__nand3_2
XANTENNA__11697__A2 _11721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20956__A2 _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22985_ _22985_/A vssd1 vssd1 vccd1 vccd1 _23324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12102__B _19193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1086 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21936_ _21936_/A _21936_/B _21936_/C vssd1 vssd1 vccd1 vccd1 _21936_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__16388__A2 _16055_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18782__B1 _18665_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21867_ _21867_/A _21867_/B vssd1 vssd1 vccd1 vccd1 _23560_/D sky130_fd_sc_hd__nor2_1
XFILLER_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19326__A2 _18439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11815_/A vssd1 vssd1 vccd1 vccd1 _12281_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20818_ _20653_/Y _20636_/X _20631_/X _20624_/X vssd1 vssd1 vccd1 vccd1 _20820_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21798_ _21794_/Y _21798_/B _21798_/C vssd1 vssd1 vccd1 vccd1 _21801_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__21431__A _21431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23537_ _23538_/CLK _23537_/D vssd1 vssd1 vccd1 vccd1 _23537_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12475__D _18531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20749_ _20752_/B vssd1 vssd1 vccd1 vccd1 _21157_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_184_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19539__C _19700_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13359__C1 _23326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14270_ _14312_/B vssd1 vssd1 vccd1 vccd1 _14777_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23468_ _23571_/CLK _23480_/Q vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__20047__A _20047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13221_ _13221_/A vssd1 vssd1 vccd1 vccd1 _13732_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14571__A1 _13264_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22419_ _22754_/A _13599_/X _22405_/A _22418_/X vssd1 vssd1 vccd1 vccd1 _22419_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14571__B2 _11784_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23399_ _23432_/CLK _23399_/D vssd1 vssd1 vccd1 vccd1 _23399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16848__B1 _19703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13152_ _12766_/X _12709_/X _13116_/Y _13114_/X vssd1 vssd1 vccd1 vccd1 _13168_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_124_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16312__A2 _16311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ _12424_/A vssd1 vssd1 vccd1 vccd1 _12103_/X sky130_fd_sc_hd__buf_4
X_17960_ _17960_/A _17960_/B _18016_/D vssd1 vssd1 vccd1 vccd1 _17960_/X sky130_fd_sc_hd__and3_1
X_13083_ _12908_/B _12908_/C _12908_/A vssd1 vssd1 vccd1 vccd1 _13083_/Y sky130_fd_sc_hd__a21oi_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__23508__D input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ _12015_/Y _12027_/Y _12033_/Y vssd1 vssd1 vccd1 vccd1 _12049_/B sky130_fd_sc_hd__o21ai_1
X_16911_ _16911_/A _16911_/B vssd1 vssd1 vccd1 vccd1 _16911_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17891_ _17891_/A _18017_/B _18017_/C _19957_/D vssd1 vssd1 vccd1 vccd1 _17896_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_144_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16076__A1 _16020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19630_ _19916_/B _19916_/C vssd1 vssd1 vccd1 vccd1 _19630_/Y sky130_fd_sc_hd__nand2_1
X_16842_ _12509_/A _15972_/X _16828_/A _17064_/A _16832_/Y vssd1 vssd1 vccd1 vccd1
+ _16843_/B sky130_fd_sc_hd__o221ai_1
XFILLER_120_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19014__A1 _16437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19561_ _19555_/Y _19556_/X _19559_/Y _19560_/Y vssd1 vssd1 vccd1 vccd1 _19562_/C
+ sky130_fd_sc_hd__o22ai_1
XFILLER_19_733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19014__B2 _19191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16773_ _17009_/A _17009_/B _17010_/C _17026_/D vssd1 vssd1 vccd1 vccd1 _17008_/A
+ sky130_fd_sc_hd__nand4_1
X_13985_ _15251_/A _14386_/A _14797_/A _13985_/D vssd1 vssd1 vccd1 vccd1 _13985_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18512_ _18500_/X _17627_/A _12460_/Y _18503_/Y _18505_/Y vssd1 vssd1 vccd1 vccd1
+ _18514_/B sky130_fd_sc_hd__o221ai_2
XFILLER_20_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ _12936_/A vssd1 vssd1 vccd1 vccd1 _12936_/X sky130_fd_sc_hd__buf_2
X_15724_ _15651_/Y _15670_/X _15946_/A vssd1 vssd1 vccd1 vccd1 _15724_/Y sky130_fd_sc_hd__o21ai_1
X_19492_ _19492_/A _19492_/B _19492_/C vssd1 vssd1 vccd1 vccd1 _19577_/B sky130_fd_sc_hd__nand3_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21372__A2 _21440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18443_ _18443_/A vssd1 vssd1 vccd1 vccd1 _19859_/A sky130_fd_sc_hd__clkbuf_4
X_12867_ _12867_/A _12867_/B _12867_/C vssd1 vssd1 vccd1 vccd1 _13034_/A sky130_fd_sc_hd__nand3_4
X_15655_ _15774_/A vssd1 vssd1 vccd1 vccd1 _15655_/X sky130_fd_sc_hd__buf_2
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _11805_/B _11805_/C _11805_/A vssd1 vssd1 vccd1 vccd1 _11818_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14606_ _23581_/Q _14520_/X _14545_/X _14883_/C vssd1 vssd1 vccd1 vccd1 _14606_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18374_ _20368_/B vssd1 vssd1 vccd1 vccd1 _20366_/B sky130_fd_sc_hd__clkbuf_2
X_15586_ _15586_/A _23514_/Q _15586_/C vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__and3_1
XFILLER_61_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _23455_/Q vssd1 vssd1 vccd1 vccd1 _13056_/A sky130_fd_sc_hd__inv_2
XANTENNA__17328__B2 _17154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _16549_/D _17323_/X _17324_/X _17326_/B _17326_/C vssd1 vssd1 vccd1 vccd1
+ _17327_/A sky130_fd_sc_hd__a32o_1
XFILLER_109_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14537_ _14657_/A vssd1 vssd1 vccd1 vccd1 _14545_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11749_ _11789_/B vssd1 vssd1 vccd1 vccd1 _11749_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21698__D _21704_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17256_ _17039_/B _17439_/A _19694_/A _17252_/Y _17450_/C vssd1 vssd1 vccd1 vccd1
+ _17267_/B sky130_fd_sc_hd__o2111ai_4
X_14468_ _14468_/A _14478_/C vssd1 vssd1 vccd1 vccd1 _14474_/A sky130_fd_sc_hd__nand2_1
XFILLER_175_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16551__A2 _16364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13419_ _13415_/X _22420_/B _22420_/C _13486_/B _13431_/A vssd1 vssd1 vccd1 vccd1
+ _13419_/X sky130_fd_sc_hd__o32a_1
X_16207_ _15920_/A _15920_/B _15631_/B _15634_/C vssd1 vssd1 vccd1 vccd1 _16865_/A
+ sky130_fd_sc_hd__a31o_1
X_17187_ _17187_/A _17187_/B vssd1 vssd1 vccd1 vccd1 _17189_/A sky130_fd_sc_hd__nand2_1
X_14399_ _14334_/Y _14381_/Y _14333_/X vssd1 vssd1 vccd1 vccd1 _14400_/C sky130_fd_sc_hd__o21ai_1
XFILLER_183_980 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16138_ _19199_/D _16056_/X _16172_/A _16137_/X vssd1 vssd1 vccd1 vccd1 _16168_/C
+ sky130_fd_sc_hd__a31o_2
XFILLER_155_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15993__B _17235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16303__A2 _15862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14314__A1 _14097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16069_ _17248_/C _19199_/D _16070_/C _16070_/B vssd1 vssd1 vccd1 vccd1 _16075_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19828_ _19682_/B _19672_/C _19673_/Y vssd1 vssd1 vccd1 vccd1 _19836_/B sky130_fd_sc_hd__a21oi_1
XFILLER_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19005__A1 _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19759_ _19745_/Y _19752_/Y _19757_/Y _19758_/Y vssd1 vssd1 vccd1 vccd1 _19771_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13018__B _23447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22770_ _22789_/A _22789_/B _22770_/C vssd1 vssd1 vccd1 vccd1 _22772_/B sky130_fd_sc_hd__and3_1
XFILLER_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18764__B1 _17761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21721_ _23577_/Q _21721_/B vssd1 vssd1 vccd1 vccd1 _21722_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15233__B _15233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21652_ _21616_/X _21617_/X _21665_/A _21631_/Y vssd1 vssd1 vccd1 vccd1 _21654_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_40_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18516__B1 _12463_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20603_ _13208_/B _13208_/A _20605_/A _20465_/C _20605_/B vssd1 vssd1 vccd1 vccd1
+ _20607_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_33_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21583_ _21542_/X _21631_/C _21631_/B vssd1 vssd1 vccd1 vccd1 _21625_/C sky130_fd_sc_hd__o21ai_1
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15887__C _15887_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23322_ _23325_/CLK _23322_/D vssd1 vssd1 vccd1 vccd1 _23322_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20534_ _20525_/X _20526_/X _20530_/Y _20533_/Y vssd1 vssd1 vccd1 vccd1 _20534_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_192_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19656__A _19656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18819__A1 _12004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23253_ _23253_/A vssd1 vssd1 vccd1 vccd1 _23444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20465_ _20465_/A _21018_/A _20465_/C _20465_/D vssd1 vssd1 vccd1 vccd1 _20607_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18819__B2 _19504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22204_ _22208_/A _22208_/B _22208_/C _22074_/X _22203_/Y vssd1 vssd1 vccd1 vccd1
+ _22207_/B sky130_fd_sc_hd__a32oi_4
XANTENNA__19375__B _19569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23184_ input40/X _23184_/B input6/X _23184_/D vssd1 vssd1 vccd1 vccd1 _23241_/A
+ sky130_fd_sc_hd__and4_2
X_20396_ _20411_/A vssd1 vssd1 vccd1 vccd1 _20396_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22091__A3 _21987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22135_ _22135_/A _22135_/B vssd1 vssd1 vccd1 vccd1 _22136_/D sky130_fd_sc_hd__nand2_1
XFILLER_133_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22066_ _13642_/X _22126_/A _21919_/Y _22167_/C _22130_/A vssd1 vssd1 vccd1 vccd1
+ _22211_/B sky130_fd_sc_hd__o221a_2
XFILLER_0_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17326__D _17326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19391__A _19391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21017_ _21017_/A _21017_/B _21017_/C vssd1 vssd1 vccd1 vccd1 _21019_/C sky130_fd_sc_hd__nand3_2
XFILLER_43_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_bq_clk_i clkbuf_3_7_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_bq_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_114_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13770_ _13658_/Y _13766_/Y _13257_/A _13765_/A vssd1 vssd1 vccd1 vccd1 _13770_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_16_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22968_ input40/X input39/X input6/X _22968_/D vssd1 vssd1 vccd1 vccd1 _23025_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12721_ _12677_/A _12680_/A _12851_/C vssd1 vssd1 vccd1 vccd1 _12722_/A sky130_fd_sc_hd__o21ai_4
XFILLER_128_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21919_ _22292_/A _22293_/A _21919_/C vssd1 vssd1 vccd1 vccd1 _21919_/Y sky130_fd_sc_hd__nand3_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11842__A2 _11841_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22899_ _20583_/A input7/X _22907_/S vssd1 vssd1 vccd1 vccd1 _22900_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18735__A _19279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20984__B _20984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16230__A1 _16480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15440_ _15439_/A _14749_/X _15439_/B vssd1 vssd1 vccd1 vccd1 _15441_/B sky130_fd_sc_hd__a21oi_1
X_12652_ _12652_/A vssd1 vssd1 vccd1 vccd1 _12652_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21161__A _21268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _23383_/Q vssd1 vssd1 vccd1 vccd1 _11656_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15371_ _15446_/A _15371_/B vssd1 vssd1 vccd1 vccd1 _15427_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12583_ _23286_/Q vssd1 vssd1 vccd1 vccd1 _20493_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_169_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17110_ _17118_/A vssd1 vssd1 vccd1 vccd1 _17302_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_128_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14322_ _14407_/A _15017_/D _15253_/B _14459_/D vssd1 vssd1 vccd1 vccd1 _14324_/A
+ sky130_fd_sc_hd__and4_1
X_18090_ _18090_/A _18090_/B vssd1 vssd1 vccd1 vccd1 _18104_/A sky130_fd_sc_hd__nor2_1
XFILLER_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_969 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17041_ _17449_/A _17041_/B _17041_/C _20317_/C vssd1 vssd1 vccd1 vccd1 _17041_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14253_ _14253_/A _14253_/B vssd1 vssd1 vccd1 vccd1 _14253_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _13205_/C _13205_/A _12921_/A _13203_/Y vssd1 vssd1 vccd1 vccd1 _20464_/B
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19483__A1 _17627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14184_ _14184_/A _14184_/B vssd1 vssd1 vccd1 vccd1 _14984_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17086__A _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13135_ _13196_/B _13135_/B vssd1 vssd1 vccd1 vccd1 _13135_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ _19186_/A _18992_/B _19186_/B vssd1 vssd1 vccd1 vccd1 _19044_/A sky130_fd_sc_hd__nand3_2
XFILLER_124_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _17943_/A vssd1 vssd1 vccd1 vccd1 _18154_/A sky130_fd_sc_hd__clkbuf_2
X_13066_ _13131_/A _13179_/A _12833_/B _12836_/B vssd1 vssd1 vccd1 vccd1 _13066_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21039__C _21174_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17236__D _19949_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ _12017_/A vssd1 vssd1 vccd1 vccd1 _15904_/A sky130_fd_sc_hd__buf_2
X_17874_ _17874_/A _17874_/B vssd1 vssd1 vccd1 vccd1 _17874_/Y sky130_fd_sc_hd__nor2_1
X_19613_ _19764_/A _19620_/A _19612_/X vssd1 vssd1 vccd1 vccd1 _19613_/Y sky130_fd_sc_hd__a21oi_4
X_16825_ _16147_/A _16632_/X _16824_/Y vssd1 vssd1 vccd1 vccd1 _16825_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_38_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19538__A2 _12283_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19544_ _19542_/X _19543_/Y _19538_/X vssd1 vssd1 vccd1 vccd1 _19560_/C sky130_fd_sc_hd__a21oi_2
XFILLER_111_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16756_ _16757_/A _16757_/B _16757_/C _16488_/A vssd1 vssd1 vccd1 vccd1 _16763_/A
+ sky130_fd_sc_hd__a22o_1
X_13968_ _13972_/A vssd1 vssd1 vccd1 vccd1 _14797_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15707_ _15707_/A _15707_/B _15814_/A _15815_/A vssd1 vssd1 vccd1 vccd1 _15709_/A
+ sky130_fd_sc_hd__nand4_4
X_19475_ _19345_/X _19346_/Y _19735_/A vssd1 vssd1 vccd1 vccd1 _19475_/X sky130_fd_sc_hd__o21a_2
X_12919_ _13133_/C _21268_/A vssd1 vssd1 vccd1 vccd1 _12921_/A sky130_fd_sc_hd__nand2_2
X_13899_ _23353_/Q vssd1 vssd1 vccd1 vccd1 _14188_/C sky130_fd_sc_hd__buf_2
X_16687_ _16675_/A _16904_/A _16900_/A vssd1 vssd1 vccd1 vccd1 _16693_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__20894__B _20894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18426_ _18420_/X _18425_/Y _18430_/A vssd1 vssd1 vccd1 vccd1 _18429_/A sky130_fd_sc_hd__o21bai_1
X_15638_ _15665_/B vssd1 vssd1 vccd1 vccd1 _15648_/A sky130_fd_sc_hd__buf_2
XANTENNA__13035__A1 _13122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22167__A _22380_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18357_ _18395_/A _18394_/B _18394_/A vssd1 vssd1 vccd1 vccd1 _18403_/A sky130_fd_sc_hd__nand3_1
XFILLER_159_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15569_ _23508_/Q _15569_/B _23507_/Q vssd1 vssd1 vccd1 vccd1 _15571_/A sky130_fd_sc_hd__nand3b_1
XFILLER_147_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17308_ _17140_/B _17305_/Y _17307_/Y vssd1 vssd1 vccd1 vccd1 _17318_/A sky130_fd_sc_hd__o21ai_1
X_18288_ _18288_/A _18288_/B _18288_/C vssd1 vssd1 vccd1 vccd1 _18289_/B sky130_fd_sc_hd__nand3_1
XFILLER_30_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17721__A1 _16683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17239_ _17246_/B vssd1 vssd1 vccd1 vccd1 _17239_/X sky130_fd_sc_hd__buf_2
XANTENNA__13301__B _21891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20250_ _20307_/B _20307_/C vssd1 vssd1 vccd1 vccd1 _20250_/Y sky130_fd_sc_hd__nand2_2
XFILLER_116_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20181_ _20181_/A _20180_/Y vssd1 vssd1 vccd1 vccd1 _20182_/B sky130_fd_sc_hd__or2b_1
XFILLER_116_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17237__B1 _17077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22822_ _22820_/Y _22821_/Y _22784_/A vssd1 vssd1 vccd1 vccd1 _22822_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22753_ _22713_/C _22569_/C _22569_/A _22800_/C vssd1 vssd1 vccd1 vccd1 _22756_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21704_ _21704_/A _21704_/B _21704_/C _21704_/D vssd1 vssd1 vccd1 vccd1 _21705_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_503 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22684_ _22631_/Y _22632_/Y _22683_/Y vssd1 vssd1 vccd1 vccd1 _22749_/A sky130_fd_sc_hd__o21ai_1
XFILLER_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_536 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21635_ _21635_/A _21635_/B _21635_/C _21428_/X vssd1 vssd1 vccd1 vccd1 _21635_/X
+ sky130_fd_sc_hd__or4b_1
XANTENNA__22508__C _22508_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21566_ _21566_/A _21566_/B _21566_/C vssd1 vssd1 vccd1 vccd1 _21568_/A sky130_fd_sc_hd__and3_2
XFILLER_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16515__A2 _16458_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23305_ _23336_/CLK _23305_/D vssd1 vssd1 vccd1 vccd1 _23305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20517_ _13027_/A _13027_/B _20556_/C _13038_/Y vssd1 vssd1 vccd1 vccd1 _20523_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_197_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21497_ _21497_/A vssd1 vssd1 vccd1 vccd1 _21548_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16920__C1 _23428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16803__A _16807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23236_ _23236_/A vssd1 vssd1 vccd1 vccd1 _23436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20448_ _20448_/A _20448_/B vssd1 vssd1 vccd1 vccd1 _20451_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16279__A1 _16281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23167_ _23406_/Q input23/X _23167_/S vssd1 vssd1 vccd1 vccd1 _23168_/A sky130_fd_sc_hd__mux2_1
X_20379_ _20379_/A _20379_/B vssd1 vssd1 vccd1 vccd1 _20381_/A sky130_fd_sc_hd__xnor2_1
XFILLER_134_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_67 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22118_ _22118_/A _22118_/B vssd1 vssd1 vccd1 vccd1 _22118_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23098_ _23375_/Q input24/X _23106_/S vssd1 vssd1 vccd1 vccd1 _23099_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20979__B _20984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12304__A3 _12289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22049_ _22049_/A _22049_/B vssd1 vssd1 vccd1 vccd1 _22479_/B sky130_fd_sc_hd__nand2_2
X_14940_ _14944_/A _14944_/B vssd1 vssd1 vccd1 vccd1 _14947_/B sky130_fd_sc_hd__xnor2_1
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input27_A wb_dat_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14871_ _14868_/Y _14883_/B _14621_/X _14089_/Y vssd1 vssd1 vccd1 vccd1 _14871_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_169_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16610_ _16610_/A _16647_/A _16647_/C _16610_/D vssd1 vssd1 vccd1 vccd1 _16655_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13822_ _13627_/Y _13821_/Y _13626_/Y vssd1 vssd1 vccd1 vccd1 _13822_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17590_ _17590_/A vssd1 vssd1 vccd1 vccd1 _17591_/A sky130_fd_sc_hd__buf_4
XANTENNA__12068__A2 _11969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20210__D _20210_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16541_ _16512_/Y _16540_/Y _16531_/A _16558_/A vssd1 vssd1 vccd1 vccd1 _16565_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_28_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13753_ _13727_/Y _13729_/Y _13730_/Y _13752_/Y vssd1 vssd1 vccd1 vccd1 _13754_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12928__D _21182_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18465__A _18465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12704_ _12704_/A vssd1 vssd1 vccd1 vccd1 _12704_/X sky130_fd_sc_hd__buf_2
X_19260_ _20320_/A vssd1 vssd1 vccd1 vccd1 _19903_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16472_ _16472_/A _16472_/B _16472_/C vssd1 vssd1 vccd1 vccd1 _16477_/B sky130_fd_sc_hd__nand3_1
X_13684_ _23480_/Q vssd1 vssd1 vccd1 vccd1 _22220_/C sky130_fd_sc_hd__buf_2
XANTENNA__23521__D _23521_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18211_ _18211_/A _18211_/B _18211_/C _18211_/D vssd1 vssd1 vccd1 vccd1 _18286_/A
+ sky130_fd_sc_hd__or4_2
X_15423_ _15422_/A _15427_/A _15420_/Y _15421_/X vssd1 vssd1 vccd1 vccd1 _15424_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_12635_ _23291_/Q _23290_/Q vssd1 vssd1 vccd1 vccd1 _12742_/A sky130_fd_sc_hd__nor2_1
XFILLER_188_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19191_ _19191_/A vssd1 vssd1 vccd1 vccd1 _19649_/A sky130_fd_sc_hd__buf_2
XFILLER_19_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18142_ _18141_/C _18141_/A _23531_/Q vssd1 vssd1 vccd1 vccd1 _18143_/B sky130_fd_sc_hd__a21oi_1
X_15354_ _15352_/Y _15350_/A _15353_/X vssd1 vssd1 vccd1 vccd1 _15354_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12566_ _12564_/Y _12565_/X _23539_/Q vssd1 vssd1 vccd1 vccd1 _12566_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_180_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14305_ _14306_/B _14306_/C _14306_/A vssd1 vssd1 vccd1 vccd1 _14842_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13121__B _13121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18073_ _18253_/B _18072_/Y _18140_/B vssd1 vssd1 vccd1 vccd1 _18137_/A sky130_fd_sc_hd__o21ai_1
X_15285_ _15283_/X _15395_/A vssd1 vssd1 vccd1 vccd1 _15288_/A sky130_fd_sc_hd__and2b_1
XFILLER_144_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _12497_/A vssd1 vssd1 vccd1 vccd1 _17964_/C sky130_fd_sc_hd__buf_2
XFILLER_89_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output95_A _23269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17024_ _17024_/A vssd1 vssd1 vccd1 vccd1 _17024_/Y sky130_fd_sc_hd__inv_2
X_14236_ _14236_/A _14236_/B vssd1 vssd1 vccd1 vccd1 _14306_/C sky130_fd_sc_hd__nand2_1
XFILLER_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15974__D _15974_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14167_ _14167_/A _15019_/A _14360_/A _14167_/D vssd1 vssd1 vccd1 vccd1 _14167_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_152_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13126_/B _13126_/C _13117_/X vssd1 vssd1 vccd1 vccd1 _13172_/B sky130_fd_sc_hd__a21bo_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _14184_/A _14184_/B _14097_/X vssd1 vssd1 vccd1 vccd1 _14098_/X sky130_fd_sc_hd__a21o_1
X_18975_ _18975_/A vssd1 vssd1 vccd1 vccd1 _18975_/X sky130_fd_sc_hd__clkbuf_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21992__C _22226_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16690__A1 _16360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17926_ _17922_/X _17924_/X _17925_/Y vssd1 vssd1 vccd1 vccd1 _18129_/B sky130_fd_sc_hd__o21a_1
X_13049_ _13049_/A vssd1 vssd1 vccd1 vccd1 _13078_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17857_ _17852_/Y _17857_/B _17857_/C vssd1 vssd1 vccd1 vccd1 _17999_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__17234__A3 _17766_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11592__A _11634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16442__A1 _15884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16808_ _16808_/A _16808_/B vssd1 vssd1 vccd1 vccd1 _17435_/A sky130_fd_sc_hd__nor2_4
XANTENNA__16442__B2 _16311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17788_ _17788_/A _17788_/B vssd1 vssd1 vccd1 vccd1 _17792_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23272__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19527_ _19476_/Y _19477_/Y _19519_/Y _19526_/Y vssd1 vssd1 vccd1 vccd1 _19527_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__12464__C1 _16140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16739_ _16739_/A _16739_/B _16739_/C vssd1 vssd1 vccd1 vccd1 _16740_/A sky130_fd_sc_hd__nand3_1
XFILLER_62_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19458_ _19457_/X _19291_/Y _19456_/A vssd1 vssd1 vccd1 vccd1 _19459_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18409_ _18409_/A vssd1 vssd1 vccd1 vccd1 _23596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ _19389_/A _19389_/B _19389_/C vssd1 vssd1 vccd1 vccd1 _19600_/A sky130_fd_sc_hd__nand3_2
XFILLER_148_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_327 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12767__B1 _13122_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21420_ _21350_/X _21254_/Y _23566_/Q _21349_/B vssd1 vssd1 vccd1 vccd1 _21420_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_147_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19695__A1 _12243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19695__B2 _17565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21351_ _21254_/Y _21350_/X _21257_/Y _21259_/X vssd1 vssd1 vccd1 vccd1 _21352_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_148_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12519__B1 _12518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20302_ _20120_/X _20205_/X _20307_/A _20250_/Y _20301_/Y vssd1 vssd1 vccd1 vccd1
+ _20303_/C sky130_fd_sc_hd__o221ai_2
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15181__A1 _15310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21282_ _21282_/A vssd1 vssd1 vccd1 vccd1 _21432_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_162_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23021_ _23341_/Q input22/X _23023_/S vssd1 vssd1 vccd1 vccd1 _23022_/A sky130_fd_sc_hd__mux2_1
X_20233_ _20167_/A _20167_/B _20232_/Y vssd1 vssd1 vccd1 vccd1 _20233_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_1002 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20164_ _20269_/B _20164_/B _20164_/C vssd1 vssd1 vccd1 vccd1 _20229_/C sky130_fd_sc_hd__and3_1
XFILLER_131_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17454__A _19543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20095_ _20095_/A _20172_/B _20095_/C vssd1 vssd1 vccd1 vccd1 _20096_/C sky130_fd_sc_hd__nand3_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_12_0_bq_clk_i_A clkbuf_3_6_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12598__A _13052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22805_ _22802_/Y _22803_/X _22840_/B vssd1 vssd1 vccd1 vccd1 _22805_/X sky130_fd_sc_hd__a21o_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20997_ _20997_/A vssd1 vssd1 vccd1 vccd1 _21132_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22736_ _21854_/A _21854_/B _22630_/X _22687_/Y _22738_/A vssd1 vssd1 vccd1 vccd1
+ _22736_/X sky130_fd_sc_hd__o221a_1
XANTENNA__16197__B1 _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12470__A2 _18506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_64 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21190__B1 _20957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22667_ _22670_/A _22725_/A _22670_/C _22667_/D vssd1 vssd1 vccd1 vccd1 _22667_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__15944__B1 _15859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12420_ _12455_/C vssd1 vssd1 vccd1 vccd1 _18511_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13222__A _23333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21618_ _21616_/X _21617_/X _21614_/Y _21630_/A _21666_/B vssd1 vssd1 vccd1 vccd1
+ _21618_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_187_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22598_ _22598_/A _22676_/A vssd1 vssd1 vccd1 vccd1 _22599_/A sky130_fd_sc_hd__nand2_1
X_12351_ _16528_/B vssd1 vssd1 vccd1 vccd1 _14735_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_181_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21549_ _21545_/X _21547_/X _21548_/X _21504_/A vssd1 vssd1 vccd1 vccd1 _21551_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15070_ _15220_/A _15220_/B _15289_/C vssd1 vssd1 vccd1 vccd1 _15072_/A sky130_fd_sc_hd__and3_1
XFILLER_107_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _12282_/A _12282_/B _18798_/B vssd1 vssd1 vccd1 vccd1 _12282_/X sky130_fd_sc_hd__and3_2
XANTENNA__20055__A _20055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ _14027_/A vssd1 vssd1 vccd1 vccd1 _14191_/C sky130_fd_sc_hd__clkbuf_2
X_23219_ _23241_/A vssd1 vssd1 vccd1 vccd1 _23228_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_49_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14053__A _23496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22993__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16672__A1 _17133_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18760_ _18601_/A _18932_/B _18759_/Y _17967_/A _12260_/D vssd1 vssd1 vccd1 vccd1
+ _18760_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_122_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16672__B2 _19161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15972_ _16030_/A vssd1 vssd1 vccd1 vccd1 _15972_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__23516__D input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17711_ _17467_/X _17710_/X _17598_/Y vssd1 vssd1 vccd1 vccd1 _17711_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_121_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14923_ _14923_/A _14926_/B _14923_/C vssd1 vssd1 vccd1 vccd1 _14923_/X sky130_fd_sc_hd__and3_1
X_18691_ _18673_/X _17643_/A _18674_/X _18675_/X vssd1 vssd1 vccd1 vccd1 _18784_/C
+ sky130_fd_sc_hd__o31ai_2
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17642_ _17642_/A vssd1 vssd1 vccd1 vccd1 _17643_/A sky130_fd_sc_hd__buf_2
X_14854_ _14836_/Y _14828_/Y _14840_/C vssd1 vssd1 vccd1 vccd1 _14957_/B sky130_fd_sc_hd__o21a_1
XFILLER_63_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13805_ _13793_/A _13793_/B _13804_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17573_ _16356_/A _17565_/X _17583_/A vssd1 vssd1 vccd1 vccd1 _17578_/A sky130_fd_sc_hd__o21ai_1
XFILLER_63_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13116__B _21177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14785_ _14220_/A _14221_/B _14784_/Y vssd1 vssd1 vccd1 vccd1 _14789_/C sky130_fd_sc_hd__a21o_1
X_11997_ _11713_/A _11713_/B _11847_/A vssd1 vssd1 vccd1 vccd1 _11997_/X sky130_fd_sc_hd__a21o_1
XANTENNA__23170__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19312_ _19184_/A _19165_/Y _19305_/Y vssd1 vssd1 vccd1 vccd1 _19312_/Y sky130_fd_sc_hd__o21ai_1
X_16524_ _16523_/X _16496_/X _16502_/X _16503_/Y vssd1 vssd1 vccd1 vccd1 _16530_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13736_ _13736_/A _13736_/B _22192_/C _22192_/D vssd1 vssd1 vccd1 vccd1 _13736_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__12461__A2 _11936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16727__A2 _16724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19243_ _19239_/X _19240_/Y _19226_/A _19242_/Y vssd1 vssd1 vccd1 vccd1 _19244_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_182_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16455_ _16380_/Y _16405_/B _16450_/Y _16454_/Y vssd1 vssd1 vccd1 vccd1 _16539_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__15935__B1 _17885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ _13467_/X _13320_/X _13341_/X vssd1 vssd1 vccd1 vccd1 _13668_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__19126__B1 _18607_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _15382_/A _15382_/B _15382_/C vssd1 vssd1 vccd1 vccd1 _15406_/X sky130_fd_sc_hd__a21o_1
X_19174_ _16437_/A _18455_/A _18461_/C _19499_/A _12323_/A vssd1 vssd1 vccd1 vccd1
+ _19182_/B sky130_fd_sc_hd__o32a_1
X_12618_ _12618_/A vssd1 vssd1 vccd1 vccd1 _12788_/B sky130_fd_sc_hd__clkbuf_4
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _16377_/X _16384_/X _16457_/D _17243_/D _16316_/Y vssd1 vssd1 vccd1 vccd1
+ _16386_/X sky130_fd_sc_hd__o2111a_1
XANTENNA__12213__A2 _12151_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13598_ _13598_/A _13598_/B vssd1 vssd1 vccd1 vccd1 _13676_/A sky130_fd_sc_hd__nand2_1
XFILLER_129_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21987__C _21987_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18125_ _18123_/A _18123_/B _18123_/C vssd1 vssd1 vccd1 vccd1 _18126_/A sky130_fd_sc_hd__a21o_1
XFILLER_185_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12549_ _12303_/Y _12547_/X _12548_/Y vssd1 vssd1 vccd1 vccd1 _12549_/Y sky130_fd_sc_hd__a21oi_1
X_15337_ _15337_/A _15337_/B vssd1 vssd1 vccd1 vccd1 _15442_/D sky130_fd_sc_hd__xor2_4
XFILLER_184_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16443__A _17134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15985__C _15985_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18056_ _18051_/Y _18055_/Y _23530_/Q vssd1 vssd1 vccd1 vccd1 _18144_/C sky130_fd_sc_hd__o21bai_1
XANTENNA__19429__A1 _19116_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15268_ _15259_/Y _15260_/X _15261_/X _15264_/Y _15267_/Y vssd1 vssd1 vccd1 vccd1
+ _15270_/A sky130_fd_sc_hd__a32oi_2
XFILLER_160_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17007_ _16768_/A _16768_/B _17010_/A _17009_/A _17022_/A vssd1 vssd1 vccd1 vccd1
+ _17008_/B sky130_fd_sc_hd__a41oi_1
XFILLER_6_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14910__A1 _14777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14219_ _14220_/A _14220_/B _14219_/C _14219_/D vssd1 vssd1 vccd1 vccd1 _14224_/A
+ sky130_fd_sc_hd__nand4_1
X_15199_ _14029_/X _14015_/B _15298_/B _14777_/A _15225_/A vssd1 vssd1 vccd1 vccd1
+ _15199_/Y sky130_fd_sc_hd__o2111ai_1
XANTENNA__22984__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14269__A3 _14876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18958_ _19900_/D _18958_/B _18958_/C _19674_/B vssd1 vssd1 vccd1 vccd1 _18958_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17909_ _17909_/A _17909_/B _17909_/C vssd1 vssd1 vccd1 vccd1 _17916_/A sky130_fd_sc_hd__nand3_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18889_ _18889_/A _18889_/B vssd1 vssd1 vccd1 vccd1 _18889_/Y sky130_fd_sc_hd__nor2_2
XFILLER_67_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20211__A2 _20320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13307__A _23322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20920_ _20920_/A vssd1 vssd1 vccd1 vccd1 _20934_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13229__A1 _13226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15225__C _15225_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20851_ _20862_/A _20862_/B _20869_/B vssd1 vssd1 vccd1 vccd1 _20851_/Y sky130_fd_sc_hd__o21ai_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18168__A1 _20151_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_650 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__23161__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23570_ _23575_/CLK _23570_/D vssd1 vssd1 vccd1 vccd1 _23570_/Q sky130_fd_sc_hd__dfxtp_1
X_20782_ _20782_/A _20782_/B _20782_/C vssd1 vssd1 vccd1 vccd1 _20783_/B sky130_fd_sc_hd__nand3_1
X_22521_ _22521_/A _22861_/C _22521_/C vssd1 vssd1 vccd1 vccd1 _22521_/X sky130_fd_sc_hd__and3_1
XFILLER_179_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22452_ _22452_/A _22452_/B vssd1 vssd1 vccd1 vccd1 _22452_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19648__B _19651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21403_ _21236_/A _21236_/B _21236_/C _21335_/A _21402_/Y vssd1 vssd1 vccd1 vccd1
+ _21404_/B sky130_fd_sc_hd__a311oi_4
XFILLER_157_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22383_ _13470_/X _22461_/A _22393_/A vssd1 vssd1 vccd1 vccd1 _22383_/X sky130_fd_sc_hd__o21a_1
XFILLER_198_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21334_ _21333_/A _21333_/B _21333_/C _21333_/D vssd1 vssd1 vccd1 vccd1 _21335_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_108_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13165__B1 _21440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21265_ _21514_/A _12981_/C _21162_/Y vssd1 vssd1 vccd1 vccd1 _21265_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23004_ _21852_/A input13/X _23012_/S vssd1 vssd1 vccd1 vccd1 _23005_/A sky130_fd_sc_hd__mux2_1
XANTENNA__22975__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20216_ _18211_/A _20139_/Y _20081_/D _20271_/D _20215_/X vssd1 vssd1 vccd1 vccd1
+ _20216_/X sky130_fd_sc_hd__o311a_1
XANTENNA__23186__A _23254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21196_ _21196_/A vssd1 vssd1 vccd1 vccd1 _21387_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22521__C _22521_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20147_ _20146_/A _20146_/B _20146_/C _20146_/D vssd1 vssd1 vccd1 vccd1 _20148_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13468__A1 _13465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20078_ _20078_/A vssd1 vssd1 vccd1 vccd1 _20172_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11920_ _23591_/Q vssd1 vssd1 vccd1 vccd1 _23256_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _11851_/A vssd1 vssd1 vccd1 vccd1 _12378_/A sky130_fd_sc_hd__buf_2
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23152__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _13911_/C _14657_/A _14698_/A _14569_/X vssd1 vssd1 vccd1 vccd1 _14570_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11782_ _18812_/A vssd1 vssd1 vccd1 vccd1 _11999_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22964__S _22966_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16247__B _16254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13521_ _13732_/B vssd1 vssd1 vccd1 vccd1 _21815_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_186_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22719_ _22717_/A _22717_/B _22717_/C _22789_/B vssd1 vssd1 vccd1 vccd1 _22722_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11651__B1 _23587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15917__B1 _11741_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13452_ _13516_/A _13516_/B vssd1 vssd1 vccd1 vccd1 _13513_/A sky130_fd_sc_hd__xnor2_1
X_16240_ _16251_/B vssd1 vssd1 vccd1 vccd1 _16240_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12403_ _12403_/A _23387_/Q _23386_/Q _23388_/Q vssd1 vssd1 vccd1 vccd1 _19155_/C
+ sky130_fd_sc_hd__nor4_4
XFILLER_12_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16171_ _17062_/B vssd1 vssd1 vccd1 vccd1 _17445_/A sky130_fd_sc_hd__buf_2
X_13383_ _21909_/C vssd1 vssd1 vccd1 vccd1 _13804_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_194_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12334_ _12339_/C _12334_/B vssd1 vssd1 vccd1 vccd1 _12336_/C sky130_fd_sc_hd__nand2_1
X_15122_ _15163_/A _15188_/A _15164_/A _15164_/B vssd1 vssd1 vccd1 vccd1 _15127_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19930_ _19442_/Y _19443_/Y _19926_/X _19275_/Y _19929_/Y vssd1 vssd1 vccd1 vccd1
+ _20184_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_126_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15053_ _15053_/A _15053_/B vssd1 vssd1 vccd1 vccd1 _15064_/A sky130_fd_sc_hd__nand2_1
XFILLER_142_728 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12265_ _18952_/D _12265_/B _12265_/C _17134_/B vssd1 vssd1 vccd1 vccd1 _12273_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_99_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20426__C1 _20368_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22966__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14004_ _13997_/Y _13991_/Y _14003_/Y vssd1 vssd1 vccd1 vccd1 _14005_/B sky130_fd_sc_hd__o21ai_1
XFILLER_123_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19861_ _19850_/Y _19851_/X _19860_/X vssd1 vssd1 vccd1 vccd1 _19864_/A sky130_fd_sc_hd__o21ai_1
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12196_ _12211_/A _12206_/A _12196_/C vssd1 vssd1 vccd1 vccd1 _12199_/D sky130_fd_sc_hd__nand3_2
Xoutput60 _14660_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput71 _14702_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput82 _14584_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[6] sky130_fd_sc_hd__buf_2
X_18812_ _18812_/A _18812_/B _18812_/C vssd1 vssd1 vccd1 vccd1 _18813_/A sky130_fd_sc_hd__nor3_2
Xoutput93 _23267_/Q vssd1 vssd1 vccd1 vccd1 y[5] sky130_fd_sc_hd__buf_2
XANTENNA__15607__A _23429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19792_ _19792_/A vssd1 vssd1 vccd1 vccd1 _23527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14511__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18743_ _19288_/A _18747_/B _18747_/A vssd1 vssd1 vccd1 vccd1 _18745_/A sky130_fd_sc_hd__nand3_1
XFILLER_110_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15955_ _23589_/Q _16815_/B _16800_/A _23592_/Q vssd1 vssd1 vccd1 vccd1 _15956_/C
+ sky130_fd_sc_hd__nor4_1
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14906_ _14968_/A _14968_/B _14908_/C _14968_/C vssd1 vssd1 vccd1 vccd1 _14909_/A
+ sky130_fd_sc_hd__a22o_1
X_18674_ _15882_/X _19040_/A _12214_/X _16604_/X vssd1 vssd1 vccd1 vccd1 _18674_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_110_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15886_ _15886_/A _15886_/B _15886_/C vssd1 vssd1 vccd1 vccd1 _15890_/B sky130_fd_sc_hd__nand3_2
XFILLER_48_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17625_ _19664_/B _17625_/B _17625_/C vssd1 vssd1 vccd1 vccd1 _17625_/Y sky130_fd_sc_hd__nand3_1
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14837_ _14828_/Y _14831_/Y _14836_/Y vssd1 vssd1 vccd1 vccd1 _14844_/A sky130_fd_sc_hd__o21ai_1
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23143__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11870__A _16044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17556_ _17485_/A _17487_/B _17553_/Y _17806_/A vssd1 vssd1 vccd1 vccd1 _17556_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14768_ _23361_/Q vssd1 vssd1 vccd1 vccd1 _15112_/D sky130_fd_sc_hd__inv_2
XFILLER_16_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16507_ _16507_/A _16507_/B vssd1 vssd1 vccd1 vccd1 _16558_/A sky130_fd_sc_hd__xor2_4
XFILLER_147_1072 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13719_ _13705_/D _13709_/A _13566_/Y _13482_/Y vssd1 vssd1 vccd1 vccd1 _13720_/D
+ sky130_fd_sc_hd__a22o_1
X_17487_ _17487_/A _17487_/B vssd1 vssd1 vccd1 vccd1 _17487_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14699_ _23040_/D vssd1 vssd1 vccd1 vccd1 _14699_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19226_ _19226_/A vssd1 vssd1 vccd1 vccd1 _19256_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16438_ _16437_/X _16398_/X _16399_/X vssd1 vssd1 vccd1 vccd1 _16438_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19157_ _19157_/A _20369_/C _19157_/C vssd1 vssd1 vccd1 vccd1 _19304_/A sky130_fd_sc_hd__nand3_2
X_16369_ _16369_/A _16369_/B _16369_/C vssd1 vssd1 vccd1 vccd1 _16404_/A sky130_fd_sc_hd__nand3_2
XFILLER_118_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20407__B _20407_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18108_ _18108_/A _18108_/B vssd1 vssd1 vccd1 vccd1 _18110_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19088_ _18907_/A _19088_/B _19088_/C vssd1 vssd1 vccd1 vccd1 _19109_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__23460__CLK _23462_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18039_ _18038_/A _18123_/A _18038_/C vssd1 vssd1 vccd1 vccd1 _18043_/B sky130_fd_sc_hd__a21o_1
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12206__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18086__B1 _18002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21050_ _21277_/A _21181_/A _21050_/C _21050_/D vssd1 vssd1 vccd1 vccd1 _21179_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_98_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_815 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20001_ _19941_/X _19942_/Y _20000_/Y vssd1 vssd1 vccd1 vccd1 _20011_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__16636__A1 _15861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21952_ _21947_/A _21982_/B _21982_/A vssd1 vssd1 vccd1 vccd1 _21953_/C sky130_fd_sc_hd__a21o_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20903_ _20903_/A _20903_/B vssd1 vssd1 vccd1 vccd1 _21072_/A sky130_fd_sc_hd__nand2_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21883_ _21883_/A _21883_/B _21883_/C vssd1 vssd1 vccd1 vccd1 _21884_/B sky130_fd_sc_hd__nand3_4
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23134__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20834_ _20836_/A _20837_/A _20843_/B vssd1 vssd1 vccd1 vccd1 _20839_/A sky130_fd_sc_hd__a21o_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1112 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23553_ _23558_/CLK _23553_/D vssd1 vssd1 vccd1 vccd1 _23553_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19659__A _20046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20765_ _20765_/A _20765_/B vssd1 vssd1 vccd1 vccd1 _20766_/B sky130_fd_sc_hd__or2_1
XFILLER_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22504_ _22504_/A _22504_/B vssd1 vssd1 vccd1 vccd1 _22509_/B sky130_fd_sc_hd__nand2_1
XFILLER_168_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23484_ _23499_/CLK _23496_/Q vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
X_20696_ _20711_/A vssd1 vssd1 vccd1 vccd1 _20715_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__18282__B _18335_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22435_ _22435_/A _22435_/B vssd1 vssd1 vccd1 vccd1 _22436_/B sky130_fd_sc_hd__nand2_1
XFILLER_195_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17116__A2 _17243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20317__B _20317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19510__B1 _19307_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13500__A _23475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22366_ _22362_/Y _22496_/A _22365_/X vssd1 vssd1 vccd1 vccd1 _22366_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__18864__A2 _18840_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21317_ _21317_/A _21317_/B _21317_/C _21317_/D vssd1 vssd1 vccd1 vccd1 _21317_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_108_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12116__A _19364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22297_ _22297_/A _22297_/B vssd1 vssd1 vccd1 vccd1 _22297_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12050_ _11903_/A _11975_/Y _11912_/D vssd1 vssd1 vccd1 vccd1 _12057_/B sky130_fd_sc_hd__o21ai_1
X_21248_ _21246_/X _21247_/X _21240_/Y vssd1 vssd1 vccd1 vccd1 _21248_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_116_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18616__A2 _17980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20959__B1 _12815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14331__A _14331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21179_ _21179_/A _21179_/B _21179_/C _21179_/D vssd1 vssd1 vccd1 vccd1 _21186_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18092__A3 _17567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19841__B _19868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17642__A _17642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ _15864_/A _17626_/A _15852_/A vssd1 vssd1 vccd1 vccd1 _16070_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__15850__A2 _16370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19041__A2 _20081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12952_ _12952_/A vssd1 vssd1 vccd1 vccd1 _12952_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_22 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17052__A1 _16447_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17052__B2 _16523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _11903_/A _11912_/C _11912_/D vssd1 vssd1 vccd1 vccd1 _11905_/B sky130_fd_sc_hd__nand3_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _23418_/Q vssd1 vssd1 vccd1 vccd1 _15672_/C sky130_fd_sc_hd__inv_2
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12756_/A _12882_/Y _13151_/B vssd1 vssd1 vccd1 vccd1 _12884_/B sky130_fd_sc_hd__a21oi_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _16684_/X _16683_/X _18503_/B _18503_/A _17233_/A vssd1 vssd1 vccd1 vccd1
+ _17410_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _23112_/D vssd1 vssd1 vccd1 vccd1 _14640_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18390_ _18392_/A _18392_/B _18356_/A _18356_/B _18355_/A vssd1 vssd1 vccd1 vccd1
+ _18400_/A sky130_fd_sc_hd__a221o_1
X_11834_ _11834_/A _11834_/B vssd1 vssd1 vccd1 vccd1 _18597_/B sky130_fd_sc_hd__nand2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17341_/A _17341_/B _17341_/C vssd1 vssd1 vccd1 vccd1 _17350_/D sky130_fd_sc_hd__nand3_2
XFILLER_42_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19569__A _19569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14553_ _23415_/Q vssd1 vssd1 vccd1 vccd1 _14553_/X sky130_fd_sc_hd__buf_2
X_11765_ _11868_/A vssd1 vssd1 vccd1 vccd1 _11766_/B sky130_fd_sc_hd__buf_4
XFILLER_159_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13504_ _21764_/C vssd1 vssd1 vccd1 vccd1 _22553_/C sky130_fd_sc_hd__clkbuf_2
X_17272_ _17039_/B _17439_/A _17269_/X vssd1 vssd1 vccd1 vccd1 _17272_/Y sky130_fd_sc_hd__o21ai_1
X_14484_ _14486_/A _14486_/B _14486_/C vssd1 vssd1 vccd1 vccd1 _14487_/A sky130_fd_sc_hd__a21o_1
X_11696_ _11860_/C _11720_/A _11724_/A _11694_/X _11695_/X vssd1 vssd1 vccd1 vccd1
+ _12239_/A sky130_fd_sc_hd__o41a_1
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19011_ _19011_/A _19700_/A _19700_/B vssd1 vssd1 vccd1 vccd1 _19012_/B sky130_fd_sc_hd__and3_2
XFILLER_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16223_ _16180_/Y _16181_/X _16219_/Y _16222_/Y vssd1 vssd1 vccd1 vccd1 _16242_/A
+ sky130_fd_sc_hd__o211ai_4
X_13435_ _13419_/X _13443_/A _13432_/Y _13434_/Y vssd1 vssd1 vccd1 vccd1 _13460_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_186_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14506__A _16821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19501__B1 _19321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16154_ _12086_/A _15884_/X _15971_/X _16598_/B _16590_/A vssd1 vssd1 vccd1 vccd1
+ _16154_/Y sky130_fd_sc_hd__o221ai_4
X_13366_ _13783_/C _13366_/B vssd1 vssd1 vccd1 vccd1 _13366_/Y sky130_fd_sc_hd__nor2_2
XFILLER_177_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15105_ _14992_/Y _15419_/B _14469_/C _15000_/Y vssd1 vssd1 vccd1 vccd1 _15107_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12317_ _11747_/X _11749_/X _16549_/B _12273_/B _12260_/Y vssd1 vssd1 vccd1 vccd1
+ _12318_/A sky130_fd_sc_hd__a32o_1
XFILLER_177_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16085_ _19363_/C vssd1 vssd1 vccd1 vccd1 _17414_/A sky130_fd_sc_hd__buf_4
XFILLER_115_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13297_ _22363_/A vssd1 vssd1 vccd1 vccd1 _22569_/B sky130_fd_sc_hd__clkbuf_2
X_19913_ _19768_/Y _19640_/Y _19928_/B _19911_/Y vssd1 vssd1 vccd1 vccd1 _19925_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ _15036_/A _15036_/B _15036_/C vssd1 vssd1 vccd1 vccd1 _15050_/B sky130_fd_sc_hd__nand3_2
X_12248_ _16198_/C vssd1 vssd1 vccd1 vccd1 _16372_/A sky130_fd_sc_hd__buf_4
XFILLER_174_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12352__A1 _11931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__B2 _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19844_ _20209_/A _18000_/A _19841_/Y _19843_/Y vssd1 vssd1 vccd1 vccd1 _19855_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14879__C _14879_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ _12167_/X _12168_/X _11948_/A _11951_/A _12178_/Y vssd1 vssd1 vccd1 vccd1
+ _12181_/B sky130_fd_sc_hd__o221ai_4
XFILLER_3_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14241__A _15356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19775_ _19770_/X _19771_/X _19772_/Y _19626_/X _19774_/Y vssd1 vssd1 vccd1 vccd1
+ _19775_/Y sky130_fd_sc_hd__o221ai_4
X_16987_ _16987_/A _17374_/C vssd1 vssd1 vccd1 vccd1 _16997_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18726_ _18914_/A _18914_/B _18914_/C vssd1 vssd1 vccd1 vccd1 _18726_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_110_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15938_ _16921_/C _17625_/B _17625_/C _16281_/A _15925_/Y vssd1 vssd1 vccd1 vccd1
+ _16251_/D sky130_fd_sc_hd__a32o_1
XFILLER_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12655__A2 _12648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18657_ _18972_/B _18972_/C _18657_/C vssd1 vssd1 vccd1 vccd1 _18657_/Y sky130_fd_sc_hd__nand3_4
XFILLER_37_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15869_ _19703_/B vssd1 vssd1 vccd1 vccd1 _20142_/A sky130_fd_sc_hd__buf_4
XFILLER_92_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17608_ _17613_/A _16478_/X _17605_/Y _17606_/X _17607_/X vssd1 vssd1 vccd1 vccd1
+ _17770_/B sky130_fd_sc_hd__o311ai_4
XFILLER_18_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18588_ _18588_/A _18733_/B _18733_/C vssd1 vssd1 vccd1 vccd1 _18589_/B sky130_fd_sc_hd__nand3_1
XFILLER_17_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _17504_/Y _17677_/C _17510_/Y vssd1 vssd1 vccd1 vccd1 _17539_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18543__A1 _18721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15800__A _15928_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20550_ _20728_/A _20714_/A _20547_/X _20549_/Y vssd1 vssd1 vccd1 vccd1 _20551_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_137_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19209_ _12053_/X _17408_/X _19201_/C _19201_/A vssd1 vssd1 vccd1 vccd1 _19221_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_193_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20481_ _20498_/A _20481_/B vssd1 vssd1 vccd1 vccd1 _20482_/B sky130_fd_sc_hd__nand2_1
XFILLER_158_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_bq_clk_i clkbuf_4_9_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 _23588_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22220_ _22220_/A _22263_/B _22220_/C _22220_/D vssd1 vssd1 vccd1 vccd1 _22221_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_164_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_555 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16857__A1 _15691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22151_ _22267_/A _22268_/A _22145_/C _22150_/Y _22381_/B vssd1 vssd1 vccd1 vccd1
+ _22151_/Y sky130_fd_sc_hd__a32oi_4
XANTENNA__17727__A _19949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21102_ _21101_/B _21101_/C _21101_/A vssd1 vssd1 vccd1 vccd1 _21102_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22082_ _22069_/Y _22074_/A _22203_/A _22203_/B vssd1 vssd1 vccd1 vccd1 _22083_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_21033_ _21243_/A _21243_/B _21019_/C vssd1 vssd1 vccd1 vccd1 _21345_/A sky130_fd_sc_hd__a21oi_2
XFILLER_120_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16609__B2 _17454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20956__A3 _20953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22984_ _13379_/X input35/X _22990_/S vssd1 vssd1 vccd1 vccd1 _22985_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21935_ _21933_/X _21934_/Y _21939_/A _21940_/B vssd1 vssd1 vccd1 vccd1 _21936_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_76_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18782__A1 _18627_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21866_ _23270_/Q _21971_/B _21861_/Y _21864_/Y vssd1 vssd1 vccd1 vccd1 _21867_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _20817_/A _20817_/B vssd1 vssd1 vccd1 vccd1 _20820_/A sky130_fd_sc_hd__nand2_1
X_21797_ _13466_/A _13765_/X _22365_/C _21792_/Y _13561_/A vssd1 vssd1 vccd1 vccd1
+ _21798_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23536_ _23558_/CLK _23536_/D vssd1 vssd1 vccd1 vccd1 _23536_/Q sky130_fd_sc_hd__dfxtp_2
X_20748_ _20748_/A _20748_/B _20748_/C vssd1 vssd1 vccd1 vccd1 _20752_/B sky130_fd_sc_hd__nand3_1
XFILLER_10_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21431__B _21431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19539__D _19700_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23467_ _23571_/CLK _23479_/Q vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfxtp_1
XFILLER_195_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20679_ _20529_/B _20674_/Y _20673_/A _20673_/B _20676_/Y vssd1 vssd1 vccd1 vccd1
+ _20679_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13220_ _23318_/Q _22018_/A _13259_/A vssd1 vssd1 vccd1 vccd1 _13221_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__13230__A _13659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22418_ _22303_/Y _22300_/Y _22301_/Y _22405_/C vssd1 vssd1 vccd1 vccd1 _22418_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_195_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23398_ _23398_/CLK _23398_/D vssd1 vssd1 vccd1 vccd1 _23398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16848__A1 _17057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13151_ _13151_/A _13151_/B _13151_/C vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__or3_2
XANTENNA__16848__B2 _16027_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22349_ _22445_/C _22445_/D vssd1 vssd1 vccd1 vccd1 _22349_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ _18445_/A _19193_/C vssd1 vssd1 vccd1 vccd1 _12424_/A sky130_fd_sc_hd__nand2_1
XANTENNA__23043__A0 _14298_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21159__A _21159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13082_ _13085_/A _13085_/B _13091_/A vssd1 vssd1 vccd1 vccd1 _20594_/A sky130_fd_sc_hd__o21ai_1
XFILLER_151_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19798__B1 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16910_ _16911_/B _16908_/X _16909_/Y vssd1 vssd1 vccd1 vccd1 _16934_/A sky130_fd_sc_hd__o21ai_2
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12033_ _12159_/A _12159_/B _12159_/C vssd1 vssd1 vccd1 vccd1 _12033_/Y sky130_fd_sc_hd__nand3_2
XFILLER_151_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17890_ _17643_/X _17635_/A _17889_/Y vssd1 vssd1 vccd1 vccd1 _18017_/C sky130_fd_sc_hd__o21ai_1
XFILLER_137_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16841_ _16841_/A _16841_/B vssd1 vssd1 vccd1 vccd1 _16843_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19560_ _19560_/A _19560_/B _19560_/C vssd1 vssd1 vccd1 vccd1 _19560_/Y sky130_fd_sc_hd__nor3_4
XFILLER_77_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19014__A2 _12103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16772_ _16774_/B vssd1 vssd1 vccd1 vccd1 _17026_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13984_ _13984_/A vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__buf_2
XFILLER_92_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_840 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18511_ _18511_/A _18511_/B vssd1 vssd1 vccd1 vccd1 _18514_/A sky130_fd_sc_hd__nand2_1
XFILLER_92_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15723_ _15723_/A _15723_/B _15723_/C vssd1 vssd1 vccd1 vccd1 _15946_/A sky130_fd_sc_hd__nand3_2
X_19491_ _19491_/A _19491_/B vssd1 vssd1 vccd1 vccd1 _19492_/C sky130_fd_sc_hd__nor2_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12935_ _12935_/A vssd1 vssd1 vccd1 vccd1 _12936_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _18442_/A vssd1 vssd1 vccd1 vccd1 _18443_/A sky130_fd_sc_hd__buf_2
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _16677_/B _16677_/C vssd1 vssd1 vccd1 vccd1 _15774_/A sky130_fd_sc_hd__nand2_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _12728_/B _12855_/Y _21065_/A _21174_/B _12852_/Y vssd1 vssd1 vccd1 vccd1
+ _12867_/C sky130_fd_sc_hd__o2111ai_4
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _23360_/Q vssd1 vssd1 vccd1 vccd1 _14883_/C sky130_fd_sc_hd__clkbuf_4
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _18373_/A vssd1 vssd1 vccd1 vccd1 _18376_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11817_ _12297_/A _12297_/D vssd1 vssd1 vccd1 vccd1 _12287_/C sky130_fd_sc_hd__nand2_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15585_ _23511_/Q _23512_/Q _23513_/Q _15585_/D vssd1 vssd1 vccd1 vccd1 _15586_/A
+ sky130_fd_sc_hd__or4_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _20957_/A _12796_/X _12703_/X _12706_/Y vssd1 vssd1 vccd1 vccd1 _12812_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_109_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17391_/C vssd1 vssd1 vccd1 vccd1 _17324_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14536_ _23040_/D vssd1 vssd1 vccd1 vccd1 _14657_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _11745_/A _11618_/C _11606_/X _11828_/B _11743_/A vssd1 vssd1 vccd1 vccd1
+ _11789_/B sky130_fd_sc_hd__o311ai_4
XFILLER_30_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17255_ _19381_/B vssd1 vssd1 vccd1 vccd1 _19694_/A sky130_fd_sc_hd__buf_4
X_14467_ _14464_/Y _14465_/X _14461_/X _14463_/Y vssd1 vssd1 vccd1 vccd1 _14478_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_186_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11679_ _23583_/Q vssd1 vssd1 vccd1 vccd1 _11724_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16551__A3 _16364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16206_ _15907_/B _15902_/Y _15910_/X _15899_/X vssd1 vssd1 vccd1 vccd1 _16206_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_174_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13418_ _13418_/A vssd1 vssd1 vccd1 vccd1 _13431_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17186_ _17186_/A vssd1 vssd1 vccd1 vccd1 _17187_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11579__B _16815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14398_ _14381_/A _14381_/B _14457_/A _14388_/X _14806_/A vssd1 vssd1 vccd1 vccd1
+ _14400_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_992 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _16860_/A _17098_/C _16308_/C _16634_/C vssd1 vssd1 vccd1 vccd1 _16137_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__13484__B1_N _13264_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13349_ _13394_/A vssd1 vssd1 vccd1 vccd1 _13349_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16451__A _16458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15993__C _17450_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22172__B _22392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16068_ _19659_/C vssd1 vssd1 vccd1 vccd1 _19199_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_170_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15019_ _15019_/A vssd1 vssd1 vccd1 vccd1 _15265_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__20399__A1 _20371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16601__D _18859_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17264__A1 _17610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19827_ _19827_/A vssd1 vssd1 vccd1 vccd1 _19939_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19758_ _19554_/X _19534_/D _19532_/X vssd1 vssd1 vccd1 vccd1 _19758_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19556__A3 _19358_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18709_ _18717_/C _18709_/B _18709_/C vssd1 vssd1 vccd1 vccd1 _18902_/A sky130_fd_sc_hd__nand3b_1
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19689_ _19796_/A _19796_/B vssd1 vssd1 vccd1 vccd1 _19740_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18764__A1 _12378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21720_ _21705_/X _21679_/X _23577_/Q vssd1 vssd1 vccd1 vccd1 _21728_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__13315__A _21925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15233__C _15233_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__22628__A _22628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21651_ _21631_/Y _21694_/C _21665_/A vssd1 vssd1 vccd1 vccd1 _21654_/A sky130_fd_sc_hd__a21o_1
XFILLER_36_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22848__B1 _22858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18516__A1 _12353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20602_ _20607_/A _20605_/A _20605_/B vssd1 vssd1 vccd1 vccd1 _20608_/B sky130_fd_sc_hd__nand3b_1
XFILLER_21_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21582_ _21570_/A _21569_/Y _21614_/C vssd1 vssd1 vccd1 vccd1 _21631_/B sky130_fd_sc_hd__o21a_1
XFILLER_71_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23321_ _23321_/CLK _23321_/D vssd1 vssd1 vccd1 vccd1 _23321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20533_ _20533_/A _20533_/B vssd1 vssd1 vccd1 vccd1 _20533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13050__A _13052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23252_ _23444_/Q input30/X _23254_/S vssd1 vssd1 vccd1 vccd1 _23253_/A sky130_fd_sc_hd__mux2_1
X_20464_ _20464_/A _20464_/B _20464_/C _20464_/D vssd1 vssd1 vccd1 vccd1 _20465_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_193_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18819__A2 _12006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22203_ _22203_/A _22203_/B vssd1 vssd1 vccd1 vccd1 _22203_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13985__A _15251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23183_ _23183_/A vssd1 vssd1 vccd1 vccd1 _23413_/D sky130_fd_sc_hd__clkbuf_1
X_20395_ _20420_/A _20395_/B vssd1 vssd1 vccd1 vccd1 _23535_/D sky130_fd_sc_hd__xnor2_1
XFILLER_3_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22134_ _22521_/A _22476_/C _22521_/C vssd1 vssd1 vccd1 vccd1 _22135_/B sky130_fd_sc_hd__and3_1
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22065_ _22173_/A vssd1 vssd1 vccd1 vccd1 _22167_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_0_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21016_ _21012_/X _21006_/Y _21015_/X vssd1 vssd1 vccd1 vccd1 _21243_/B sky130_fd_sc_hd__a21o_1
XFILLER_102_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22967_ _22967_/A vssd1 vssd1 vccd1 vccd1 _23317_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15018__B1 _15225_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13225__A _13732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ _12652_/X _12651_/X _12654_/Y _12661_/B vssd1 vssd1 vccd1 vccd1 _12734_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_21918_ _21934_/A _21918_/B _21934_/B vssd1 vssd1 vccd1 vccd1 _21939_/B sky130_fd_sc_hd__nand3_1
X_22898_ _22966_/S vssd1 vssd1 vccd1 vccd1 _22907_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_167_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18735__B _19280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20984__C _20984_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16230__A2 _16741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12651_ _12728_/A vssd1 vssd1 vccd1 vccd1 _12651_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21849_ _21852_/A _23482_/Q vssd1 vssd1 vccd1 vccd1 _21850_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18507__A1 _12460_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11602_ _18653_/C vssd1 vssd1 vccd1 vccd1 _11773_/C sky130_fd_sc_hd__buf_2
XFILLER_90_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21161__B _21271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15370_ _15370_/A vssd1 vssd1 vccd1 vccd1 _15446_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12582_ _23287_/Q vssd1 vssd1 vccd1 vccd1 _12618_/A sky130_fd_sc_hd__buf_2
XANTENNA__17715__C1 _19957_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14321_ _14911_/C vssd1 vssd1 vccd1 vccd1 _15253_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_183_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19847__A _20320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23519_ _23566_/CLK _23519_/D vssd1 vssd1 vccd1 vccd1 _23519_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_183_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17040_ _17040_/A vssd1 vssd1 vccd1 vccd1 _20317_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_128_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14252_ _14858_/A _14806_/C _15116_/B _14252_/D vssd1 vssd1 vccd1 vccd1 _14361_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__15741__A1 _16798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18470__B _18997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13203_ _13203_/A vssd1 vssd1 vccd1 vccd1 _13203_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13895__A _23504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14183_ _14183_/A vssd1 vssd1 vccd1 vccd1 _15175_/C sky130_fd_sc_hd__buf_2
XFILLER_87_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19483__A2 _19190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23521__CLK _23582_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13134_ _13133_/D _13133_/A _13151_/A _12785_/X vssd1 vssd1 vccd1 vccd1 _13135_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_98_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18991_ _18792_/Y _18806_/B _18796_/X _18790_/X vssd1 vssd1 vccd1 vccd1 _19186_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ _17942_/A _23529_/Q _17942_/C vssd1 vssd1 vccd1 vccd1 _18144_/B sky130_fd_sc_hd__nand3_2
X_13065_ _13063_/Y _13064_/Y _13061_/Y vssd1 vssd1 vccd1 vccd1 _13065_/Y sky130_fd_sc_hd__a21oi_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12016_ _12016_/A _12016_/B vssd1 vssd1 vccd1 vccd1 _12016_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17873_ _17773_/A _17758_/Y _17869_/Y _17872_/Y vssd1 vssd1 vccd1 vccd1 _17873_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19612_ _19614_/A _20371_/B _19614_/B _19381_/X vssd1 vssd1 vccd1 vccd1 _19612_/X
+ sky130_fd_sc_hd__a31o_1
X_16824_ _16447_/Y _16146_/A _16627_/A _16810_/A _16814_/A vssd1 vssd1 vccd1 vccd1
+ _16824_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_94_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19543_ _19543_/A _19543_/B _19811_/A _19709_/A vssd1 vssd1 vccd1 vccd1 _19543_/Y
+ sky130_fd_sc_hd__nand4_1
X_16755_ _16755_/A _16755_/B vssd1 vssd1 vccd1 vccd1 _16755_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13967_ _13948_/X _14029_/A _13908_/C vssd1 vssd1 vccd1 vccd1 _13972_/A sky130_fd_sc_hd__o21ai_1
XFILLER_59_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20002__B1 _19888_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15706_ _15706_/A _15707_/B _16591_/C _16591_/D vssd1 vssd1 vccd1 vccd1 _15908_/B
+ sky130_fd_sc_hd__nand4_4
X_19474_ _19470_/Y _19471_/Y _19472_/Y _19473_/Y vssd1 vssd1 vccd1 vccd1 _19592_/A
+ sky130_fd_sc_hd__o22ai_1
X_12918_ _20773_/D vssd1 vssd1 vccd1 vccd1 _21268_/A sky130_fd_sc_hd__buf_2
X_16686_ _16686_/A vssd1 vssd1 vccd1 vccd1 _17230_/A sky130_fd_sc_hd__clkbuf_4
X_13898_ _23352_/Q _23350_/Q _23351_/Q _14011_/B vssd1 vssd1 vccd1 vccd1 _13901_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_62_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18425_ _18407_/A _18407_/B _18407_/D _18424_/Y vssd1 vssd1 vccd1 vccd1 _18425_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_185_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15637_ _15761_/A _16187_/C _15637_/C _15637_/D vssd1 vssd1 vccd1 vccd1 _15639_/A
+ sky130_fd_sc_hd__nand4_4
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _12849_/A vssd1 vssd1 vccd1 vccd1 _12862_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22167__B _22479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18356_ _18356_/A _18356_/B vssd1 vssd1 vccd1 vccd1 _18394_/A sky130_fd_sc_hd__nand2_1
XANTENNA__21071__B _21276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15980__A1 _15889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15568_ _15574_/A vssd1 vssd1 vccd1 vccd1 _15569_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17307_ _17307_/A _17307_/B vssd1 vssd1 vccd1 vccd1 _17307_/Y sky130_fd_sc_hd__nand2_2
XFILLER_30_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14519_ _14633_/A _14633_/B _14633_/C _14519_/D vssd1 vssd1 vccd1 vccd1 _14551_/A
+ sky130_fd_sc_hd__and4bb_1
X_18287_ _18288_/A _18288_/B _18288_/C vssd1 vssd1 vccd1 vccd1 _18345_/A sky130_fd_sc_hd__a21o_1
XFILLER_119_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15499_ _15499_/A _15499_/B vssd1 vssd1 vccd1 vccd1 _15501_/C sky130_fd_sc_hd__xnor2_1
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17238_ _17238_/A _17238_/B _17238_/C vssd1 vssd1 vccd1 vccd1 _17246_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13301__C _22558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17169_ _17350_/A _17170_/B _17170_/C vssd1 vssd1 vccd1 vccd1 _17169_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_143_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20180_ _20171_/X _20179_/X _20173_/Y _20177_/Y vssd1 vssd1 vccd1 vccd1 _20180_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_143_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12214__A _12324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20241__B1 _20243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18985__A1 _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15525__A _15525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22821_ _22821_/A _22821_/B _22821_/C vssd1 vssd1 vccd1 vccd1 _22821_/Y sky130_fd_sc_hd__nand3_1
XFILLER_38_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13274__A2 _13732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14471__B2 _14469_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22752_ _22751_/X _22726_/B _22723_/B vssd1 vssd1 vccd1 vccd1 _22772_/A sky130_fd_sc_hd__a21oi_1
XFILLER_198_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21703_ _21700_/Y _21711_/A _21717_/B _21723_/A vssd1 vssd1 vccd1 vccd1 _23554_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22683_ _22683_/A _22683_/B vssd1 vssd1 vccd1 vccd1 _22683_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_515 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12884__A _20669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16356__A _16356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21634_ _21668_/B _21595_/B _21595_/C _21594_/A vssd1 vssd1 vccd1 vccd1 _21643_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_40_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16075__B _16075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1081 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11588__A2 _11960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21565_ _21565_/A _21565_/B vssd1 vssd1 vccd1 vccd1 _21566_/C sky130_fd_sc_hd__or2_1
XFILLER_139_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20516_ _20516_/A vssd1 vssd1 vccd1 vccd1 _20728_/A sky130_fd_sc_hd__clkbuf_2
X_23304_ _23336_/CLK _23304_/D vssd1 vssd1 vccd1 vccd1 _23304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21496_ _21559_/A _21559_/B vssd1 vssd1 vccd1 vccd1 _21509_/A sky130_fd_sc_hd__or2_1
XANTENNA__16920__B1 _16780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23235_ _23436_/Q input21/X _23239_/S vssd1 vssd1 vccd1 vccd1 _23236_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20447_ _20031_/X _20453_/B _23558_/Q vssd1 vssd1 vccd1 vccd1 _20448_/B sky130_fd_sc_hd__o21ai_1
XFILLER_181_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16279__A2 _16281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11947__B _16140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23166_ _23166_/A vssd1 vssd1 vccd1 vccd1 _23405_/D sky130_fd_sc_hd__clkbuf_1
X_20378_ _20378_/A _20378_/B vssd1 vssd1 vccd1 vccd1 _20379_/B sky130_fd_sc_hd__nand2_1
XFILLER_133_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22117_ _22106_/B _22439_/D _22118_/B _22117_/D vssd1 vssd1 vccd1 vccd1 _22117_/Y
+ sky130_fd_sc_hd__nand4b_1
XANTENNA__20480__B1 _14655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23097_ _23097_/A vssd1 vssd1 vccd1 vccd1 _23106_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17228__A1 _11971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20979__C _20984_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22048_ _21738_/C _13339_/X _14614_/X _21898_/B vssd1 vssd1 vccd1 vccd1 _22049_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_134_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14870_ _14868_/Y _14883_/B _14621_/X vssd1 vssd1 vccd1 vccd1 _14870_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_78_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13821_ _13552_/A _13599_/A _13610_/Y _13609_/X _13616_/Y vssd1 vssd1 vccd1 vccd1
+ _13821_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16540_ _16558_/A _16530_/A _16538_/Y _16539_/X vssd1 vssd1 vccd1 vccd1 _16540_/Y
+ sky130_fd_sc_hd__o22ai_1
X_13752_ _13744_/Y _13749_/Y _13751_/Y vssd1 vssd1 vccd1 vccd1 _13752_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12703_ _12622_/X _12624_/X _13151_/B vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__a21o_1
X_16471_ _16518_/C _16483_/B _16483_/A vssd1 vssd1 vccd1 vccd1 _16471_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13683_ _13544_/A _13303_/C _13303_/A vssd1 vssd1 vccd1 vccd1 _13864_/A sky130_fd_sc_hd__o21bai_1
XFILLER_188_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18210_ _18132_/B _18124_/Y _18155_/A _18155_/B vssd1 vssd1 vccd1 vccd1 _18210_/Y
+ sky130_fd_sc_hd__a22oi_4
X_15422_ _15422_/A _15427_/A _15420_/Y _15421_/X vssd1 vssd1 vccd1 vccd1 _15424_/B
+ sky130_fd_sc_hd__or4bb_1
X_19190_ _19190_/A vssd1 vssd1 vccd1 vccd1 _19668_/A sky130_fd_sc_hd__buf_2
XANTENNA__12225__B1 _12227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12634_ _12709_/A vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__buf_2
XFILLER_169_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18141_ _18141_/A _23531_/Q _18141_/C vssd1 vssd1 vccd1 vccd1 _18263_/B sky130_fd_sc_hd__and3_1
XFILLER_180_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15353_ _15353_/A _15353_/B _15353_/C vssd1 vssd1 vccd1 vccd1 _15353_/X sky130_fd_sc_hd__and3_1
XFILLER_169_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12565_ _19090_/A _12565_/B _12565_/C vssd1 vssd1 vccd1 vccd1 _12565_/X sky130_fd_sc_hd__and3_2
XFILLER_54_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater159_A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14304_ _14310_/B _14304_/B vssd1 vssd1 vccd1 vccd1 _14306_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18072_ _18072_/A _18072_/B _18072_/C _18072_/D vssd1 vssd1 vccd1 vccd1 _18072_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_102_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15284_ _15211_/B _15282_/Y _15392_/A _15392_/B vssd1 vssd1 vccd1 vccd1 _15395_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_89_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12496_ _12181_/A _12181_/B _12181_/C _12211_/C vssd1 vssd1 vccd1 vccd1 _18559_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17023_ _16979_/A _16979_/B _16979_/C vssd1 vssd1 vccd1 vccd1 _17024_/A sky130_fd_sc_hd__a21o_1
X_14235_ _14235_/A _14235_/B vssd1 vssd1 vccd1 vccd1 _14236_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14514__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output88_A _23582_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ _14162_/B _14331_/C _14331_/A _14167_/A _14167_/D vssd1 vssd1 vccd1 vccd1
+ _14166_/X sky130_fd_sc_hd__a32o_1
XFILLER_113_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11751__A2 _16360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _13114_/X _13115_/X _13116_/Y vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__a21bo_1
XFILLER_152_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _14097_/A vssd1 vssd1 vccd1 vccd1 _14097_/X sky130_fd_sc_hd__buf_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _11736_/A _18490_/A _18984_/B vssd1 vssd1 vccd1 vccd1 _18975_/A sky130_fd_sc_hd__o21ai_2
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23038__S _23038_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17925_ _17924_/C _17922_/A _17814_/B vssd1 vssd1 vccd1 vccd1 _17925_/Y sky130_fd_sc_hd__o21ai_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16690__A2 _15655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13048_ _13048_/A _13048_/B _13048_/C vssd1 vssd1 vccd1 vccd1 _13049_/A sky130_fd_sc_hd__nand3_1
XFILLER_140_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17856_ _17980_/A _17465_/X _17982_/A _17988_/A vssd1 vssd1 vccd1 vccd1 _17857_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16807_ _16807_/A _16807_/B vssd1 vssd1 vccd1 vccd1 _17434_/A sky130_fd_sc_hd__nand2_4
XANTENNA__16442__A2 _12373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_607 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17787_ _12237_/X _16742_/A _17646_/X _17407_/Y _17406_/Y vssd1 vssd1 vccd1 vccd1
+ _17788_/B sky130_fd_sc_hd__o32a_1
X_14999_ _15096_/A _15096_/B vssd1 vssd1 vccd1 vccd1 _14999_/Y sky130_fd_sc_hd__nand2_2
XFILLER_35_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19526_ _19526_/A _19526_/B _19578_/A _19578_/B vssd1 vssd1 vccd1 vccd1 _19526_/Y
+ sky130_fd_sc_hd__nand4_2
X_16738_ _16725_/Y _16737_/Y _16721_/Y _16724_/X vssd1 vssd1 vccd1 vccd1 _16739_/C
+ sky130_fd_sc_hd__o22ai_1
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19457_ _19457_/A _23544_/Q _19457_/C vssd1 vssd1 vccd1 vccd1 _19457_/X sky130_fd_sc_hd__and3_1
X_16669_ _16669_/A _16669_/B vssd1 vssd1 vccd1 vccd1 _17134_/C sky130_fd_sc_hd__nand2_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_824 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18408_ _18406_/Y _18408_/B vssd1 vssd1 vccd1 vccd1 _18409_/A sky130_fd_sc_hd__and2b_1
XFILLER_167_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19388_ _19573_/A _19573_/B _19568_/A _19569_/A vssd1 vssd1 vccd1 vccd1 _19389_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__13413__C1 _22388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19144__A1 _18944_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18339_ _18339_/A _18339_/B _18339_/C vssd1 vssd1 vccd1 vccd1 _18341_/A sky130_fd_sc_hd__nand3_1
XFILLER_33_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20829__A2 _12815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19695__A2 _17846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21350_ _21246_/X _21247_/X _21345_/C _21256_/Y vssd1 vssd1 vccd1 vccd1 _21350_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_135_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16363__D1 _16462_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__A1 _12374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20301_ _20293_/X _20294_/X _20343_/A vssd1 vssd1 vccd1 vccd1 _20301_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_163_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12519__B2 _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21281_ _21281_/A vssd1 vssd1 vccd1 vccd1 _21432_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23020_ _23020_/A vssd1 vssd1 vccd1 vccd1 _23340_/D sky130_fd_sc_hd__clkbuf_1
X_20232_ _20232_/A vssd1 vssd1 vccd1 vccd1 _20232_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_815 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1014 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20163_ _20217_/B vssd1 vssd1 vccd1 vccd1 _20269_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_104_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20094_ _20095_/A _20078_/A _20095_/C vssd1 vssd1 vccd1 vccd1 _20096_/B sky130_fd_sc_hd__a21o_1
XANTENNA__17454__B _17454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17630__A1 _17410_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11933__D _18531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22804_ _22756_/A _22764_/B _22829_/A _22829_/B vssd1 vssd1 vccd1 vccd1 _22840_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_77_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20996_ _21000_/A _21000_/B _20997_/A _21131_/B vssd1 vssd1 vccd1 vccd1 _20996_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22088__A _22089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12110__C _19193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22735_ _22698_/Y _22731_/Y _22810_/B vssd1 vssd1 vccd1 vccd1 _22738_/A sky130_fd_sc_hd__o21ba_1
XFILLER_198_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16086__A _19363_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_98 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22666_ _22725_/A _22670_/C _22237_/A _22484_/X vssd1 vssd1 vccd1 vccd1 _22666_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_185_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14318__B _15120_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21617_ _21617_/A vssd1 vssd1 vccd1 vccd1 _21617_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22597_ _22549_/A _22549_/B _22598_/A _22676_/A vssd1 vssd1 vccd1 vccd1 _22597_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_138_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12350_ _12372_/A _12372_/B vssd1 vssd1 vccd1 vccd1 _12350_/Y sky130_fd_sc_hd__nand2_1
X_21548_ _21668_/A _21548_/B _21637_/C _21548_/D vssd1 vssd1 vccd1 vccd1 _21548_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_194_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12281_ _12281_/A vssd1 vssd1 vccd1 vccd1 _12374_/A sky130_fd_sc_hd__buf_2
X_21479_ _21482_/B _21482_/C vssd1 vssd1 vccd1 vccd1 _21528_/B sky130_fd_sc_hd__nand2_1
XFILLER_153_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20055__B _20055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14020_ _14243_/A _14901_/A vssd1 vssd1 vccd1 vccd1 _14020_/Y sky130_fd_sc_hd__nand2_2
XFILLER_88_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23218_ _23218_/A vssd1 vssd1 vccd1 vccd1 _23428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17645__A _19670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_62 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23149_ _23149_/A vssd1 vssd1 vccd1 vccd1 _23397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15971_ _16598_/A vssd1 vssd1 vccd1 vccd1 _15971_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18949__A1 _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17710_ _17760_/A vssd1 vssd1 vccd1 vccd1 _17710_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14922_ _14926_/B _14926_/C _14926_/A vssd1 vssd1 vccd1 vccd1 _14922_/Y sky130_fd_sc_hd__a21oi_1
X_18690_ _18784_/B vssd1 vssd1 vccd1 vccd1 _18773_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_979 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17641_ _17641_/A _17641_/B _17641_/C vssd1 vssd1 vccd1 vccd1 _17788_/A sky130_fd_sc_hd__nand3_1
X_14853_ _14853_/A _14853_/B vssd1 vssd1 vccd1 vccd1 _15065_/B sky130_fd_sc_hd__nand2_1
XFILLER_75_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18476__A _18476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17380__A _23525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13804_ _21927_/A _13804_/B vssd1 vssd1 vccd1 vccd1 _13804_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17572_ _17566_/X _17575_/A _17571_/Y vssd1 vssd1 vccd1 vccd1 _17583_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12446__B1 _19180_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14784_ _14180_/B _14180_/C _14180_/A vssd1 vssd1 vccd1 vccd1 _14784_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20508__A1 _20502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_10_0_bq_clk_i clkbuf_3_5_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 _23598_/CLK
+ sky130_fd_sc_hd__clkbuf_8
X_11996_ _12183_/A _12187_/A _19019_/B _16027_/A vssd1 vssd1 vccd1 vccd1 _11996_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_189_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19311_ _19158_/A _19304_/X _19306_/X _19310_/Y vssd1 vssd1 vccd1 vccd1 _19320_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_95_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16523_ _16523_/A _16523_/B _16523_/C _16523_/D vssd1 vssd1 vccd1 vccd1 _16523_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_90_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13735_ _13563_/A _22192_/D _13563_/C _22192_/C _13736_/B vssd1 vssd1 vccd1 vccd1
+ _13735_/X sky130_fd_sc_hd__a32o_1
XFILLER_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14509__A _16167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19242_ _19410_/C _19146_/A _19241_/Y vssd1 vssd1 vccd1 vccd1 _19242_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_189_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16454_ _16404_/A _16405_/A _16452_/Y _16453_/X vssd1 vssd1 vccd1 vccd1 _16454_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_13666_ _13666_/A _13666_/B vssd1 vssd1 vccd1 vccd1 _13668_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19126__A1 _12184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15405_ _15350_/A _15353_/X _15352_/Y vssd1 vssd1 vccd1 vccd1 _15431_/A sky130_fd_sc_hd__a21boi_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _20493_/B vssd1 vssd1 vccd1 vccd1 _12667_/B sky130_fd_sc_hd__clkbuf_4
X_19173_ _11713_/A _11713_/B _19670_/B vssd1 vssd1 vccd1 vccd1 _19173_/X sky130_fd_sc_hd__a21o_2
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _17845_/C vssd1 vssd1 vccd1 vccd1 _17243_/D sky130_fd_sc_hd__buf_2
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13597_ _13538_/A _13538_/B _13477_/X vssd1 vssd1 vccd1 vccd1 _13598_/B sky130_fd_sc_hd__o21ai_1
X_18124_ _18133_/A vssd1 vssd1 vccd1 vccd1 _18124_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15336_ _15395_/A _15288_/B _15283_/X vssd1 vssd1 vccd1 vccd1 _15337_/B sky130_fd_sc_hd__a21oi_2
XFILLER_157_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12548_ _12547_/A _12303_/Y _12547_/B vssd1 vssd1 vccd1 vccd1 _12548_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16443__B _16499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18055_ _18198_/C _18140_/B _18054_/Y vssd1 vssd1 vccd1 vccd1 _18055_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15267_ _15388_/C _15267_/B _15267_/C _15420_/C vssd1 vssd1 vccd1 vccd1 _15267_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_144_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12479_ _18524_/B vssd1 vssd1 vccd1 vccd1 _12480_/B sky130_fd_sc_hd__clkinv_2
XFILLER_172_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11709__C1 _16619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17006_ _23519_/Q _17011_/A _17011_/B vssd1 vssd1 vccd1 vccd1 _17006_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_160_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14218_ _14218_/A _14218_/B _14218_/C vssd1 vssd1 vccd1 vccd1 _14218_/Y sky130_fd_sc_hd__nand3_2
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15198_ _15093_/B _15093_/A _15196_/X vssd1 vssd1 vccd1 vccd1 _15225_/A sky130_fd_sc_hd__a21o_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14149_ _14149_/A vssd1 vssd1 vccd1 vccd1 _14407_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_879 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16663__A2 _18461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18957_ _19123_/C vssd1 vssd1 vccd1 vccd1 _19900_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15075__A _15075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17908_ _17868_/Y _17873_/Y _17881_/Y _17902_/B vssd1 vssd1 vccd1 vccd1 _17909_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18888_ _18889_/A _18889_/B _18884_/Y _18885_/Y vssd1 vssd1 vccd1 vccd1 _18893_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20211__A3 _20320_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17839_ _17838_/B _17838_/C _17838_/A vssd1 vssd1 vccd1 vccd1 _18038_/C sky130_fd_sc_hd__a21oi_2
XFILLER_39_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20850_ _20733_/Y _20717_/A _20846_/Y _20849_/Y vssd1 vssd1 vccd1 vccd1 _20869_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18168__A2 _17753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19365__A1 _19218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19509_ _19509_/A vssd1 vssd1 vccd1 vccd1 _19868_/A sky130_fd_sc_hd__buf_2
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20781_ _20782_/A _20782_/B _20781_/C vssd1 vssd1 vccd1 vccd1 _20920_/A sky130_fd_sc_hd__nand3_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_790 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22520_ _22716_/D vssd1 vssd1 vccd1 vccd1 _22861_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__15926__A1 _12052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22451_ _22451_/A _22451_/B _22451_/C vssd1 vssd1 vccd1 vccd1 _22451_/Y sky130_fd_sc_hd__nand3_1
XFILLER_124_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19648__C _19652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16634__A _18755_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21402_ _21402_/A _21402_/B vssd1 vssd1 vccd1 vccd1 _21402_/Y sky130_fd_sc_hd__nand2_1
XFILLER_194_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13977__B _13977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22382_ _22386_/A _22386_/B _22384_/A _22283_/X vssd1 vssd1 vccd1 vccd1 _22393_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_198_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21333_ _21333_/A _21333_/B _21333_/C _21333_/D vssd1 vssd1 vccd1 vccd1 _21402_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_135_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19945__A _20142_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13165__A1 _20773_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21264_ _21354_/A vssd1 vssd1 vccd1 vccd1 _21264_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18628__B1 _18465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19664__B _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20215_ _20215_/A _20215_/B _20215_/C vssd1 vssd1 vccd1 vccd1 _20215_/X sky130_fd_sc_hd__and3_1
XANTENNA__12912__A1 _12902_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23003_ _23025_/A vssd1 vssd1 vccd1 vccd1 _23012_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__13993__A _23495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17465__A _17465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21195_ _21191_/Y _21192_/Y _21431_/C _21196_/A _21194_/Y vssd1 vssd1 vccd1 vccd1
+ _21195_/X sky130_fd_sc_hd__o2111a_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22090__B _22096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16800__C _23593_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20146_ _20146_/A _20146_/B _20146_/C _20146_/D vssd1 vssd1 vccd1 vccd1 _20148_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_132_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_998 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19053__B1 _18846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20077_ _19986_/B _20073_/X _20076_/X _20070_/Y _20172_/A vssd1 vssd1 vccd1 vccd1
+ _20078_/A sky130_fd_sc_hd__o2111ai_2
XANTENNA__12676__B1 _12675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12402__A _19011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12121__B _12121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _18500_/A _11848_/X _18474_/A vssd1 vssd1 vccd1 vccd1 _11850_/Y sky130_fd_sc_hd__o21ai_2
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19356__A1 _12378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11960__B _11960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11781_ _15718_/A vssd1 vssd1 vccd1 vccd1 _12262_/B sky130_fd_sc_hd__clkbuf_4
X_20979_ _20979_/A _20984_/B _20984_/C vssd1 vssd1 vccd1 vccd1 _20980_/C sky130_fd_sc_hd__nand3_1
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13520_ _13520_/A vssd1 vssd1 vccd1 vccd1 _13547_/A sky130_fd_sc_hd__buf_2
XFILLER_198_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22718_ _22722_/B vssd1 vssd1 vccd1 vccd1 _22718_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15917__A1 _11738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16244__A2_N _16254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13451_ _13257_/A _13269_/X _13450_/Y _13284_/Y vssd1 vssd1 vccd1 vccd1 _13516_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_186_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22649_ _22649_/A _22649_/B _22649_/C vssd1 vssd1 vccd1 vccd1 _22712_/A sky130_fd_sc_hd__nand3_2
XFILLER_139_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12402_ _19011_/A vssd1 vssd1 vccd1 vccd1 _19180_/D sky130_fd_sc_hd__buf_2
XANTENNA__14990__C _15094_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16170_ _16170_/A _16650_/A vssd1 vssd1 vccd1 vccd1 _16175_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_884 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13382_ _23473_/Q vssd1 vssd1 vccd1 vccd1 _21909_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15121_ _15121_/A vssd1 vssd1 vccd1 vccd1 _15164_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__20674__B1 _23454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12333_ _12339_/A _12339_/B vssd1 vssd1 vccd1 vccd1 _12334_/B sky130_fd_sc_hd__nand2_1
XFILLER_126_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15052_ _15049_/B _15052_/B _15052_/C vssd1 vssd1 vccd1 vccd1 _15053_/B sky130_fd_sc_hd__nand3b_1
X_12264_ _16049_/D vssd1 vssd1 vccd1 vccd1 _17134_/B sky130_fd_sc_hd__buf_4
XFILLER_123_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23262__CLK _23584_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14003_ _14003_/A _14253_/B vssd1 vssd1 vccd1 vccd1 _14003_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18095__B2 _20210_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19860_ _20081_/A _19482_/B _19953_/A _20210_/C _19674_/Y vssd1 vssd1 vccd1 vccd1
+ _19860_/X sky130_fd_sc_hd__o32a_1
X_12195_ _12211_/A _12206_/A _12196_/C vssd1 vssd1 vccd1 vccd1 _12199_/C sky130_fd_sc_hd__a21o_1
XFILLER_122_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput61 _14663_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput72 _14705_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[26] sky130_fd_sc_hd__buf_2
X_18811_ _23394_/Q _18811_/B _18811_/C vssd1 vssd1 vccd1 vccd1 _18812_/C sky130_fd_sc_hd__nand3b_2
Xoutput83 _14591_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[7] sky130_fd_sc_hd__buf_2
Xoutput94 _23268_/Q vssd1 vssd1 vccd1 vccd1 y[6] sky130_fd_sc_hd__buf_2
X_19791_ _19789_/Y _19791_/B vssd1 vssd1 vccd1 vccd1 _19792_/A sky130_fd_sc_hd__and2b_2
XFILLER_1_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_732 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18742_ _18739_/Y _18740_/Y _18741_/Y _18589_/Y _12567_/A vssd1 vssd1 vccd1 vccd1
+ _18747_/A sky130_fd_sc_hd__a32oi_4
X_15954_ _19364_/C _16821_/A _19364_/B vssd1 vssd1 vccd1 vccd1 _16119_/A sky130_fd_sc_hd__nand3_4
XFILLER_95_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12312__A _17149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14905_ _14058_/X _15366_/A _14872_/Y _14874_/A vssd1 vssd1 vccd1 vccd1 _14968_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18673_ _18673_/A vssd1 vssd1 vccd1 vccd1 _18673_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15885_ _15882_/X _15884_/X _15843_/A _15852_/X _15754_/X vssd1 vssd1 vccd1 vccd1
+ _15886_/C sky130_fd_sc_hd__o221ai_1
XFILLER_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17624_ _17460_/B _17457_/Y _17467_/X _17454_/Y vssd1 vssd1 vccd1 vccd1 _17637_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_14836_ _14298_/C _15054_/A _14007_/B _14835_/X vssd1 vssd1 vccd1 vccd1 _14836_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _17555_/A vssd1 vssd1 vccd1 vccd1 _17806_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__22159__C _22159_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14767_ _14783_/B vssd1 vssd1 vccd1 vccd1 _14857_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14239__A _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11979_ _18469_/D vssd1 vssd1 vccd1 vccd1 _18998_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_17_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_790 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16506_ _16440_/Y _16505_/Y _16463_/Y _16465_/Y vssd1 vssd1 vccd1 vccd1 _16507_/B
+ sky130_fd_sc_hd__a22oi_4
X_13718_ _21892_/A _13487_/Y _13482_/Y _13709_/A _13705_/D vssd1 vssd1 vccd1 vccd1
+ _13720_/C sky130_fd_sc_hd__o2111ai_1
X_17486_ _17654_/A _17654_/B _17481_/C _17481_/D vssd1 vssd1 vccd1 vccd1 _17486_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14698_ _14698_/A vssd1 vssd1 vccd1 vccd1 _14698_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19225_ _19148_/X _19151_/Y _19215_/Y _19224_/Y vssd1 vssd1 vccd1 vccd1 _19226_/A
+ sky130_fd_sc_hd__o211ai_4
X_16437_ _16437_/A vssd1 vssd1 vccd1 vccd1 _16437_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_72_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1068 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13649_ _13633_/X _13637_/X _13645_/A _13645_/B vssd1 vssd1 vccd1 vccd1 _13649_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_82_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19156_ _19156_/A _19156_/B _19156_/C vssd1 vssd1 vccd1 vccd1 _20369_/C sky130_fd_sc_hd__nand3_4
X_16368_ _16364_/X _16399_/A _12238_/A _16398_/A vssd1 vssd1 vccd1 vccd1 _16369_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__13797__B _13797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18107_ _18179_/B _18106_/C _18106_/A vssd1 vssd1 vccd1 vccd1 _18108_/B sky130_fd_sc_hd__a21o_1
XFILLER_145_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15319_ _15419_/C _15419_/D _15319_/C vssd1 vssd1 vccd1 vccd1 _15366_/C sky130_fd_sc_hd__nand3_1
X_19087_ _19087_/A _19087_/B _19087_/C _19263_/A vssd1 vssd1 vccd1 vccd1 _19088_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_184_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16299_ _16366_/A vssd1 vssd1 vccd1 vccd1 _16389_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18038_ _18038_/A _18123_/A _18038_/C vssd1 vssd1 vccd1 vccd1 _18043_/C sky130_fd_sc_hd__nand3_1
XFILLER_160_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20704__A _23457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18086__A1 _12506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17285__A _17285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20000_ _20003_/C _20003_/D vssd1 vssd1 vccd1 vccd1 _20000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16097__B1 _16335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16636__A2 _16370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19989_ _19850_/Y _19860_/X _19943_/B vssd1 vssd1 vccd1 vccd1 _19991_/B sky130_fd_sc_hd__o21ai_2
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20142__C _20142_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21951_ _21982_/A _22089_/A _21982_/B vssd1 vssd1 vccd1 vccd1 _21953_/B sky130_fd_sc_hd__nand3_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ _20902_/A _20902_/B _20902_/C vssd1 vssd1 vccd1 vccd1 _20903_/B sky130_fd_sc_hd__nand3_1
XFILLER_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21882_ _21882_/A _21882_/B _21882_/C vssd1 vssd1 vccd1 vccd1 _21884_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19338__A1 _19966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22069__C _22208_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20833_ _20841_/A _20841_/B vssd1 vssd1 vccd1 vccd1 _20843_/B sky130_fd_sc_hd__nand2_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18010__A1 _12088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23552_ _23558_/CLK _23552_/D vssd1 vssd1 vccd1 vccd1 _23552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19659__B _20047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20764_ _20608_/A _20608_/B _20608_/C _20611_/A vssd1 vssd1 vccd1 vccd1 _20765_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_126_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16021__B1 _16020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22503_ _13803_/A _13803_/B _21829_/A vssd1 vssd1 vccd1 vccd1 _22505_/B sky130_fd_sc_hd__a21o_1
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23483_ _23499_/CLK _23495_/Q vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20695_ _20695_/A _20695_/B _20695_/C vssd1 vssd1 vccd1 vccd1 _20711_/A sky130_fd_sc_hd__nand3_1
XFILLER_196_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16364__A _16364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_862 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22434_ _22434_/A _22457_/A _22524_/A _22434_/D vssd1 vssd1 vccd1 vccd1 _22435_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_149_884 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20317__C _20317_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19675__A _19675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22365_ _22508_/A _22508_/B _22365_/C vssd1 vssd1 vccd1 vccd1 _22365_/X sky130_fd_sc_hd__and3_1
XFILLER_184_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21316_ _21306_/A _21307_/D _21315_/X vssd1 vssd1 vccd1 vccd1 _21317_/D sky130_fd_sc_hd__a21o_1
XANTENNA__23197__A _23254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22296_ _22476_/A _22476_/B _22562_/B vssd1 vssd1 vccd1 vccd1 _22297_/B sky130_fd_sc_hd__nand3_2
XFILLER_190_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21247_ _21353_/A vssd1 vssd1 vccd1 vccd1 _21247_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21178_ _21281_/A _21282_/A _21178_/C _21279_/D vssd1 vssd1 vccd1 vccd1 _21179_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14638__A1 _14632_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_946 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20129_ _20102_/A _20102_/B _20111_/C vssd1 vssd1 vccd1 vccd1 _20183_/A sky130_fd_sc_hd__o21a_1
XFILLER_133_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19841__C _19949_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21908__B1 _22043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12951_ _12640_/X _12637_/X _12696_/A _12724_/A vssd1 vssd1 vccd1 vccd1 _12952_/A
+ sky130_fd_sc_hd__o211ai_2
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_34 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17052__A2 _17975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _11902_/A _11902_/B _11902_/C vssd1 vssd1 vccd1 vccd1 _11912_/D sky130_fd_sc_hd__nand3_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15670_ _12373_/A _15802_/B _15655_/X _15669_/X _15641_/Y vssd1 vssd1 vccd1 vccd1
+ _15670_/X sky130_fd_sc_hd__o311a_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12882_ _20894_/A _12756_/B _12875_/B vssd1 vssd1 vccd1 vccd1 _12882_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _23362_/Q vssd1 vssd1 vccd1 vccd1 _14621_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ _11745_/A _23382_/Q _11656_/B _11608_/A _11746_/A vssd1 vssd1 vccd1 vccd1
+ _11834_/B sky130_fd_sc_hd__o311ai_4
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17334_/A _17334_/B _17350_/B _17339_/X vssd1 vssd1 vccd1 vccd1 _17341_/C
+ sky130_fd_sc_hd__a31oi_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _23184_/D vssd1 vssd1 vccd1 vccd1 _14698_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12821__B1 _12770_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ _11764_/A vssd1 vssd1 vccd1 vccd1 _11868_/A sky130_fd_sc_hd__buf_2
XFILLER_198_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22276__A _22276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ _13450_/Y _13496_/X _22392_/C _13712_/D _13502_/X vssd1 vssd1 vccd1 vccd1
+ _13507_/A sky130_fd_sc_hd__o2111a_1
XFILLER_53_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17271_ _16447_/Y _17744_/A _17433_/A vssd1 vssd1 vccd1 vccd1 _17271_/X sky130_fd_sc_hd__o21a_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18488__A1_N _18458_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14483_ _14483_/A _14486_/C _14486_/B _14486_/A vssd1 vssd1 vccd1 vccd1 _14483_/Y
+ sky130_fd_sc_hd__nand4_1
X_11695_ _11808_/A _23587_/Q vssd1 vssd1 vccd1 vccd1 _11695_/X sky130_fd_sc_hd__and2_1
XFILLER_158_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19010_ _19010_/A vssd1 vssd1 vccd1 vccd1 _19700_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16222_ _16222_/A _16233_/A vssd1 vssd1 vccd1 vccd1 _16222_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16705__C _16706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13434_ _13434_/A _13434_/B vssd1 vssd1 vccd1 vccd1 _13434_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16153_ _16153_/A _16153_/B vssd1 vssd1 vccd1 vccd1 _16590_/A sky130_fd_sc_hd__nand2_2
XFILLER_154_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13365_ _13323_/X _13338_/X _13354_/C _13354_/B _13366_/B vssd1 vssd1 vccd1 vccd1
+ _13365_/Y sky130_fd_sc_hd__a41oi_4
XFILLER_154_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15104_ _15104_/A vssd1 vssd1 vccd1 vccd1 _15419_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_bq_clk_i clkbuf_0_bq_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_12316_ _17134_/B vssd1 vssd1 vccd1 vccd1 _16549_/B sky130_fd_sc_hd__buf_2
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16084_ _16084_/A _16084_/B _16084_/C vssd1 vssd1 vccd1 vccd1 _16297_/B sky130_fd_sc_hd__nand3_2
X_13296_ _21882_/B vssd1 vssd1 vccd1 vccd1 _22363_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14877__A1 _14883_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_846 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19912_ _19771_/X _19794_/Y _19911_/Y vssd1 vssd1 vccd1 vccd1 _19925_/A sky130_fd_sc_hd__o21bai_1
X_15035_ _15035_/A _15035_/B _15077_/B _15035_/D vssd1 vssd1 vccd1 vccd1 _15036_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19265__B1 _12353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ _11676_/X _11980_/B _11999_/A _11840_/X _12245_/X vssd1 vssd1 vccd1 vccd1
+ _12247_/Y sky130_fd_sc_hd__a311oi_4
XANTENNA__14522__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20243__B _20243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output70_A _14697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__A2 _11931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19843_ _19949_/A _20142_/C _19848_/B vssd1 vssd1 vccd1 vccd1 _19843_/Y sky130_fd_sc_hd__nand3_1
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12178_ _15882_/A _12171_/Y _12177_/Y vssd1 vssd1 vccd1 vccd1 _12178_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_150_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14629__A1 _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15826__B1 _12020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19774_ _19442_/Y _19443_/Y _19275_/Y _19773_/X vssd1 vssd1 vccd1 vccd1 _19774_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16986_ _17025_/A _16982_/X _16994_/D vssd1 vssd1 vccd1 vccd1 _17374_/C sky130_fd_sc_hd__o21ai_2
XFILLER_114_1050 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18725_ _18728_/A _18728_/B _18725_/C _18725_/D vssd1 vssd1 vccd1 vccd1 _19091_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_7_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15937_ _15937_/A vssd1 vssd1 vccd1 vccd1 _17625_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_595 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15353__A _15353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15868_ _15868_/A vssd1 vssd1 vccd1 vccd1 _19703_/B sky130_fd_sc_hd__buf_2
X_18656_ _12004_/X _12006_/X _20046_/A _20047_/A vssd1 vssd1 vccd1 vccd1 _18656_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_97_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18791__A2 _18484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17607_ _17243_/D _20138_/A _20138_/B _18077_/A _17243_/B vssd1 vssd1 vccd1 vccd1
+ _17607_/X sky130_fd_sc_hd__a32o_1
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14819_ _14819_/A _23504_/Q vssd1 vssd1 vccd1 vccd1 _14821_/C sky130_fd_sc_hd__nand2_1
XFILLER_92_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13065__B1 _13061_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18587_ _18576_/A _18570_/Y _18573_/Y vssd1 vssd1 vccd1 vccd1 _18733_/C sky130_fd_sc_hd__o21ai_2
XFILLER_17_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15799_ _15799_/A vssd1 vssd1 vccd1 vccd1 _17414_/D sky130_fd_sc_hd__buf_4
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17538_ _17934_/A vssd1 vssd1 vccd1 vccd1 _17538_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18543__A2 _18541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17469_ _17469_/A vssd1 vssd1 vccd1 vccd1 _17473_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__15800__B _17414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13368__A1 _13349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19208_ _19194_/X _19196_/Y _19207_/X vssd1 vssd1 vccd1 vccd1 _19221_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20480_ _12748_/X _20479_/X _14655_/A _20494_/D vssd1 vssd1 vccd1 vccd1 _20482_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_146_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19139_ _19139_/A _19139_/B vssd1 vssd1 vccd1 vccd1 _19140_/C sky130_fd_sc_hd__nand2_1
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22150_ _22144_/A _22168_/A _22144_/C _22141_/D _13486_/B vssd1 vssd1 vccd1 vccd1
+ _22150_/Y sky130_fd_sc_hd__a41oi_4
XFILLER_173_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21101_ _21101_/A _21101_/B _21101_/C vssd1 vssd1 vccd1 vccd1 _21101_/Y sky130_fd_sc_hd__nand3_1
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16719__A2_N _16176_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22081_ _22076_/X _22077_/Y _22069_/Y _22074_/X vssd1 vssd1 vccd1 vccd1 _22083_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_160_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21032_ _21025_/A _21029_/X _21031_/Y vssd1 vssd1 vccd1 vccd1 _21147_/A sky130_fd_sc_hd__o21ai_1
XFILLER_99_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19646__A2_N _16033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22983_ _22983_/A vssd1 vssd1 vccd1 vccd1 _23323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21934_ _21934_/A _21934_/B vssd1 vssd1 vccd1 vccd1 _21934_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_26 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21865_ _21861_/Y _21864_/Y _23270_/Q _21971_/B vssd1 vssd1 vccd1 vccd1 _21867_/A
+ sky130_fd_sc_hd__a211oi_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20816_ _20819_/C _20819_/D vssd1 vssd1 vccd1 vccd1 _20817_/B sky130_fd_sc_hd__nand2_1
XFILLER_196_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21796_ _13826_/X _21795_/X _13818_/B vssd1 vssd1 vccd1 vccd1 _21798_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__22096__A _22830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18534__A2 _17456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23535_ _23558_/CLK _23535_/D vssd1 vssd1 vccd1 vccd1 _23535_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16545__A1 _16531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20747_ _20868_/A _20867_/A _20747_/C vssd1 vssd1 vccd1 vccd1 _20748_/C sky130_fd_sc_hd__nand3_1
XFILLER_184_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13359__A1 _23325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22618__B2 _22858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23466_ _23571_/CLK _23478_/Q vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfxtp_1
X_20678_ _20678_/A _20678_/B vssd1 vssd1 vccd1 vccd1 _20678_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15918__A_N _15921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22417_ _22417_/A _22417_/B _22417_/C vssd1 vssd1 vccd1 vccd1 _22428_/D sky130_fd_sc_hd__nand3_1
XANTENNA__12031__A1 _12051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23397_ _23397_/CLK _23397_/D vssd1 vssd1 vccd1 vccd1 _23397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16848__A2 _18607_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ _13172_/A _13172_/B _13172_/C vssd1 vssd1 vccd1 vccd1 _13171_/A sky130_fd_sc_hd__a21oi_1
X_22348_ _21973_/C _22348_/B _22348_/C _22348_/D vssd1 vssd1 vccd1 vccd1 _22348_/Y
+ sky130_fd_sc_hd__nand4b_1
XFILLER_151_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12101_ _18447_/B vssd1 vssd1 vccd1 vccd1 _19193_/C sky130_fd_sc_hd__buf_2
XFILLER_128_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__23043__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12246__B1_N _12245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13081_ _13072_/Y _13075_/Y _20595_/B vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__o21ai_1
X_22279_ _22279_/A _22386_/A vssd1 vssd1 vccd1 vccd1 _22279_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__19798__A1 _19203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_762 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19798__B2 _19218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ _12032_/A _12032_/B vssd1 vssd1 vccd1 vccd1 _12159_/C sky130_fd_sc_hd__nand2_1
XFILLER_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16840_ _16840_/A _18755_/D _18755_/C vssd1 vssd1 vccd1 vccd1 _16841_/B sky130_fd_sc_hd__and3_1
XFILLER_66_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16481__B1 _16479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16771_ _16771_/A _16771_/B _16771_/C vssd1 vssd1 vccd1 vccd1 _17010_/C sky130_fd_sc_hd__nand3_1
XFILLER_19_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13983_ _23502_/Q _23501_/Q vssd1 vssd1 vccd1 vccd1 _15251_/A sky130_fd_sc_hd__and2_1
XFILLER_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18510_ _18511_/A _18511_/B _18510_/C _18510_/D vssd1 vssd1 vccd1 vccd1 _18518_/A
+ sky130_fd_sc_hd__nand4_2
X_15722_ _11868_/A _16200_/A _15908_/A _15908_/B _15721_/X vssd1 vssd1 vccd1 vccd1
+ _15723_/C sky130_fd_sc_hd__o221ai_4
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11845__A1 _12353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12934_ _13113_/A _13113_/C _12933_/X vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__18222__B2 _18330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19490_ _19670_/C _19480_/X _19847_/C _19482_/Y _20062_/B vssd1 vssd1 vccd1 vccd1
+ _19492_/B sky130_fd_sc_hd__o2111ai_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ _18439_/X _18440_/X _18788_/A vssd1 vssd1 vccd1 vccd1 _18442_/A sky130_fd_sc_hd__o21ai_1
XFILLER_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_727 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23450__CLK _23462_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15653_ _15621_/X _15618_/X _16661_/C _16866_/A vssd1 vssd1 vccd1 vccd1 _15802_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__B _22035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12865_ _21039_/B vssd1 vssd1 vccd1 vccd1 _21174_/B sky130_fd_sc_hd__buf_2
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18484__A _18484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14604_ _23424_/Q vssd1 vssd1 vccd1 vccd1 _15605_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _23536_/Q vssd1 vssd1 vccd1 vccd1 _18398_/A sky130_fd_sc_hd__inv_2
X_11816_ _11717_/B _11717_/C _12238_/A _11815_/X vssd1 vssd1 vccd1 vccd1 _12297_/D
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15584_ _23513_/Q _15584_/B vssd1 vssd1 vccd1 vccd1 _23501_/D sky130_fd_sc_hd__xor2_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12796_ _12796_/A vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__buf_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17391_/B vssd1 vssd1 vccd1 vccd1 _17323_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14535_ _14535_/A _14538_/B _14538_/C _14538_/A vssd1 vssd1 vccd1 vccd1 _23040_/D
+ sky130_fd_sc_hd__nor4b_2
XFILLER_57_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11789_/A vssd1 vssd1 vccd1 vccd1 _11747_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__15423__A1_N _15422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17254_ _17434_/A _17435_/A _17057_/A _18947_/A vssd1 vssd1 vccd1 vccd1 _17439_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_175_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14466_ _14461_/X _14463_/Y _14464_/Y _14465_/X vssd1 vssd1 vccd1 vccd1 _14468_/A
+ sky130_fd_sc_hd__a211o_1
X_11678_ _11686_/B _11676_/X _11677_/X vssd1 vssd1 vccd1 vccd1 _11852_/A sky130_fd_sc_hd__o21a_4
XANTENNA__18931__B _18931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16205_ _15902_/B _16202_/Y _16217_/B vssd1 vssd1 vccd1 vccd1 _16205_/Y sky130_fd_sc_hd__o21ai_1
X_13417_ _13417_/A _13423_/A vssd1 vssd1 vccd1 vccd1 _13418_/A sky130_fd_sc_hd__nand2_1
X_17185_ _16957_/A _16957_/B _17183_/Y _17184_/Y vssd1 vssd1 vccd1 vccd1 _17185_/Y
+ sky130_fd_sc_hd__a22oi_4
X_14397_ _14381_/B _14395_/B _14436_/A vssd1 vssd1 vccd1 vccd1 _14400_/A sky130_fd_sc_hd__o21ai_1
XFILLER_155_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16136_ _16136_/A vssd1 vssd1 vccd1 vccd1 _16174_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13348_ _21744_/C vssd1 vssd1 vccd1 vccd1 _13348_/X sky130_fd_sc_hd__buf_2
XFILLER_6_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16451__B _16451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_868 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16067_ _17041_/B vssd1 vssd1 vccd1 vccd1 _17248_/C sky130_fd_sc_hd__buf_2
XANTENNA__23034__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13279_ _13279_/A vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__buf_2
XANTENNA__14252__A _14858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15018_ _14243_/A _14901_/X _15254_/B _15225_/C _15253_/B vssd1 vssd1 vccd1 vccd1
+ _15020_/C sky130_fd_sc_hd__a32o_1
XFILLER_116_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22793__B1 _22237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19826_ _19835_/A _19836_/A _19825_/X _19673_/Y vssd1 vssd1 vccd1 vccd1 _19827_/A
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_151_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17264__A2 _17285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19757_ _19757_/A _19757_/B _19757_/C vssd1 vssd1 vccd1 vccd1 _19757_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__21348__A1 _21542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16969_ _17202_/A _16969_/B _16969_/C vssd1 vssd1 vccd1 vccd1 _16969_/X sky130_fd_sc_hd__and3_1
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18708_ _18708_/A _18708_/B vssd1 vssd1 vccd1 vccd1 _18709_/C sky130_fd_sc_hd__nand2_1
X_19688_ _19688_/A _19688_/B vssd1 vssd1 vccd1 vccd1 _19796_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12500__A _23593_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18764__A2 _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22909__A _22966_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18639_ _18639_/A _18639_/B vssd1 vssd1 vccd1 vccd1 _18639_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21650_ _21650_/A _21650_/B vssd1 vssd1 vccd1 vccd1 _21665_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_708 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18516__A2 _17643_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20601_ _20597_/C _20614_/A _20614_/B vssd1 vssd1 vccd1 vccd1 _20605_/B sky130_fd_sc_hd__nand3b_2
XFILLER_177_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12261__A1 _18673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21581_ _21616_/A _21617_/A _21529_/X _21575_/Y _21572_/Y vssd1 vssd1 vccd1 vccd1
+ _21625_/B sky130_fd_sc_hd__o221ai_1
XANTENNA__16527__A1 _12346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23320_ input5/X _23320_/D vssd1 vssd1 vccd1 vccd1 _23320_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13331__A _13660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20532_ _20532_/A _20532_/B _23455_/Q vssd1 vssd1 vccd1 vccd1 _20533_/B sky130_fd_sc_hd__and3_1
XFILLER_166_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22644__A _22644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20463_ _20612_/A _20613_/A vssd1 vssd1 vccd1 vccd1 _21018_/A sky130_fd_sc_hd__or2_1
X_23251_ _23251_/A vssd1 vssd1 vccd1 vccd1 _23443_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13050__B _23454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_256 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22202_ _22215_/A _22215_/B _22201_/Y vssd1 vssd1 vccd1 vccd1 _22207_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__21284__B1 _20957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20394_ _20420_/B _20394_/B vssd1 vssd1 vccd1 vccd1 _20395_/B sky130_fd_sc_hd__nand2_1
XFILLER_174_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23182_ _23413_/Q input31/X _23182_/S vssd1 vssd1 vccd1 vccd1 _23183_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22133_ _22123_/Y _22126_/X _22132_/X _22128_/Y vssd1 vssd1 vccd1 vccd1 _22136_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_134_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22064_ _22064_/A _22064_/B _22064_/C vssd1 vssd1 vccd1 vccd1 _22173_/A sky130_fd_sc_hd__nand3_1
XFILLER_82_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21015_ _21014_/X _21002_/Y _20999_/X vssd1 vssd1 vccd1 vccd1 _21015_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_1_0_bq_clk_i_A clkbuf_2_1_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_798 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22966_ _23317_/Q input31/X _22966_/S vssd1 vssd1 vccd1 vccd1 _22967_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15018__B2 _15253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21917_ _22487_/A _21750_/Y _22270_/C _21916_/Y vssd1 vssd1 vccd1 vccd1 _21934_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13225__B _13732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22897_ _22953_/A vssd1 vssd1 vccd1 vccd1 _22966_/S sky130_fd_sc_hd__buf_2
XFILLER_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12650_ _13121_/A _13121_/B _20781_/C vssd1 vssd1 vccd1 vccd1 _12728_/A sky130_fd_sc_hd__nand3_1
XFILLER_167_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21848_ _21852_/A _23482_/Q vssd1 vssd1 vccd1 vccd1 _21850_/A sky130_fd_sc_hd__or2_1
XFILLER_167_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18507__A2 _18503_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16536__B _16536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11601_ _23397_/Q vssd1 vssd1 vccd1 vccd1 _18653_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _20799_/A _13019_/C _13019_/B vssd1 vssd1 vccd1 vccd1 _20532_/A sky130_fd_sc_hd__o21ai_4
XFILLER_168_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21779_ _13616_/A _13616_/B _13620_/X vssd1 vssd1 vccd1 vccd1 _21779_/X sky130_fd_sc_hd__a21o_1
XFILLER_196_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14320_ _14911_/B vssd1 vssd1 vccd1 vccd1 _15017_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23518_ _23518_/CLK input43/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_196_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19847__B _20320_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22554__A _22554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ _14243_/A _14901_/A _14374_/D _14806_/C _14867_/C vssd1 vssd1 vccd1 vccd1
+ _14251_/Y sky130_fd_sc_hd__a32oi_4
XFILLER_172_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23449_ _23559_/CLK hold17/X vssd1 vssd1 vccd1 vccd1 _23449_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15741__A2 _14553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202_ _13202_/A vssd1 vssd1 vccd1 vccd1 _13208_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_87_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14182_ _14181_/X _14178_/Y _14177_/A vssd1 vssd1 vccd1 vccd1 _14187_/A sky130_fd_sc_hd__o21ai_1
XFILLER_178_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15168__A _15233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20483__D1 _21054_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13133_ _13133_/A _21548_/B _13133_/C _13133_/D vssd1 vssd1 vccd1 vccd1 _13196_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__18691__A1 _18673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18990_ _18971_/X _18981_/A _19509_/A _18975_/A _15928_/C vssd1 vssd1 vccd1 vccd1
+ _18992_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_151_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17941_ _18207_/A _18208_/A _18253_/A _18253_/B _17933_/X vssd1 vssd1 vccd1 vccd1
+ _17942_/C sky130_fd_sc_hd__o221ai_4
X_13064_ _13058_/Y _13059_/X _13051_/X vssd1 vssd1 vccd1 vccd1 _13064_/Y sky130_fd_sc_hd__o21ai_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18479__A _18479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12015_ _12011_/X _12013_/Y _12029_/B vssd1 vssd1 vccd1 vccd1 _12015_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_39_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17872_ _17874_/A _17874_/B _17867_/Y vssd1 vssd1 vccd1 vccd1 _17872_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_repeater104_A _23479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19611_ _20320_/A vssd1 vssd1 vccd1 vccd1 _20371_/B sky130_fd_sc_hd__clkbuf_2
X_16823_ _16814_/X _16821_/Y _16822_/X vssd1 vssd1 vccd1 vccd1 _16823_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19542_ _19542_/A vssd1 vssd1 vccd1 vccd1 _19542_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16754_ _16988_/A _16989_/A _16778_/A _16792_/A vssd1 vssd1 vccd1 vccd1 _16998_/C
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_98_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13966_ _13966_/A vssd1 vssd1 vccd1 vccd1 _13966_/X sky130_fd_sc_hd__buf_2
XFILLER_185_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12917_ _23456_/Q vssd1 vssd1 vccd1 vccd1 _20773_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15705_ _16187_/A _16187_/B _16187_/C _15688_/A vssd1 vssd1 vccd1 vccd1 _16591_/C
+ sky130_fd_sc_hd__a31o_2
X_19473_ _19471_/B _19470_/A _19471_/A vssd1 vssd1 vccd1 vccd1 _19473_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16685_ _16683_/X _16684_/X _15660_/A vssd1 vssd1 vccd1 vccd1 _16686_/A sky130_fd_sc_hd__o21ai_2
X_13897_ _23365_/Q vssd1 vssd1 vccd1 vccd1 _14011_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18424_ _18417_/A _18398_/C _18398_/A vssd1 vssd1 vccd1 vccd1 _18424_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12848_ _20473_/C _20473_/A vssd1 vssd1 vccd1 vccd1 _12849_/A sky130_fd_sc_hd__nand2_1
X_15636_ _23420_/Q _23421_/Q _23422_/Q vssd1 vssd1 vccd1 vccd1 _15637_/C sky130_fd_sc_hd__nor3_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18355_ _18355_/A _18355_/B vssd1 vssd1 vccd1 vccd1 _18356_/B sky130_fd_sc_hd__nor2_1
XFILLER_15_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15350__B _15353_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15567_ _15567_/A vssd1 vssd1 vccd1 vccd1 _23285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _12779_/A _12779_/B _12779_/C vssd1 vssd1 vccd1 vccd1 _12975_/B sky130_fd_sc_hd__nand3_2
XFILLER_187_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15980__A2 _15971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17306_ _16032_/X _16033_/X _17631_/A _17712_/D vssd1 vssd1 vccd1 vccd1 _17307_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14518_ _14549_/A vssd1 vssd1 vccd1 vccd1 _14518_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18286_ _18286_/A _18286_/B vssd1 vssd1 vccd1 vccd1 _18288_/C sky130_fd_sc_hd__xnor2_1
XFILLER_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15498_ _15498_/A _15497_/Y vssd1 vssd1 vccd1 vccd1 _15499_/B sky130_fd_sc_hd__or2b_1
XFILLER_30_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17237_ _17068_/X _17069_/X _17077_/B _17070_/X vssd1 vssd1 vccd1 vccd1 _17238_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_14449_ _15118_/A vssd1 vssd1 vccd1 vccd1 _14472_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16462__A _19512_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17168_ _16934_/X _16936_/Y _17166_/A vssd1 vssd1 vccd1 vccd1 _17170_/C sky130_fd_sc_hd__o21a_1
XFILLER_66_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16119_ _16119_/A _16153_/A vssd1 vssd1 vccd1 vccd1 _16119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17099_ _17098_/Y _17096_/X _11935_/X _15655_/X vssd1 vssd1 vccd1 vccd1 _17099_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_116_879 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20241__A1 _20290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19809_ _17610_/A _18455_/A _18461_/C _17613_/A _19668_/A vssd1 vssd1 vccd1 vccd1
+ _19809_/X sky130_fd_sc_hd__o32a_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18985__A2 _18490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13326__A _13663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22820_ _22820_/A _22820_/B vssd1 vssd1 vccd1 vccd1 _22820_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23191__A0 _15662_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14471__A2 _15233_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22751_ _22718_/X _22722_/C _22722_/A vssd1 vssd1 vccd1 vccd1 _22751_/X sky130_fd_sc_hd__a21o_1
XFILLER_198_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21702_ _21717_/A _21717_/B _21723_/A vssd1 vssd1 vccd1 vccd1 _21711_/A sky130_fd_sc_hd__o21a_1
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22682_ _22680_/X _22679_/Y _22633_/Y _22605_/A vssd1 vssd1 vccd1 vccd1 _22683_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_25_579 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21633_ _21633_/A vssd1 vssd1 vccd1 vccd1 _21668_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__18852__A _18959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_916 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16075__C _16075_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13982__A1 _13960_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21564_ _21564_/A _21564_/B _21564_/C vssd1 vssd1 vccd1 vccd1 _21565_/B sky130_fd_sc_hd__and3_1
XFILLER_138_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23303_ _23398_/CLK _23303_/D vssd1 vssd1 vccd1 vccd1 _23303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23246__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20515_ _20515_/A _20515_/B _20515_/C vssd1 vssd1 vccd1 vccd1 _20516_/A sky130_fd_sc_hd__nand3_1
X_21495_ _21495_/A _21495_/B _21495_/C vssd1 vssd1 vccd1 vccd1 _21559_/B sky130_fd_sc_hd__and3_1
XANTENNA__16372__A _16372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16920__A1 _14631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_971 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13734__A1 _13415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23234_ _23234_/A vssd1 vssd1 vccd1 vccd1 _23435_/D sky130_fd_sc_hd__clkbuf_1
X_20446_ _20446_/A _20446_/B _20446_/C vssd1 vssd1 vccd1 vccd1 _20453_/B sky130_fd_sc_hd__and3_1
XFILLER_109_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12942__C1 _21121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23165_ _23405_/Q input22/X _23167_/S vssd1 vssd1 vccd1 vccd1 _23166_/A sky130_fd_sc_hd__mux2_1
X_20377_ _20376_/A _20376_/B _20401_/B vssd1 vssd1 vccd1 vccd1 _20378_/B sky130_fd_sc_hd__o21ai_1
XFILLER_192_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22116_ _23273_/Q _22112_/A _22115_/B vssd1 vssd1 vccd1 vccd1 _22451_/B sky130_fd_sc_hd__o21ai_1
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23096_ _23096_/A vssd1 vssd1 vccd1 vccd1 _23374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17228__A2 _11972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22047_ _14614_/X _22047_/B _22186_/C vssd1 vssd1 vccd1 vccd1 _22049_/A sky130_fd_sc_hd__nand3b_1
XFILLER_47_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16436__B1 _15749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1075 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13820_ _13799_/X _13813_/X _13819_/Y vssd1 vssd1 vccd1 vccd1 _13820_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__13236__A _23477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13751_ _13738_/X _13750_/X _13747_/X _13748_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_18_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22949_ _23309_/Q input22/X _22951_/S vssd1 vssd1 vccd1 vccd1 _22950_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ _23447_/Q vssd1 vssd1 vccd1 vccd1 _13151_/B sky130_fd_sc_hd__clkinv_2
XFILLER_188_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16470_ _16394_/A _16517_/C _16415_/B vssd1 vssd1 vccd1 vccd1 _16483_/A sky130_fd_sc_hd__a21o_1
XANTENNA__21172__B _21453_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13682_ _13682_/A _13682_/B _13682_/C vssd1 vssd1 vccd1 vccd1 _13692_/B sky130_fd_sc_hd__nand3_1
XFILLER_71_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15421_ _15420_/C _14990_/A _14990_/B _15420_/D _15420_/A vssd1 vssd1 vccd1 vccd1
+ _15421_/X sky130_fd_sc_hd__a32o_1
XFILLER_54_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12633_ _12633_/A vssd1 vssd1 vccd1 vccd1 _12709_/A sky130_fd_sc_hd__buf_2
XANTENNA__19858__A _19858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14067__A _14777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18140_ _18252_/A _18140_/B _18140_/C vssd1 vssd1 vccd1 vccd1 _18141_/C sky130_fd_sc_hd__nand3b_1
X_15352_ _15348_/Y _15324_/A _15508_/A _15109_/X _15110_/X vssd1 vssd1 vccd1 vccd1
+ _15352_/Y sky130_fd_sc_hd__o2111ai_2
XFILLER_54_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12564_ _19090_/A _19089_/B _12563_/Y vssd1 vssd1 vccd1 vccd1 _12564_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_180_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18361__B1 _23535_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18481__B _18481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303_ _14303_/A _14310_/D vssd1 vssd1 vccd1 vccd1 _14304_/B sky130_fd_sc_hd__nand2_1
X_18071_ _18069_/Y _18070_/Y _18049_/B _18053_/A vssd1 vssd1 vccd1 vccd1 _18072_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_156_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23237__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15283_ _15221_/Y _15222_/Y _15392_/A _15392_/B _15282_/Y vssd1 vssd1 vccd1 vccd1
+ _15283_/X sky130_fd_sc_hd__o221a_1
X_12495_ _12536_/B vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13121__D _20905_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17022_ _17022_/A vssd1 vssd1 vccd1 vccd1 _17943_/A sky130_fd_sc_hd__buf_2
XFILLER_172_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14234_ _14236_/B _14235_/A _14235_/B vssd1 vssd1 vccd1 vccd1 _14306_/B sky130_fd_sc_hd__nand3b_1
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14165_ _14161_/Y _14162_/X _14164_/Y vssd1 vssd1 vccd1 vccd1 _14818_/B sky130_fd_sc_hd__o21ai_1
X_13116_ _13156_/A _21177_/B _13116_/C _13157_/B vssd1 vssd1 vccd1 vccd1 _13116_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_124_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14096_ _14096_/A vssd1 vssd1 vccd1 vccd1 _14097_/A sky130_fd_sc_hd__clkbuf_2
X_18973_ _18973_/A _18973_/B _18973_/C vssd1 vssd1 vccd1 vccd1 _18984_/B sky130_fd_sc_hd__nand3_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _17924_/A _17924_/B _17924_/C vssd1 vssd1 vccd1 vccd1 _17924_/X sky130_fd_sc_hd__or3_4
XFILLER_152_1120 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13047_ _13035_/X _13036_/X _20556_/C _20556_/A vssd1 vssd1 vccd1 vccd1 _13048_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_26_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18002__A _18002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17855_ _17855_/A vssd1 vssd1 vccd1 vccd1 _17988_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20774__A2 _20773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16806_ _17041_/B _16812_/B _16165_/A _15964_/B _16805_/X vssd1 vssd1 vccd1 vccd1
+ _17073_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_93_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17786_ _17776_/Y _17780_/Y _17782_/Y _17785_/Y vssd1 vssd1 vccd1 vccd1 _17786_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_54_619 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14998_ _15094_/B vssd1 vssd1 vccd1 vccd1 _15096_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19525_ _19525_/A _19525_/B _19525_/C _19525_/D vssd1 vssd1 vccd1 vccd1 _19578_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16737_ _16737_/A vssd1 vssd1 vccd1 vccd1 _16737_/Y sky130_fd_sc_hd__inv_2
X_13949_ _13949_/A vssd1 vssd1 vccd1 vccd1 _14029_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19456_ _19456_/A _19456_/B vssd1 vssd1 vccd1 vccd1 _19456_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16668_ _23427_/Q _16668_/B _16668_/C vssd1 vssd1 vccd1 vccd1 _16669_/B sky130_fd_sc_hd__nand3b_2
XFILLER_35_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18407_ _18407_/A _18407_/B _18407_/C _18407_/D vssd1 vssd1 vccd1 vccd1 _18408_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_50_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15619_ _23429_/Q vssd1 vssd1 vccd1 vccd1 _15665_/B sky130_fd_sc_hd__clkbuf_4
X_19387_ _19387_/A _19387_/B vssd1 vssd1 vccd1 vccd1 _19389_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13413__B1 _22264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18672__A _18868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16599_ _16153_/A _16152_/A _16588_/X vssd1 vssd1 vccd1 vccd1 _16599_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18338_ _18338_/A _18338_/B vssd1 vssd1 vccd1 vccd1 _18339_/C sky130_fd_sc_hd__xnor2_1
XFILLER_33_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11975__B1 _11902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16904__B _16908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23228__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18269_ _18269_/A _18231_/B vssd1 vssd1 vccd1 vccd1 _18288_/B sky130_fd_sc_hd__or2b_1
XFILLER_148_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16363__C1 _16499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16902__A1 _12004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20300_ _20341_/A _20300_/B vssd1 vssd1 vccd1 vccd1 _20303_/A sky130_fd_sc_hd__nand2_1
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12519__A2 _12509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21280_ _21278_/A _21453_/D _21279_/Y vssd1 vssd1 vccd1 vccd1 _21280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_144_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20231_ _20283_/A _20231_/B _20231_/C vssd1 vssd1 vccd1 vccd1 _20231_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_196_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16666__B1 _14631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20162_ _20167_/A _20167_/B _20232_/A vssd1 vssd1 vccd1 vccd1 _20162_/X sky130_fd_sc_hd__and3_1
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1086 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20093_ _19996_/A _19996_/B _19996_/C _19963_/B vssd1 vssd1 vccd1 vccd1 _20096_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_162_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12152__B1 _12093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20214__A1 _20217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14692__A2 _14672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_800 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19368__C1 _19900_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22803_ _22764_/C _22764_/A _22764_/B _22829_/B vssd1 vssd1 vccd1 vccd1 _22803_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20995_ _20995_/A _20995_/B _20995_/C vssd1 vssd1 vccd1 vccd1 _21131_/B sky130_fd_sc_hd__nand3_1
XANTENNA__22088__B _22089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12110__D _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22734_ _22734_/A vssd1 vssd1 vccd1 vccd1 _22810_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17394__B2 _17307_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16051__D1 _16046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22665_ _22582_/X _22580_/Y _22586_/Y _22664_/X vssd1 vssd1 vccd1 vccd1 _22670_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_41_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21616_ _21616_/A vssd1 vssd1 vccd1 vccd1 _21616_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17146__A1 _11882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22596_ _22499_/A _22499_/B _22499_/C _22595_/Y vssd1 vssd1 vccd1 vccd1 _22596_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21547_ _21371_/C _21548_/D _21371_/B _21637_/C _21502_/D vssd1 vssd1 vccd1 vccd1
+ _21547_/X sky130_fd_sc_hd__a32o_1
XANTENNA__14615__A _23297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13707__A1 _21778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12280_ _11611_/A _11611_/B _11717_/B _11717_/C _12279_/X vssd1 vssd1 vccd1 vccd1
+ _12280_/Y sky130_fd_sc_hd__a221oi_1
X_21478_ _21426_/X _21425_/Y _21474_/Y _21477_/Y vssd1 vssd1 vccd1 vccd1 _21482_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_112_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20055__C _20055_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23217_ _23428_/Q input12/X _23217_/S vssd1 vssd1 vccd1 vccd1 _23218_/A sky130_fd_sc_hd__mux2_1
X_20429_ _20426_/X _20427_/X _20429_/S vssd1 vssd1 vccd1 vccd1 _20430_/B sky130_fd_sc_hd__mux2_2
XFILLER_181_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23148_ _18434_/A input13/X _23156_/S vssd1 vssd1 vccd1 vccd1 _23149_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__22270__C _22270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_988 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15970_ _17590_/A _17592_/A _15860_/C _18756_/A vssd1 vssd1 vccd1 vccd1 _16598_/A
+ sky130_fd_sc_hd__o211ai_4
X_23079_ _23079_/A vssd1 vssd1 vccd1 vccd1 _23366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18949__A2 _18096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input32_A wb_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13340__C1 _13304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17606__C1 _20142_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14921_ _14923_/A vssd1 vssd1 vccd1 vccd1 _14926_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17640_ _17410_/Y _17625_/Y _19957_/D _17898_/D _17629_/Y vssd1 vssd1 vccd1 vccd1
+ _17641_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_29_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14852_ _23270_/D _14849_/Y vssd1 vssd1 vccd1 vccd1 _14962_/A sky130_fd_sc_hd__or2b_1
XFILLER_29_660 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13803_ _13803_/A _13803_/B vssd1 vssd1 vccd1 vccd1 _21927_/A sky130_fd_sc_hd__nand2_1
X_17571_ _17571_/A _17737_/A vssd1 vssd1 vccd1 vccd1 _17571_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__12446__A1 _12246_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14783_ _14788_/A _14783_/B _14788_/C vssd1 vssd1 vccd1 vccd1 _14783_/X sky130_fd_sc_hd__and3_1
XANTENNA__21166__C1 _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11995_ _12426_/B vssd1 vssd1 vccd1 vccd1 _19019_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_44_630 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20508__A2 _20504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19310_ _19304_/X _19307_/Y _19309_/Y vssd1 vssd1 vccd1 vccd1 _19310_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16522_ _16522_/A _16522_/B vssd1 vssd1 vccd1 vccd1 _16522_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13734_ _13415_/X _13701_/Y _13659_/Y _13732_/X _13707_/X vssd1 vssd1 vccd1 vccd1
+ _13739_/B sky130_fd_sc_hd__o311a_1
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19241_ _19135_/Y _19410_/C _19142_/Y vssd1 vssd1 vccd1 vccd1 _19241_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16453_ _16370_/X _16384_/X _16356_/A _16225_/X _16457_/A vssd1 vssd1 vccd1 vccd1
+ _16453_/X sky130_fd_sc_hd__o221a_1
XFILLER_32_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13665_ _13665_/A _13666_/A _13666_/B vssd1 vssd1 vccd1 vccd1 _13680_/C sky130_fd_sc_hd__nand3_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19126__A2 _12185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15404_/A _15435_/B vssd1 vssd1 vccd1 vccd1 _15433_/B sky130_fd_sc_hd__nor2_1
X_12616_ _13121_/A _13121_/B _21039_/B vssd1 vssd1 vccd1 vccd1 _12945_/B sky130_fd_sc_hd__and3_1
X_19172_ _19172_/A _19172_/B _19172_/C vssd1 vssd1 vccd1 vccd1 _19183_/B sky130_fd_sc_hd__nand3_2
XFILLER_157_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16384_ _16384_/A vssd1 vssd1 vccd1 vccd1 _16384_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13540_/A _13540_/B _13540_/C _13535_/A vssd1 vssd1 vccd1 vccd1 _13596_/Y
+ sky130_fd_sc_hd__a31oi_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18334__B1 _20320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11957__B1 _11915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12029__B _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18123_ _18123_/A _18123_/B _18123_/C vssd1 vssd1 vccd1 vccd1 _18133_/A sky130_fd_sc_hd__and3_1
XFILLER_12_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15335_ _15395_/B _15335_/B vssd1 vssd1 vccd1 vccd1 _15337_/A sky130_fd_sc_hd__nand2_2
XFILLER_157_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12547_ _12547_/A _12547_/B vssd1 vssd1 vccd1 vccd1 _12547_/X sky130_fd_sc_hd__and2_1
XFILLER_145_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16896__B1 _11830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18054_ _17943_/A _18139_/C _18138_/A _18138_/B vssd1 vssd1 vccd1 vccd1 _18054_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15266_ _15363_/D vssd1 vssd1 vccd1 vccd1 _15420_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_172_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12478_ _12478_/A _12478_/B _12478_/C vssd1 vssd1 vccd1 vccd1 _18524_/B sky130_fd_sc_hd__nand3_4
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17005_ _23519_/Q _16776_/A _23520_/Q vssd1 vssd1 vccd1 vccd1 _17014_/B sky130_fd_sc_hd__o21ai_1
X_14217_ _14222_/A _14222_/B _14217_/C vssd1 vssd1 vccd1 vccd1 _14218_/C sky130_fd_sc_hd__nand3_1
X_15197_ _14834_/A _14777_/C _14777_/A _15093_/B _15093_/A vssd1 vssd1 vccd1 vccd1
+ _15197_/X sky130_fd_sc_hd__a32o_1
XFILLER_99_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14910__A3 _14777_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21358__A _21358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148_ _14148_/A _14148_/B _14148_/C vssd1 vssd1 vccd1 vccd1 _14156_/B sky130_fd_sc_hd__nand3_2
XFILLER_113_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15356__A _15356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18956_ _18954_/Y _18955_/Y _18950_/Y _19410_/A vssd1 vssd1 vccd1 vccd1 _18956_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14079_ _14078_/Y _14865_/A _14188_/A vssd1 vssd1 vccd1 vccd1 _14752_/A sky130_fd_sc_hd__a21o_1
XFILLER_140_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17907_ _17901_/A _17901_/B _17902_/A vssd1 vssd1 vccd1 vccd1 _17909_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__15075__B _15075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18887_ _18751_/X _18752_/X _18878_/Y _18886_/Y vssd1 vssd1 vccd1 vccd1 _18897_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_117_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21944__A1 _21892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23534__CLK _23538_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17838_ _17838_/A _17838_/B _17838_/C vssd1 vssd1 vccd1 vccd1 _17911_/A sky130_fd_sc_hd__and3_1
XFILLER_55_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12211__C _12211_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17769_ _17580_/A _17580_/B _17583_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17769_/Y
+ sky130_fd_sc_hd__a22oi_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18168__A3 _17753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19508_ _19503_/X _19307_/Y _19507_/Y vssd1 vssd1 vccd1 vccd1 _19525_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__19365__A2 _15861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20780_ _20625_/B _20778_/X _20779_/X vssd1 vssd1 vccd1 vccd1 _20789_/A sky130_fd_sc_hd__o21ai_1
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19439_ _19434_/X _19435_/Y _19436_/X _19438_/Y vssd1 vssd1 vccd1 vccd1 _19439_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15926__A2 _17409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22450_ _22450_/A _22450_/B vssd1 vssd1 vccd1 vccd1 _22454_/A sky130_fd_sc_hd__nand2_2
XFILLER_10_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16634__B _18755_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21401_ _21476_/A _21476_/B vssd1 vssd1 vccd1 vccd1 _21407_/A sky130_fd_sc_hd__xnor2_2
XFILLER_109_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22381_ _22381_/A _22381_/B _22381_/C vssd1 vssd1 vccd1 vccd1 _22384_/A sky130_fd_sc_hd__nand3_1
XFILLER_124_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21332_ _21331_/B _21331_/C _21266_/X vssd1 vssd1 vccd1 vccd1 _21333_/D sky130_fd_sc_hd__a21bo_1
XFILLER_136_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13165__A2 _12979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21263_ _21263_/A vssd1 vssd1 vccd1 vccd1 _23545_/D sky130_fd_sc_hd__clkbuf_1
X_23002_ _23002_/A vssd1 vssd1 vccd1 vccd1 _23332_/D sky130_fd_sc_hd__clkbuf_1
X_20214_ _20217_/D _19862_/B _19862_/C _18077_/A _20142_/B vssd1 vssd1 vccd1 vccd1
+ _20271_/D sky130_fd_sc_hd__a32o_1
XFILLER_144_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21268__A _21268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12912__A2 _12902_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21194_ _21194_/A _21194_/B vssd1 vssd1 vccd1 vccd1 _21194_/Y sky130_fd_sc_hd__nand2_2
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20145_ _20141_/X _20143_/Y _20148_/C vssd1 vssd1 vccd1 vccd1 _20158_/A sky130_fd_sc_hd__o21bai_4
XFILLER_131_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13468__A3 _21892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ _19975_/A _19975_/B _20073_/A _20073_/B vssd1 vssd1 vccd1 vccd1 _20076_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23137__A0 _18997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_714 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_bq_clk_i clkbuf_2_3_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_bq_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13625__B1 _22484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19356__A2 _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16528__C _16536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _18972_/A vssd1 vssd1 vccd1 vccd1 _15718_/A sky130_fd_sc_hd__clkbuf_2
X_20978_ _20978_/A _20978_/B vssd1 vssd1 vccd1 vccd1 _20979_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_808 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22717_ _22717_/A _22717_/B _22717_/C _22789_/B vssd1 vssd1 vccd1 vccd1 _22722_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_14_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11651__A2 _11721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15917__A2 _11740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13450_ _13701_/A _21921_/C _13701_/C vssd1 vssd1 vccd1 vccd1 _13450_/Y sky130_fd_sc_hd__nand3_1
X_22648_ _22703_/A _22830_/D _22701_/C _22641_/B _22638_/Y vssd1 vssd1 vccd1 vccd1
+ _22649_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_139_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12401_ _16027_/B vssd1 vssd1 vccd1 vccd1 _19011_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13381_ _13423_/A vssd1 vssd1 vccd1 vccd1 _21883_/A sky130_fd_sc_hd__buf_2
X_22579_ _22577_/Y _22578_/X _22564_/X vssd1 vssd1 vccd1 vccd1 _22579_/Y sky130_fd_sc_hd__o21bai_2
XANTENNA__20066__B _20066_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15120_ _15120_/A _15120_/B _15263_/A _15120_/D vssd1 vssd1 vccd1 vccd1 _15121_/A
+ sky130_fd_sc_hd__nand4_1
X_12332_ _12273_/B _12273_/C _12273_/D _12273_/A vssd1 vssd1 vccd1 vccd1 _12339_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15051_ _15050_/A _15050_/B _15050_/C vssd1 vssd1 vccd1 vccd1 _15052_/C sky130_fd_sc_hd__a21o_1
X_12263_ _12265_/C _12265_/B _12214_/X _11898_/X vssd1 vssd1 vccd1 vccd1 _12273_/D
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_108_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14002_ _14002_/A _14162_/B _14433_/D _14003_/A vssd1 vssd1 vccd1 vccd1 _14253_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12194_ _11952_/Y _11966_/B _11937_/X vssd1 vssd1 vccd1 vccd1 _12196_/C sky130_fd_sc_hd__a21oi_1
XFILLER_150_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput62 _14666_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[17] sky130_fd_sc_hd__buf_2
X_18810_ _18810_/A _23393_/Q vssd1 vssd1 vccd1 vccd1 _18811_/C sky130_fd_sc_hd__nor2_1
XFILLER_123_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput73 _14708_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[27] sky130_fd_sc_hd__buf_2
X_19790_ _19635_/A _19788_/A _19923_/A _19788_/C _19636_/B vssd1 vssd1 vccd1 vccd1
+ _19791_/B sky130_fd_sc_hd__a221o_1
XFILLER_110_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput84 _14597_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[8] sky130_fd_sc_hd__buf_2
Xoutput95 _23269_/Q vssd1 vssd1 vccd1 vccd1 y[7] sky130_fd_sc_hd__buf_2
XFILLER_49_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18741_ _12564_/Y _18749_/A _12565_/X _18733_/C _18733_/B vssd1 vssd1 vccd1 vccd1
+ _18741_/Y sky130_fd_sc_hd__o311ai_4
XANTENNA__21906__A _21906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15953_ _17964_/C _17964_/A _15957_/C _23260_/B vssd1 vssd1 vccd1 vccd1 _19364_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_49_744 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17391__A _19653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14904_ _14904_/A vssd1 vssd1 vccd1 vccd1 _15366_/A sky130_fd_sc_hd__clkbuf_2
X_18672_ _18868_/A _18868_/B _18868_/C vssd1 vssd1 vccd1 vccd1 _18672_/Y sky130_fd_sc_hd__nand3_1
X_15884_ _15884_/A vssd1 vssd1 vccd1 vccd1 _15884_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23128__A0 _11665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17623_ _17656_/A _17656_/B vssd1 vssd1 vccd1 vccd1 _17657_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_438 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14835_ _14835_/A _15298_/B _14835_/C vssd1 vssd1 vccd1 vccd1 _14835_/X sky130_fd_sc_hd__and3_1
XFILLER_5_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _17485_/A _17430_/A _17553_/Y vssd1 vssd1 vccd1 vccd1 _17555_/A sky130_fd_sc_hd__a21oi_1
X_14766_ _14766_/A _14766_/B _14766_/C vssd1 vssd1 vccd1 vccd1 _14783_/B sky130_fd_sc_hd__nand3_1
XFILLER_32_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11978_ _23389_/Q vssd1 vssd1 vccd1 vccd1 _18469_/D sky130_fd_sc_hd__inv_2
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16505_ _12238_/X _16398_/X _16526_/C _19653_/A _16399_/X vssd1 vssd1 vccd1 vccd1
+ _16505_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_44_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13717_ _13748_/C _13715_/X _13716_/Y vssd1 vssd1 vccd1 vccd1 _13717_/Y sky130_fd_sc_hd__a21oi_1
X_17485_ _17485_/A _17485_/B _17485_/C vssd1 vssd1 vccd1 vccd1 _17654_/B sky130_fd_sc_hd__and3_1
XFILLER_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14697_ _23406_/Q _14693_/X _14677_/X _23438_/Q _14696_/X vssd1 vssd1 vccd1 vccd1
+ _14697_/X sky130_fd_sc_hd__a221o_1
XFILLER_149_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19224_ _19217_/X _19222_/X _19230_/A vssd1 vssd1 vccd1 vccd1 _19224_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_176_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16436_ _11882_/X _11883_/X _15749_/A _15749_/B vssd1 vssd1 vccd1 vccd1 _16436_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13648_ _13414_/A _13414_/B _13414_/C _13474_/A _13474_/B vssd1 vssd1 vccd1 vccd1
+ _13648_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_60_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19155_ _18799_/B _19155_/B _19155_/C _19155_/D vssd1 vssd1 vccd1 vccd1 _19156_/A
+ sky130_fd_sc_hd__nand4b_2
X_16367_ _12146_/X _12147_/X _15860_/C _15964_/B _12149_/X vssd1 vssd1 vccd1 vccd1
+ _16398_/A sky130_fd_sc_hd__o2111ai_1
X_13579_ _13709_/C vssd1 vssd1 vccd1 vccd1 _13736_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18106_ _18106_/A _18179_/B _18106_/C vssd1 vssd1 vccd1 vccd1 _18108_/A sky130_fd_sc_hd__nand3_1
XFILLER_173_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15318_ _15233_/C _15419_/C _15419_/D _15238_/Y vssd1 vssd1 vccd1 vccd1 _15321_/A
+ sky130_fd_sc_hd__a31o_1
X_19086_ _12167_/X _12168_/X _17249_/X _17250_/X _20317_/B vssd1 vssd1 vccd1 vccd1
+ _19263_/A sky130_fd_sc_hd__o221a_2
XFILLER_145_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16298_ _12146_/X _12147_/X _15862_/A _15862_/B _12149_/A vssd1 vssd1 vccd1 vccd1
+ _16366_/A sky130_fd_sc_hd__o221ai_2
XFILLER_172_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18037_ _18036_/B _18037_/B _18037_/C vssd1 vssd1 vccd1 vccd1 _18123_/A sky130_fd_sc_hd__nand3b_2
XFILLER_172_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15249_ _15249_/A _15249_/B vssd1 vssd1 vccd1 vccd1 _15250_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18086__A2 _12506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16097__A1 _16020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19988_ _19985_/A _19985_/B _19986_/A vssd1 vssd1 vccd1 vccd1 _19991_/A sky130_fd_sc_hd__o21ai_1
XFILLER_154_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20142__D _20142_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18939_ _18755_/Y _18934_/Y _19381_/D _18938_/X _18080_/A vssd1 vssd1 vccd1 vccd1
+ _19141_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_39_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21917__A1 _22487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21950_ _21875_/Y _21782_/C _21806_/X _21948_/Y _21949_/Y vssd1 vssd1 vccd1 vccd1
+ _21982_/B sky130_fd_sc_hd__o2111ai_4
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11866__C1 _19363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23119__A0 _11677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20901_ _21046_/A _21046_/B _20901_/C _23300_/Q vssd1 vssd1 vccd1 vccd1 _20903_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21881_ _22521_/A _22363_/A _22521_/C vssd1 vssd1 vccd1 vccd1 _21881_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__11881__A2 _16462_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20832_ _21121_/B _20887_/A _20887_/B vssd1 vssd1 vccd1 vccd1 _20841_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__22647__A _22647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23551_ _23558_/CLK _23551_/D vssd1 vssd1 vccd1 vccd1 _23551_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18010__A2 _18276_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20763_ _20763_/A _21030_/A vssd1 vssd1 vccd1 vccd1 _20766_/A sky130_fd_sc_hd__nand2_1
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19659__C _19659_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22502_ _22541_/A _22541_/B _22541_/C _22541_/D vssd1 vssd1 vccd1 vccd1 _22513_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_74_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23482_ _23510_/CLK hold19/X vssd1 vssd1 vccd1 vccd1 _23482_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14032__B1 _14031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20694_ _20666_/A _20666_/B _20667_/A vssd1 vssd1 vccd1 vccd1 _20695_/C sky130_fd_sc_hd__o21ai_1
XFILLER_167_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16364__B _16364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12892__B _21124_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14583__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22433_ _22457_/A _22524_/A _22457_/B vssd1 vssd1 vccd1 vccd1 _22435_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__20105__B1 _20106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14583__B2 _14031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19510__A2 _19868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22364_ _22487_/A _22364_/B _22637_/C _22636_/C vssd1 vssd1 vccd1 vccd1 _22496_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_175_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19675__B _19868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21315_ _21502_/D _21387_/B _21194_/Y _21312_/X vssd1 vssd1 vccd1 vccd1 _21315_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_124_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_760 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22295_ _22508_/A _22508_/B _22569_/B vssd1 vssd1 vccd1 vccd1 _22297_/A sky130_fd_sc_hd__nand3_1
XFILLER_105_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21246_ _21255_/A vssd1 vssd1 vccd1 vccd1 _21246_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__20959__A2 _12850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21177_ _21370_/A _21177_/B _21369_/A vssd1 vssd1 vccd1 vccd1 _21178_/C sky130_fd_sc_hd__nand3_1
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_98 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14331__C _14331_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20128_ _20128_/A _20128_/B vssd1 vssd1 vccd1 vccd1 _23530_/D sky130_fd_sc_hd__nand2_1
XFILLER_131_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22030__B1 _13486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12950_ _13177_/B _13177_/C _12674_/X vssd1 vssd1 vccd1 vccd1 _12950_/X sky130_fd_sc_hd__a21o_1
X_20059_ _20210_/C _18211_/B _20045_/Y _20048_/Y _20050_/Y vssd1 vssd1 vccd1 vccd1
+ _20060_/C sky130_fd_sc_hd__o221ai_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11901_ _12016_/A _12016_/B _12032_/A _19548_/A _16497_/A vssd1 vssd1 vccd1 vccd1
+ _11902_/C sky130_fd_sc_hd__o2111ai_4
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _12880_/Y _20528_/B vssd1 vssd1 vccd1 vccd1 _20669_/A sky130_fd_sc_hd__and2b_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19329__A2 _19482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14620_ _23426_/Q vssd1 vssd1 vccd1 vccd1 _16191_/A sky130_fd_sc_hd__clkbuf_4
X_11832_ _11672_/Y _11754_/A _11746_/B _11743_/A vssd1 vssd1 vccd1 vccd1 _11834_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18537__B1 _17593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14551_ _14551_/A vssd1 vssd1 vccd1 vccd1 _14551_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11820_/A vssd1 vssd1 vccd1 vccd1 _11766_/A sky130_fd_sc_hd__buf_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13502_ _22280_/B _13701_/C _13701_/A _13709_/C _22381_/C vssd1 vssd1 vccd1 vccd1
+ _13502_/X sky130_fd_sc_hd__a32o_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _17248_/Y _17252_/Y _17269_/X vssd1 vssd1 vccd1 vccd1 _17270_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14482_ _14410_/Y _14405_/Y _14380_/Y vssd1 vssd1 vccd1 vccd1 _14486_/A sky130_fd_sc_hd__a21bo_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11739_/B vssd1 vssd1 vccd1 vccd1 _11694_/X sky130_fd_sc_hd__buf_2
XFILLER_174_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13433_ _13433_/A _13433_/B vssd1 vssd1 vccd1 vccd1 _13434_/A sky130_fd_sc_hd__nand2_1
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11699__A _11830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16221_ _16183_/X _16193_/Y _16199_/Y vssd1 vssd1 vccd1 vccd1 _16233_/A sky130_fd_sc_hd__o21ai_1
XFILLER_174_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16705__D _16706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16152_ _16152_/A vssd1 vssd1 vccd1 vccd1 _16153_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13364_ _13364_/A vssd1 vssd1 vccd1 vccd1 _13433_/A sky130_fd_sc_hd__buf_2
XFILLER_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12315_ _12353_/A _12379_/A _12314_/Y vssd1 vssd1 vccd1 vccd1 _12360_/B sky130_fd_sc_hd__o21ai_2
X_15103_ _15000_/B _15096_/Y _15175_/C _15099_/Y _15446_/B vssd1 vssd1 vccd1 vccd1
+ _15107_/C sky130_fd_sc_hd__o2111ai_4
X_16083_ _15837_/Y _15810_/X _16062_/B _16022_/A _15895_/C vssd1 vssd1 vccd1 vccd1
+ _16084_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_182_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13295_ _23478_/Q vssd1 vssd1 vccd1 vccd1 _21882_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__16290__A _17243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23538__D _23538_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19911_ _19911_/A vssd1 vssd1 vccd1 vccd1 _19911_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _15035_/A _15035_/B _15030_/X _15031_/Y vssd1 vssd1 vccd1 vccd1 _15036_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__19265__A1 _19082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12246_ _11861_/A _19156_/C _12245_/X vssd1 vssd1 vccd1 vccd1 _12246_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_177_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19265__B2 _20368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16079__A1 _15878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19842_ _19505_/X _19504_/X _19494_/D _20369_/B vssd1 vssd1 vccd1 vccd1 _19848_/B
+ sky130_fd_sc_hd__o211ai_1
X_12177_ _12177_/A _12177_/B vssd1 vssd1 vccd1 vccd1 _12177_/Y sky130_fd_sc_hd__nand2_2
XFILLER_69_828 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12323__A _12323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output63_A _14671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15826__B2 _12018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19773_ _19613_/Y _19638_/Y _19768_/A _19625_/A _19439_/Y vssd1 vssd1 vccd1 vccd1
+ _19773_/X sky130_fd_sc_hd__o2111a_1
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16985_ _17025_/A _16984_/Y _17369_/A vssd1 vssd1 vccd1 vccd1 _16994_/D sky130_fd_sc_hd__o21ai_4
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18724_ _18722_/Y _18723_/Y _18914_/B _18914_/A vssd1 vssd1 vccd1 vccd1 _18725_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_114_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15936_ _15936_/A vssd1 vssd1 vccd1 vccd1 _17625_/B sky130_fd_sc_hd__buf_2
XANTENNA__17579__A1 _16479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18655_ _18972_/C vssd1 vssd1 vccd1 vccd1 _20047_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15353__B _15353_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _15879_/A _15879_/B _15867_/C vssd1 vssd1 vccd1 vccd1 _15867_/Y sky130_fd_sc_hd__nand3_2
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18945__A _19381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17606_ _14599_/X _16203_/Y _15791_/X _17753_/B _20142_/D vssd1 vssd1 vccd1 vccd1
+ _17606_/X sky130_fd_sc_hd__o311a_4
X_14818_ _14818_/A _14818_/B _14821_/A vssd1 vssd1 vccd1 vccd1 _14821_/B sky130_fd_sc_hd__nand3_1
XFILLER_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18586_ _18586_/A _18586_/B _18586_/C vssd1 vssd1 vccd1 vccd1 _18733_/B sky130_fd_sc_hd__nand3_2
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18528__B1 _18499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15798_ _15798_/A vssd1 vssd1 vccd1 vccd1 _17414_/C sky130_fd_sc_hd__buf_4
XFILLER_178_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17537_ _17537_/A _17537_/B vssd1 vssd1 vccd1 vccd1 _17934_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14749_ _15439_/C vssd1 vssd1 vccd1 vccd1 _14749_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17468_ _17454_/Y _17467_/X _17457_/Y _17960_/A _18172_/D vssd1 vssd1 vccd1 vccd1
+ _17562_/B sky130_fd_sc_hd__o2111ai_1
XANTENNA__15800__C _17414_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19207_ _18435_/A _11841_/Y _11948_/X _11951_/X _11849_/A vssd1 vssd1 vccd1 vccd1
+ _19207_/X sky130_fd_sc_hd__o221a_1
XFILLER_32_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16419_ _16475_/B _16475_/C _16474_/B vssd1 vssd1 vccd1 vccd1 _16472_/B sky130_fd_sc_hd__nand3_1
XANTENNA__14565__A1 _14188_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14565__B2 _11743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17399_ _17239_/X _17397_/Y _17395_/Y vssd1 vssd1 vccd1 vccd1 _17401_/A sky130_fd_sc_hd__a21oi_1
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19138_ _19138_/A _19138_/B vssd1 vssd1 vccd1 vccd1 _19139_/B sky130_fd_sc_hd__nand2_1
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19069_ _19069_/A _19069_/B _19069_/C vssd1 vssd1 vccd1 vccd1 _19069_/Y sky130_fd_sc_hd__nand3_4
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21100_ _21121_/A _21493_/C vssd1 vssd1 vccd1 vccd1 _21115_/A sky130_fd_sc_hd__nand2_1
XFILLER_191_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22080_ _21936_/B _21994_/Y _21995_/Y vssd1 vssd1 vccd1 vccd1 _22083_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__15528__B _15528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21063__A1 _12815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21031_ _21031_/A _21031_/B _21031_/C vssd1 vssd1 vccd1 vccd1 _21031_/Y sky130_fd_sc_hd__nand3_1
XFILLER_114_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13329__A _13660_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19008__A1 _19043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22982_ _13304_/X input34/X _22990_/S vssd1 vssd1 vccd1 vccd1 _22983_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22563__A1 _13547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21933_ _21747_/Y _21749_/Y _22045_/B _21910_/B _22043_/A vssd1 vssd1 vccd1 vccd1
+ _21933_/X sky130_fd_sc_hd__o311a_1
XFILLER_28_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18277__D _18277_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21864_ _21864_/A _23271_/Q _21864_/C vssd1 vssd1 vccd1 vccd1 _21864_/Y sky130_fd_sc_hd__nand3_2
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16793__A2 _16796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20815_ _12877_/Y _21278_/A _21054_/B _21065_/A _20973_/A vssd1 vssd1 vccd1 vccd1
+ _20819_/D sky130_fd_sc_hd__o2111ai_1
XFILLER_179_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21795_ _13495_/A _13620_/B _13620_/C _13465_/A _13431_/A vssd1 vssd1 vccd1 vccd1
+ _21795_/X sky130_fd_sc_hd__o32a_1
XANTENNA__19192__B1 _19210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22096__B _22096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23534_ _23538_/CLK _23534_/D vssd1 vssd1 vccd1 vccd1 _23534_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_196_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20746_ _21008_/C _20577_/Y _21008_/B vssd1 vssd1 vccd1 vccd1 _20748_/B sky130_fd_sc_hd__o21ai_1
XFILLER_196_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22079__B1 _21995_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14556__A1 _11604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23465_ _23559_/CLK _23477_/Q vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfxtp_1
XFILLER_137_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20677_ _20529_/B _20674_/Y _20676_/Y vssd1 vssd1 vccd1 vccd1 _20678_/B sky130_fd_sc_hd__o21ai_1
XFILLER_195_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22416_ _22414_/X _22415_/Y _22411_/X _22410_/Y _22541_/A vssd1 vssd1 vccd1 vccd1
+ _22417_/C sky130_fd_sc_hd__o2111ai_2
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19495__A1 _19951_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23396_ _23396_/CLK _23396_/D vssd1 vssd1 vccd1 vccd1 _23396_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12031__A2 _11846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22347_ _21981_/C _21968_/A _21970_/A _21981_/B vssd1 vssd1 vccd1 vccd1 _22348_/D
+ sky130_fd_sc_hd__a22oi_1
XFILLER_191_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16848__A3 _18607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16702__C1 _17388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11790__A1 _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ _12100_/A _12100_/B _12100_/C vssd1 vssd1 vccd1 vccd1 _18447_/B sky130_fd_sc_hd__nand3_4
XFILLER_163_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13080_ _12906_/Y _13076_/X _13077_/Y _13079_/Y vssd1 vssd1 vccd1 vccd1 _20595_/B
+ sky130_fd_sc_hd__o211ai_4
X_22278_ _22569_/A _22278_/B _22569_/C vssd1 vssd1 vccd1 vccd1 _22386_/A sky130_fd_sc_hd__nand3_4
XFILLER_3_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14342__B _14777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ _12051_/A _11846_/A _12022_/X _12025_/X _12011_/X vssd1 vssd1 vccd1 vccd1
+ _12159_/B sky130_fd_sc_hd__o221ai_2
XFILLER_88_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21229_ _21333_/A vssd1 vssd1 vccd1 vccd1 _21229_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16481__A1 _12379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16481__B2 _16480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16770_ _16576_/B _16339_/X _16575_/A vssd1 vssd1 vccd1 vccd1 _16771_/A sky130_fd_sc_hd__o21a_1
XFILLER_120_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13982_ _13960_/Y _13964_/Y _13969_/Y _13971_/X _14150_/D vssd1 vssd1 vccd1 vccd1
+ _13991_/A sky130_fd_sc_hd__o311ai_1
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ _15721_/A vssd1 vssd1 vccd1 vccd1 _15721_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _12571_/X _12796_/X _13177_/A _12766_/X vssd1 vssd1 vccd1 vccd1 _12933_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11845__A2 _11822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18440_ _18440_/A vssd1 vssd1 vccd1 vccd1 _18440_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _15652_/A vssd1 vssd1 vccd1 vccd1 _16866_/A sky130_fd_sc_hd__buf_2
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14244__B1 _14097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12864_ _12864_/A _12864_/B vssd1 vssd1 vccd1 vccd1 _21065_/A sky130_fd_sc_hd__nand2_2
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22306__B2 _22126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14603_ _12100_/B _14544_/X _14600_/X _14602_/X vssd1 vssd1 vccd1 vccd1 _14603_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _18371_/A _18371_/B vssd1 vssd1 vccd1 vccd1 _23595_/D sky130_fd_sc_hd__nor2_1
X_11815_ _11815_/A vssd1 vssd1 vccd1 vccd1 _11815_/X sky130_fd_sc_hd__buf_2
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15583_ _23511_/Q _23512_/Q _15585_/D _15574_/A vssd1 vssd1 vccd1 vccd1 _15584_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _13051_/C _13051_/A vssd1 vssd1 vccd1 vccd1 _12796_/A sky130_fd_sc_hd__nand2_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17327_/B _17322_/B _17322_/C vssd1 vssd1 vccd1 vccd1 _17330_/A sky130_fd_sc_hd__nand3b_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ _23184_/D vssd1 vssd1 vccd1 vccd1 _14534_/X sky130_fd_sc_hd__clkbuf_2
X_11746_ _11746_/A _11746_/B _11746_/C vssd1 vssd1 vccd1 vccd1 _11789_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12270__A2 _19675_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17253_ _17248_/Y _17252_/Y _16370_/X _17565_/A vssd1 vssd1 vccd1 vccd1 _17267_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_41_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14465_ _14465_/A _14465_/B _14465_/C _14465_/D vssd1 vssd1 vccd1 vccd1 _14465_/X
+ sky130_fd_sc_hd__and4_1
X_11677_ _11745_/A vssd1 vssd1 vccd1 vccd1 _11677_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16204_ _14599_/X _16203_/Y _15791_/X _16213_/A _19165_/C vssd1 vssd1 vccd1 vccd1
+ _16217_/B sky130_fd_sc_hd__o311a_1
X_13416_ _13416_/A vssd1 vssd1 vccd1 vccd1 _13486_/B sky130_fd_sc_hd__buf_2
XFILLER_128_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17184_ _17184_/A vssd1 vssd1 vccd1 vccd1 _17184_/Y sky130_fd_sc_hd__inv_2
X_14396_ _14396_/A _14396_/B _14396_/C _14760_/B vssd1 vssd1 vccd1 vccd1 _14436_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_128_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21293__A1 _21545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16135_ _16135_/A _16135_/B _16135_/C vssd1 vssd1 vccd1 vccd1 _16136_/A sky130_fd_sc_hd__nand3_1
X_13347_ _21744_/C _21902_/C _13394_/A vssd1 vssd1 vccd1 vccd1 _13620_/C sky130_fd_sc_hd__a21oi_4
XFILLER_6_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16451__C _16451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16066_ _16066_/A _16523_/C _16066_/C _19670_/A vssd1 vssd1 vccd1 vccd1 _16469_/A
+ sky130_fd_sc_hd__or4_4
X_13278_ _13741_/B _13741_/C _13469_/A vssd1 vssd1 vccd1 vccd1 _13516_/A sky130_fd_sc_hd__a21o_1
X_12229_ _12542_/A _18437_/D _12542_/B vssd1 vssd1 vccd1 vccd1 _12546_/B sky130_fd_sc_hd__nand3_1
X_15017_ _15155_/A _15225_/C _15253_/B _15017_/D vssd1 vssd1 vccd1 vccd1 _15081_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22793__A1 _22560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19825_ _20081_/B _19668_/X _19669_/X _19670_/X _19682_/B vssd1 vssd1 vccd1 vccd1
+ _19825_/X sky130_fd_sc_hd__o311a_1
XFILLER_64_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19756_ _19598_/Y _19755_/Y _19746_/Y vssd1 vssd1 vccd1 vccd1 _19757_/C sky130_fd_sc_hd__a21oi_1
X_16968_ _16704_/B _18277_/D _16749_/C _16662_/Y vssd1 vssd1 vccd1 vccd1 _16969_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_96_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18707_ _18707_/A _18707_/B vssd1 vssd1 vccd1 vccd1 _18708_/B sky130_fd_sc_hd__nor2_1
XANTENNA__23275__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18213__A2 _17323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15919_ _15937_/A vssd1 vssd1 vccd1 vccd1 _17137_/C sky130_fd_sc_hd__clkbuf_2
X_19687_ _19575_/A _19575_/B _19578_/A _19643_/Y vssd1 vssd1 vccd1 vccd1 _19796_/A
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__18675__A _18675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16899_ _11822_/A _15774_/A _16686_/A _11848_/X vssd1 vssd1 vccd1 vccd1 _16899_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18638_ _11896_/A _11896_/B _18476_/A _18484_/A _18479_/A vssd1 vssd1 vccd1 vccd1
+ _18639_/B sky130_fd_sc_hd__o221a_2
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18569_ _18569_/A vssd1 vssd1 vccd1 vccd1 _19090_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20600_ _20583_/Y _20585_/Y _21008_/A _20593_/C _20585_/A vssd1 vssd1 vccd1 vccd1
+ _20614_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_21_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21580_ _23570_/Q vssd1 vssd1 vccd1 vccd1 _21625_/A sky130_fd_sc_hd__inv_2
XANTENNA__16527__A2 _16536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12261__A2 _11898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20531_ _13053_/X _20676_/A _20670_/A vssd1 vssd1 vccd1 vccd1 _20533_/A sky130_fd_sc_hd__o21ai_1
XFILLER_162_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23250_ _23443_/Q input28/X _23250_/S vssd1 vssd1 vccd1 vccd1 _23251_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20462_ _20902_/B _23458_/Q vssd1 vssd1 vccd1 vccd1 _20613_/A sky130_fd_sc_hd__and2_1
XANTENNA__13050__C _13052_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22201_ _22177_/Y _22195_/Y _22200_/Y vssd1 vssd1 vccd1 vccd1 _22201_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23181_ _23181_/A vssd1 vssd1 vccd1 vccd1 _23412_/D sky130_fd_sc_hd__clkbuf_1
X_20393_ _20393_/A _20393_/B vssd1 vssd1 vccd1 vccd1 _20394_/B sky130_fd_sc_hd__or2_1
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_516 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22132_ _13392_/A _13392_/B _22121_/A vssd1 vssd1 vccd1 vccd1 _22132_/X sky130_fd_sc_hd__a21o_1
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22063_ _22130_/A _22136_/A _22062_/X vssd1 vssd1 vccd1 vccd1 _22211_/A sky130_fd_sc_hd__a21oi_2
XFILLER_160_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18988__B1 _19156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21014_ _21000_/A _21000_/B _21001_/Y vssd1 vssd1 vccd1 vccd1 _21014_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21276__A _21276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22965_ _22965_/A vssd1 vssd1 vccd1 vccd1 _23316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21916_ _21916_/A _22045_/A vssd1 vssd1 vccd1 vccd1 _21916_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22896_ input40/X _23184_/B input6/X _22896_/D vssd1 vssd1 vccd1 vccd1 _22953_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21847_ _21847_/A _21847_/B _21847_/C vssd1 vssd1 vccd1 vccd1 _21858_/D sky130_fd_sc_hd__nand3_4
XFILLER_130_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11600_ _18947_/B vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16536__C _17450_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12580_ _12580_/A vssd1 vssd1 vccd1 vccd1 _13019_/B sky130_fd_sc_hd__buf_2
XFILLER_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21778_ _22487_/A _22364_/B _21778_/C _21778_/D vssd1 vssd1 vccd1 vccd1 _21778_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20729_ _20523_/A _20523_/B _20523_/C _20713_/B vssd1 vssd1 vccd1 vccd1 _20729_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_8_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23517_ _23518_/CLK input42/X vssd1 vssd1 vccd1 vccd1 _23517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19847__C _19847_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14250_ _14245_/Y _14248_/Y _14253_/A _14253_/B vssd1 vssd1 vccd1 vccd1 _14255_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_139_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23448_ _23462_/CLK hold5/X vssd1 vssd1 vccd1 vccd1 _23448_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_184_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _13201_/A _13201_/B _13201_/C vssd1 vssd1 vccd1 vccd1 _13202_/A sky130_fd_sc_hd__nand3_4
XFILLER_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ _14181_/A vssd1 vssd1 vccd1 vccd1 _14181_/X sky130_fd_sc_hd__buf_2
XFILLER_87_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23379_ _23443_/CLK _23379_/D vssd1 vssd1 vccd1 vccd1 _23379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13132_ _21435_/C vssd1 vssd1 vccd1 vccd1 _21548_/B sky130_fd_sc_hd__buf_2
XFILLER_87_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16151__B1 _16447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18691__A2 _17643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17940_ _18198_/C _18256_/A _17933_/X vssd1 vssd1 vccd1 vccd1 _17942_/A sky130_fd_sc_hd__a21o_1
X_13063_ _13056_/X _12796_/A _12828_/Y _20529_/A _13054_/Y vssd1 vssd1 vccd1 vccd1
+ _13063_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17696__A1_N _23526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12014_ _11896_/A _11896_/B _11841_/Y _11840_/X _12118_/A vssd1 vssd1 vccd1 vccd1
+ _12029_/B sky130_fd_sc_hd__o221a_2
X_17871_ _17840_/Y _17842_/Y _17850_/Y vssd1 vssd1 vccd1 vccd1 _17874_/B sky130_fd_sc_hd__o21ai_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19610_ _19603_/Y _19422_/A _19606_/Y _19609_/Y vssd1 vssd1 vccd1 vccd1 _19620_/A
+ sky130_fd_sc_hd__o211ai_4
X_16822_ _15749_/A _15749_/B _16638_/X _16639_/X vssd1 vssd1 vccd1 vccd1 _16822_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_66_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19541_ _19547_/A _19537_/X _19538_/X _19542_/A vssd1 vssd1 vccd1 vccd1 _19560_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16753_ _16744_/Y _16750_/Y _16752_/Y vssd1 vssd1 vccd1 vccd1 _16792_/A sky130_fd_sc_hd__a21oi_2
X_13965_ _14029_/A vssd1 vssd1 vccd1 vccd1 _13965_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15704_ _15704_/A _15704_/B _15814_/A _15815_/A vssd1 vssd1 vccd1 vccd1 _15908_/A
+ sky130_fd_sc_hd__nand4_4
X_19472_ _19755_/A _19396_/A _19393_/Y vssd1 vssd1 vccd1 vccd1 _19472_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12916_ _13158_/A vssd1 vssd1 vccd1 vccd1 _13133_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_185_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16684_ _16684_/A vssd1 vssd1 vccd1 vccd1 _16684_/X sky130_fd_sc_hd__buf_4
XFILLER_0_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13896_ _14835_/C _14936_/B vssd1 vssd1 vccd1 vccd1 _14006_/A sky130_fd_sc_hd__nand2_1
XFILLER_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18423_ _18423_/A _18423_/B vssd1 vssd1 vccd1 vccd1 _23597_/D sky130_fd_sc_hd__nor2_1
XFILLER_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15635_ _15927_/A vssd1 vssd1 vccd1 vccd1 _16677_/B sky130_fd_sc_hd__buf_2
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12847_ _12723_/X _12725_/X _12733_/B _12728_/Y vssd1 vssd1 vccd1 vccd1 _12859_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _18305_/X _18353_/Y _18305_/A vssd1 vssd1 vccd1 vccd1 _18356_/A sky130_fd_sc_hd__o21bai_1
X_15566_ _23446_/D _15563_/Y _15566_/S vssd1 vssd1 vccd1 vccd1 _15567_/A sky130_fd_sc_hd__mux2_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12845_/A _12846_/A _12777_/A vssd1 vssd1 vccd1 vccd1 _12779_/C sky130_fd_sc_hd__a21o_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _14729_/A _11807_/X _12040_/X _17631_/A _17712_/D vssd1 vssd1 vccd1 vccd1
+ _17305_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_159_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14517_ _14519_/D _14633_/B _14633_/C _14633_/A vssd1 vssd1 vccd1 vccd1 _14549_/A
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__13151__B _13151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18285_ _18285_/A _18285_/B vssd1 vssd1 vccd1 vccd1 _18286_/B sky130_fd_sc_hd__xor2_1
XFILLER_159_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11729_ _19161_/A vssd1 vssd1 vccd1 vccd1 _16497_/A sky130_fd_sc_hd__clkbuf_4
X_15497_ _15494_/X _15497_/B _15516_/A vssd1 vssd1 vccd1 vccd1 _15497_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_30_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17236_ _17420_/B _17236_/B _17236_/C _19949_/D vssd1 vssd1 vccd1 vccd1 _17238_/B
+ sky130_fd_sc_hd__nand4_1
X_14448_ _14448_/A vssd1 vssd1 vccd1 vccd1 _15118_/A sky130_fd_sc_hd__buf_2
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16462__B _16462_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15359__A _15488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17167_ _17334_/A _17335_/A _17167_/C _17167_/D vssd1 vssd1 vccd1 vccd1 _17172_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18667__C1 _18666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14379_ _14377_/A _15358_/A _14377_/C vssd1 vssd1 vccd1 vccd1 _14380_/B sky130_fd_sc_hd__a21oi_1
XFILLER_155_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16118_ _15949_/X _16015_/Y _16002_/B _16249_/B vssd1 vssd1 vccd1 vccd1 _16248_/B
+ sky130_fd_sc_hd__o211ai_2
X_17098_ _18859_/A _17098_/B _17098_/C _17108_/B vssd1 vssd1 vccd1 vccd1 _17098_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_115_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_986 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17890__B1 _17889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16049_ _16490_/A _17414_/D _17414_/C _16049_/D vssd1 vssd1 vccd1 vccd1 _16757_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_170_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12703__B1 _13151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13604__B1_N _13603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20431__C _20431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20241__A2 _20242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19808_ _19803_/X _18003_/A _19701_/B _19807_/X vssd1 vssd1 vccd1 vccd1 _19975_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_96_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13607__A _23472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22518__A1 _22521_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15653__C1 _16866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19739_ _19560_/Y _19728_/X _19719_/Y _19893_/A vssd1 vssd1 vccd1 vccd1 _19893_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_38_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16918__A _23428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__23191__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22750_ _22750_/A _22750_/B vssd1 vssd1 vccd1 vccd1 _22774_/A sky130_fd_sc_hd__and2_1
XANTENNA__23461__D _23473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21701_ _23574_/Q _21716_/B _21716_/C vssd1 vssd1 vccd1 vccd1 _21723_/A sky130_fd_sc_hd__nand3b_1
X_22681_ _22605_/A _22633_/Y _22679_/Y _22680_/X vssd1 vssd1 vccd1 vccd1 _22683_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_53_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21632_ _21666_/A vssd1 vssd1 vccd1 vccd1 _21632_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18852__B _18959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21563_ _21564_/B _21564_/C _21564_/A vssd1 vssd1 vccd1 vccd1 _21565_/A sky130_fd_sc_hd__a21oi_1
XFILLER_139_928 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16075__D _16539_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19667__C _19675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23302_ _23398_/CLK _23302_/D vssd1 vssd1 vccd1 vccd1 _23302_/Q sky130_fd_sc_hd__dfxtp_1
X_20514_ _20507_/X _20501_/X _20510_/Y _20518_/A _20492_/B vssd1 vssd1 vccd1 vccd1
+ _20515_/C sky130_fd_sc_hd__o2111ai_1
X_21494_ _21495_/C _21495_/A _21495_/B vssd1 vssd1 vccd1 vccd1 _21559_/A sky130_fd_sc_hd__a21oi_1
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16920__A2 _16668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23233_ _23435_/Q input20/X _23239_/S vssd1 vssd1 vccd1 vccd1 _23234_/A sky130_fd_sc_hd__mux2_1
X_20445_ _20446_/A _20446_/B _20446_/C _20031_/X _23558_/Q vssd1 vssd1 vccd1 vccd1
+ _20448_/A sky130_fd_sc_hd__a311o_1
XFILLER_10_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16133__B1 _16124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23164_ _23164_/A vssd1 vssd1 vccd1 vccd1 _23404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20376_ _20376_/A _20376_/B _20401_/B vssd1 vssd1 vccd1 vccd1 _20378_/A sky130_fd_sc_hd__or3_1
XFILLER_122_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22115_ _22115_/A _22115_/B vssd1 vssd1 vccd1 vccd1 _23562_/D sky130_fd_sc_hd__xnor2_4
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23095_ _23374_/Q input23/X _23095_/S vssd1 vssd1 vccd1 vccd1 _23096_/A sky130_fd_sc_hd__mux2_1
X_22046_ _21906_/A _22037_/X _21913_/B vssd1 vssd1 vccd1 vccd1 _22046_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__19622__B2 _19380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16436__A1 _11882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16436__B2 _15749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23590__CLK _23598_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__23182__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13750_ _13739_/A _13739_/B _13739_/C _22465_/D _13743_/A vssd1 vssd1 vccd1 vccd1
+ _13750_/X sky130_fd_sc_hd__o311a_1
X_22948_ _22948_/A vssd1 vssd1 vccd1 vccd1 _23308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_86 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12701_ _13041_/B _13184_/A _12812_/A _12700_/Y vssd1 vssd1 vccd1 vccd1 _13138_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13681_ _13671_/A _13671_/B _13679_/Y _13680_/X vssd1 vssd1 vccd1 vccd1 _13682_/C
+ sky130_fd_sc_hd__o2bb2ai_1
X_22879_ _22878_/A _22887_/C _22878_/B vssd1 vssd1 vccd1 vccd1 _22887_/B sky130_fd_sc_hd__a21o_1
X_15420_ _15420_/A _15485_/D _15420_/C _15420_/D vssd1 vssd1 vccd1 vccd1 _15420_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_19_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12632_ _12632_/A vssd1 vssd1 vccd1 vccd1 _12633_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15170__C _15238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12563_ _12563_/A _12563_/B _12563_/C vssd1 vssd1 vccd1 vccd1 _12563_/Y sky130_fd_sc_hd__nor3_2
X_15351_ _15455_/A vssd1 vssd1 vccd1 vccd1 _15508_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18481__C _18481_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14302_ _14294_/B _14302_/B _14302_/C vssd1 vssd1 vccd1 vccd1 _14310_/D sky130_fd_sc_hd__nand3b_1
X_18070_ _17928_/Y _17929_/X _17930_/Y vssd1 vssd1 vccd1 vccd1 _18070_/Y sky130_fd_sc_hd__a21oi_1
X_12494_ _12494_/A _12494_/B _12494_/C vssd1 vssd1 vccd1 vccd1 _12536_/B sky130_fd_sc_hd__nand3_2
XFILLER_8_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15282_ _15282_/A _15282_/B vssd1 vssd1 vccd1 vccd1 _15282_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17021_ _16996_/Y _17381_/B _17020_/X vssd1 vssd1 vccd1 vccd1 _23583_/D sky130_fd_sc_hd__o21a_1
X_14233_ _14826_/A _14826_/B _14826_/C vssd1 vssd1 vccd1 vccd1 _14235_/B sky130_fd_sc_hd__nand3_1
XFILLER_172_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12933__B1 _13177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ _14164_/A _14164_/B vssd1 vssd1 vccd1 vccd1 _14164_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__21909__A _22064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13115_ _13115_/A _13115_/B _21174_/B vssd1 vssd1 vccd1 vccd1 _13115_/X sky130_fd_sc_hd__and3_1
X_14095_ _14078_/Y _14094_/X _14193_/C vssd1 vssd1 vccd1 vccd1 _14184_/B sky130_fd_sc_hd__a21o_2
X_18972_ _18972_/A _18972_/B _18972_/C vssd1 vssd1 vccd1 vccd1 _18981_/A sky130_fd_sc_hd__nand3_2
XFILLER_125_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20532__B _20532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _17920_/B _17920_/C _17920_/A vssd1 vssd1 vccd1 vccd1 _17924_/C sky130_fd_sc_hd__a21oi_1
XFILLER_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13001_/X _13029_/Y _13030_/Y _13031_/Y vssd1 vssd1 vccd1 vccd1 _20556_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_26_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17854_ _17855_/A _17982_/A _17982_/B vssd1 vssd1 vccd1 vccd1 _17857_/B sky130_fd_sc_hd__a21bo_1
XFILLER_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16805_ _16805_/A _17569_/A _17040_/A vssd1 vssd1 vccd1 vccd1 _16805_/X sky130_fd_sc_hd__and3_1
XANTENNA__20774__A3 _20773_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17785_ _17783_/X _17784_/Y _17782_/A vssd1 vssd1 vccd1 vccd1 _17785_/Y sky130_fd_sc_hd__o21bai_1
X_14997_ _15094_/A vssd1 vssd1 vccd1 vccd1 _15096_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19524_ _19524_/A _19524_/B _19524_/C vssd1 vssd1 vccd1 vccd1 _19578_/A sky130_fd_sc_hd__nand3_4
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16736_ _16240_/Y _16251_/X _16246_/C vssd1 vssd1 vccd1 vccd1 _16737_/A sky130_fd_sc_hd__o21ai_1
XFILLER_19_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13948_ _14044_/B vssd1 vssd1 vccd1 vccd1 _13948_/X sky130_fd_sc_hd__buf_2
X_19455_ _23544_/Q _19457_/C _19457_/A _19291_/Y vssd1 vssd1 vccd1 vccd1 _19456_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16667_ _15599_/X _16667_/B _16667_/C _16667_/D vssd1 vssd1 vccd1 vccd1 _16668_/B
+ sky130_fd_sc_hd__nand4b_4
XANTENNA__15938__B1 _16281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13879_ _14001_/A vssd1 vssd1 vccd1 vccd1 _14430_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_62_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18406_ _18407_/B _18407_/C _18407_/D _18407_/A vssd1 vssd1 vccd1 vccd1 _18406_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_62_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15618_ _15618_/A vssd1 vssd1 vccd1 vccd1 _15618_/X sky130_fd_sc_hd__buf_4
X_19386_ _19221_/Y _19216_/Y _19212_/Y vssd1 vssd1 vccd1 vccd1 _19389_/A sky130_fd_sc_hd__a21oi_2
XFILLER_72_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16598_ _16598_/A _16598_/B vssd1 vssd1 vccd1 vccd1 _16598_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18672__B _18868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18337_ _18378_/B _18337_/B vssd1 vssd1 vccd1 vccd1 _18338_/B sky130_fd_sc_hd__nand2_1
X_15549_ _15522_/A _15526_/A _15548_/Y vssd1 vssd1 vccd1 vccd1 _15558_/C sky130_fd_sc_hd__o21a_1
XANTENNA__12621__C1 _20894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18268_ _18268_/A _18268_/B vssd1 vssd1 vccd1 vccd1 _18288_/A sky130_fd_sc_hd__nand2_1
XANTENNA__23463__CLK _23559_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16902__A2 _12006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_bq_clk_i clkbuf_3_5_0_bq_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_bq_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_17219_ _17189_/B _17189_/A _17187_/B vssd1 vssd1 vccd1 vccd1 _17347_/A sky130_fd_sc_hd__o21ai_1
X_18199_ _18154_/X _18196_/X _18302_/C _23532_/Q vssd1 vssd1 vccd1 vccd1 _18199_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_175_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12506__A _12506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20230_ _20158_/B _20159_/B _20224_/Y _20225_/X vssd1 vssd1 vccd1 vccd1 _20231_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_116_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16666__A1 _16781_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22641__C _22647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20161_ _20167_/B _20232_/A _20167_/A vssd1 vssd1 vccd1 vccd1 _20161_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14721__A _14729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1098 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20092_ _20087_/Y _20175_/C _20091_/Y vssd1 vssd1 vccd1 vccd1 _20099_/B sky130_fd_sc_hd__o21ai_1
XFILLER_69_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12152__A1 _16437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_872 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12152__B2 _12151_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12241__A _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19024__A _19029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15552__A _15552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22802_ _22829_/B _22799_/Y _22801_/X vssd1 vssd1 vccd1 vccd1 _22802_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20994_ _20994_/A _20994_/B _20994_/C vssd1 vssd1 vccd1 vccd1 _20995_/C sky130_fd_sc_hd__nand3_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13652__A1 _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21704__D _21704_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22733_ _22731_/B _22732_/X _22731_/A vssd1 vssd1 vccd1 vccd1 _22734_/A sky130_fd_sc_hd__a21oi_1
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16051__C1 _16372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22664_ _21777_/A _21777_/B _21829_/A vssd1 vssd1 vccd1 vccd1 _22664_/X sky130_fd_sc_hd__a21o_1
XFILLER_198_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22385__A _22479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21615_ _21630_/A _21666_/B _21614_/Y _21694_/C vssd1 vssd1 vccd1 vccd1 _21615_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22595_ _22505_/X _22507_/Y _22511_/Y _22509_/X vssd1 vssd1 vccd1 vccd1 _22595_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_178_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17146__A2 _11883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21546_ _21546_/A vssd1 vssd1 vccd1 vccd1 _21637_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17551__C1 _17546_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19694__A _19694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13707__A2 _21987_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21477_ _21477_/A _21477_/B vssd1 vssd1 vccd1 vccd1 _21477_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11718__A1 _12323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23216_ _23216_/A vssd1 vssd1 vccd1 vccd1 _23427_/D sky130_fd_sc_hd__clkbuf_1
X_20428_ _20428_/A _20428_/B _20428_/C vssd1 vssd1 vccd1 vccd1 _20429_/S sky130_fd_sc_hd__or3_1
XANTENNA__20055__D _20055_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23147_ _23169_/A vssd1 vssd1 vccd1 vccd1 _23156_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20359_ _20359_/A _20359_/B _20359_/C _20359_/D vssd1 vssd1 vccd1 vccd1 _20359_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_945 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23078_ _23366_/Q input14/X _23084_/S vssd1 vssd1 vccd1 vccd1 _23079_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22029_ _22029_/A vssd1 vssd1 vccd1 vccd1 _22141_/C sky130_fd_sc_hd__clkbuf_2
X_14920_ _14795_/Y _14796_/Y _14797_/X _14798_/Y vssd1 vssd1 vccd1 vccd1 _14923_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__17606__B1 _17753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input25_A wb_dat_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851_ _14853_/A _14501_/B _14749_/X _14845_/Y _14850_/Y vssd1 vssd1 vccd1 vccd1
+ _23271_/D sky130_fd_sc_hd__a41o_1
XANTENNA__16558__A _16558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19359__B1 _19358_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _13802_/A _13802_/B vssd1 vssd1 vccd1 vccd1 _13803_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17570_ _17249_/X _17250_/X _16056_/X _20317_/B vssd1 vssd1 vccd1 vccd1 _17737_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_1_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21166__B1 _21387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12446__A2 _12247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14782_ _14788_/A _14857_/A _14788_/C vssd1 vssd1 vccd1 vccd1 _14782_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11994_ _12099_/D _12121_/A vssd1 vssd1 vccd1 vccd1 _12426_/B sky130_fd_sc_hd__nand2_2
XFILLER_17_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16521_ _16566_/B _16566_/C _16566_/A vssd1 vssd1 vccd1 vccd1 _16759_/B sky130_fd_sc_hd__a21o_1
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13733_ _13707_/X _13731_/X _13732_/X vssd1 vssd1 vccd1 vccd1 _13739_/A sky130_fd_sc_hd__a21oi_2
XFILLER_189_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19240_ _19240_/A _19240_/B vssd1 vssd1 vccd1 vccd1 _19240_/Y sky130_fd_sc_hd__nand2_2
XFILLER_182_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ _16457_/A _16457_/B _16451_/X vssd1 vssd1 vccd1 vccd1 _16452_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13664_ _13769_/A _13497_/A _13663_/Y _13661_/Y vssd1 vssd1 vccd1 vccd1 _13666_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15403_ _15403_/A vssd1 vssd1 vccd1 vccd1 _15404_/A sky130_fd_sc_hd__inv_2
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19171_ _18978_/B _18975_/X _19158_/A _18971_/X vssd1 vssd1 vccd1 vccd1 _19172_/C
+ sky130_fd_sc_hd__o2bb2ai_4
X_12615_ _20784_/C vssd1 vssd1 vccd1 vccd1 _21039_/B sky130_fd_sc_hd__clkbuf_2
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16383_ _16225_/X _17285_/A _16318_/A vssd1 vssd1 vccd1 vccd1 _16383_/X sky130_fd_sc_hd__o21a_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18334__A1 _20369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13595_ _13540_/A _13540_/C _13540_/B vssd1 vssd1 vccd1 vccd1 _13595_/Y sky130_fd_sc_hd__a21oi_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18334__B2 _18157_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18122_ _18134_/B vssd1 vssd1 vccd1 vccd1 _18122_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11957__B2 _17642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _15292_/B _15292_/A _15279_/B _15332_/X vssd1 vssd1 vccd1 vccd1 _15335_/B
+ sky130_fd_sc_hd__o211ai_4
X_12546_ _12546_/A _12546_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12565_/C sky130_fd_sc_hd__and3_1
XFILLER_184_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18053_ _18053_/A _18129_/A vssd1 vssd1 vccd1 vccd1 _18138_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16443__D _19503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15265_ _15265_/A vssd1 vssd1 vccd1 vccd1 _15363_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_184_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12477_ _12478_/A _12478_/B _12478_/C vssd1 vssd1 vccd1 vccd1 _12480_/A sky130_fd_sc_hd__a21oi_1
X_17004_ _23521_/Q vssd1 vssd1 vccd1 vccd1 _17014_/A sky130_fd_sc_hd__inv_2
XANTENNA_output93_A _23267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _14220_/A _14220_/B _14221_/B vssd1 vssd1 vccd1 vccd1 _14218_/B sky130_fd_sc_hd__nand3_1
XFILLER_125_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15196_ _14981_/X _14976_/Y _14985_/X _15090_/Y vssd1 vssd1 vccd1 vccd1 _15196_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14147_ _14222_/A _14222_/B _14217_/C _14218_/A vssd1 vssd1 vccd1 vccd1 _14148_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21358__B _21358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18955_ _18942_/B _18942_/A _18944_/C vssd1 vssd1 vccd1 vccd1 _18955_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15320__B2 _15422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078_ _14078_/A _14189_/A _14864_/B _14191_/C vssd1 vssd1 vccd1 vccd1 _14078_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12134__B2 _19363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13157__A _21279_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17906_ _17782_/A _17782_/B _17784_/Y vssd1 vssd1 vccd1 vccd1 _17909_/A sky130_fd_sc_hd__a21oi_1
XFILLER_140_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13029_ _13029_/A _13029_/B vssd1 vssd1 vccd1 vccd1 _13029_/Y sky130_fd_sc_hd__nand2_1
X_18886_ _18879_/Y _18882_/Y _18884_/Y _18885_/Y vssd1 vssd1 vccd1 vccd1 _18886_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_117_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17837_ _17708_/Y _17805_/Y _17805_/A vssd1 vssd1 vccd1 vccd1 _17920_/A sky130_fd_sc_hd__o21ai_2
XFILLER_55_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1047 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17768_ _17773_/A _17773_/B _17765_/X _17767_/X vssd1 vssd1 vccd1 vccd1 _17768_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_81_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19507_ _19656_/A _19491_/B _19649_/B _18656_/Y vssd1 vssd1 vccd1 vccd1 _19507_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16719_ _16010_/X _16176_/Y _16253_/B _16253_/A vssd1 vssd1 vccd1 vccd1 _16719_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_17699_ _17699_/A vssd1 vssd1 vccd1 vccd1 _17928_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19438_ _19638_/A _19616_/A _19616_/B vssd1 vssd1 vccd1 vccd1 _19438_/Y sky130_fd_sc_hd__nand3_1
XFILLER_179_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19369_ _19369_/A _19369_/B _19369_/C vssd1 vssd1 vccd1 vccd1 _19568_/A sky130_fd_sc_hd__nand3_2
XFILLER_163_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21400_ _21400_/A _21400_/B vssd1 vssd1 vccd1 vccd1 _21476_/B sky130_fd_sc_hd__and2_1
XFILLER_31_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16634__C _16634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20132__A1 _20133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22380_ _22637_/A _22637_/B _22380_/C vssd1 vssd1 vccd1 vccd1 _22386_/B sky130_fd_sc_hd__nand3_1
XFILLER_198_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18876__A2 _18875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21331_ _21266_/X _21331_/B _21331_/C vssd1 vssd1 vccd1 vccd1 _21333_/C sky130_fd_sc_hd__nand3b_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12236__A _16408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18089__B1 _12088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21262_ _21260_/Y _21262_/B vssd1 vssd1 vccd1 vccd1 _21263_/A sky130_fd_sc_hd__and2b_1
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13165__A3 _20773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19825__A1 _20081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19664__D _19969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23001_ _22142_/B input12/X _23001_/S vssd1 vssd1 vccd1 vccd1 _23002_/A sky130_fd_sc_hd__mux2_1
X_20213_ _19700_/A _19700_/B _20268_/D _20287_/A _20212_/C vssd1 vssd1 vccd1 vccd1
+ _20277_/B sky130_fd_sc_hd__a32o_1
XFILLER_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19019__A _19327_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21193_ _21493_/A _21493_/B _21193_/C vssd1 vssd1 vccd1 vccd1 _21194_/B sky130_fd_sc_hd__nand3_1
XFILLER_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20144_ _20050_/Y _20056_/B _20048_/Y _20045_/Y vssd1 vssd1 vccd1 vccd1 _20148_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__22090__D _22090_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16091__A1_N _16469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20075_ _20070_/Y _20172_/A _20074_/X vssd1 vssd1 vccd1 vccd1 _20095_/A sky130_fd_sc_hd__a21o_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23137__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16811__A1 _15742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13625__A1 _13486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15713__C _15713_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20977_ _20977_/A _20984_/A vssd1 vssd1 vccd1 vccd1 _20980_/B sky130_fd_sc_hd__nand2_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22716_ _22716_/A _22789_/A _22716_/C _22716_/D vssd1 vssd1 vccd1 vccd1 _22789_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17772__C1 _17771_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19201__B _19709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22647_ _22647_/A vssd1 vssd1 vccd1 vccd1 _22701_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19513__B1 _19656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ _12491_/A _12491_/B _12217_/B vssd1 vssd1 vccd1 vccd1 _12400_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13530__A _21921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13380_ _13602_/C _13264_/B _13379_/X vssd1 vssd1 vccd1 vccd1 _13423_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11969__B _11969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22578_ _13547_/A _22461_/A _22635_/A vssd1 vssd1 vccd1 vccd1 _22578_/X sky130_fd_sc_hd__o21a_1
XFILLER_142_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12331_ _12360_/A _12360_/B _12318_/A _12321_/A _12330_/X vssd1 vssd1 vccd1 vccd1
+ _12336_/B sky130_fd_sc_hd__a41o_1
XANTENNA__20674__A2 _12637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21529_ _21529_/A vssd1 vssd1 vccd1 vccd1 _21529_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12146__A _16802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23073__A0 _23364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12262_ _12475_/B _12262_/B _12306_/A _18531_/A vssd1 vssd1 vccd1 vccd1 _12265_/C
+ sky130_fd_sc_hd__nand4_1
X_15050_ _15050_/A _15050_/B _15050_/C vssd1 vssd1 vccd1 vccd1 _15052_/B sky130_fd_sc_hd__nand3_1
XFILLER_154_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14001_ _14001_/A vssd1 vssd1 vccd1 vccd1 _14433_/D sky130_fd_sc_hd__buf_2
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12193_ _12183_/X _12188_/Y _12191_/Y _12192_/Y vssd1 vssd1 vccd1 vccd1 _12206_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_134_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput63 _14671_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput74 _14711_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput85 _14603_/X vssd1 vssd1 vccd1 vccd1 wb_dat_o[9] sky130_fd_sc_hd__buf_2
Xoutput96 _23579_/Q vssd1 vssd1 vccd1 vccd1 y[8] sky130_fd_sc_hd__buf_2
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18740_ _18579_/Y _18574_/X _18588_/A vssd1 vssd1 vccd1 vccd1 _18740_/Y sky130_fd_sc_hd__o21ai_1
X_15952_ _15742_/X _16447_/B _19703_/C vssd1 vssd1 vccd1 vccd1 _15998_/A sky130_fd_sc_hd__o21ai_4
XFILLER_95_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14903_ _14903_/A _14903_/B vssd1 vssd1 vccd1 vccd1 _14968_/A sky130_fd_sc_hd__nand2_1
XFILLER_49_756 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17391__B _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18671_ _18670_/Y _18627_/Y _18465_/X vssd1 vssd1 vccd1 vccd1 _18868_/C sky130_fd_sc_hd__o21ai_2
X_15883_ _15883_/A vssd1 vssd1 vccd1 vccd1 _15884_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16288__A _17845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__23128__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ _17622_/A _17622_/B _17622_/C vssd1 vssd1 vccd1 vccd1 _17656_/B sky130_fd_sc_hd__nand3_1
X_14834_ _14834_/A vssd1 vssd1 vccd1 vccd1 _15298_/B sky130_fd_sc_hd__buf_2
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18004__B1 _18211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _17553_/A _17791_/A vssd1 vssd1 vccd1 vccd1 _17553_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11627__B1 _16815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _14174_/B _14887_/A _14183_/A _14753_/Y _15301_/A vssd1 vssd1 vccd1 vccd1
+ _14766_/B sky130_fd_sc_hd__o2111ai_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11977_ _23387_/Q _11977_/B _23388_/Q vssd1 vssd1 vccd1 vccd1 _18469_/B sky130_fd_sc_hd__nor3_4
XFILLER_91_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16504_ _16389_/X _16523_/D _16496_/X _16502_/X _16503_/Y vssd1 vssd1 vccd1 vccd1
+ _16530_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_32_612 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15920__A _15920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13716_ _13711_/A _13711_/B _13711_/C vssd1 vssd1 vccd1 vccd1 _13716_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__20362__A1 _20031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17484_ _17485_/A _17485_/B _17485_/C vssd1 vssd1 vccd1 vccd1 _17654_/A sky130_fd_sc_hd__a21oi_1
X_14696_ _23374_/Q _14688_/X _14695_/X vssd1 vssd1 vccd1 vccd1 _14696_/X sky130_fd_sc_hd__o21a_1
XFILLER_189_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19223_ _19176_/Y _19179_/Y _19189_/A vssd1 vssd1 vccd1 vccd1 _19230_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16435_ _16435_/A _16435_/B _16435_/C vssd1 vssd1 vccd1 vccd1 _16765_/A sky130_fd_sc_hd__nand3_2
XFILLER_20_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13647_ _13419_/X _13443_/A _13432_/Y _13434_/Y vssd1 vssd1 vccd1 vccd1 _13647_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19154_ _16054_/A _16055_/A _19505_/A _19504_/A _19502_/A vssd1 vssd1 vccd1 vccd1
+ _19309_/A sky130_fd_sc_hd__o221ai_4
XFILLER_169_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16366_ _16366_/A _16366_/B vssd1 vssd1 vccd1 vccd1 _16399_/A sky130_fd_sc_hd__nand2_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13578_ _13556_/X _13557_/Y _13577_/Y vssd1 vssd1 vccd1 vccd1 _13578_/Y sky130_fd_sc_hd__o21ai_1
X_18105_ _18179_/A _18104_/B _18090_/A _18090_/B vssd1 vssd1 vccd1 vccd1 _18106_/C
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_158_886 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15317_ _15317_/A vssd1 vssd1 vccd1 vccd1 _15419_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19085_ _19087_/A _19087_/B _18617_/X _18928_/X vssd1 vssd1 vccd1 vccd1 _19088_/B
+ sky130_fd_sc_hd__o2bb2ai_2
X_12529_ _12529_/A _12529_/B _12529_/C vssd1 vssd1 vccd1 vccd1 _12540_/C sky130_fd_sc_hd__nand3_1
XFILLER_9_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16297_ _16297_/A _16297_/B vssd1 vssd1 vccd1 vccd1 _16297_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18036_ _18036_/A _18036_/B vssd1 vssd1 vccd1 vccd1 _18038_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15541__A1 _15225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15248_ _15250_/C _15250_/D _15247_/Y vssd1 vssd1 vccd1 vccd1 _15270_/B sky130_fd_sc_hd__a21o_1
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14271__A _14777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ _15179_/A _15179_/B _15179_/C vssd1 vssd1 vccd1 vccd1 _15249_/B sky130_fd_sc_hd__nand3_1
XFILLER_113_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19987_ _19987_/A _19987_/B _19987_/C vssd1 vssd1 vccd1 vccd1 _19987_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__18678__A _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17582__A _17845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18938_ _18938_/A vssd1 vssd1 vccd1 vccd1 _18938_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
.ends

