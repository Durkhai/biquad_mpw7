VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bqmain
  CLASS BLOCK ;
  FOREIGN bqmain ;
  ORIGIN 0.000 0.000 ;
  SIZE 547.300 BY 558.020 ;
  PIN bq_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END bq_clk_i
  PIN nreset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 554.020 22.450 558.020 ;
    END
  END nreset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 546.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 546.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 546.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 546.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 546.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 546.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 546.960 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 4.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END wb_adr_i[24]
  PIN wb_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END wb_adr_i[25]
  PIN wb_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END wb_adr_i[26]
  PIN wb_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END wb_adr_i[27]
  PIN wb_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END wb_adr_i[28]
  PIN wb_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END wb_adr_i[29]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END wb_adr_i[30]
  PIN wb_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END wb_adr_i[31]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wb_dat_o[9]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END wb_rst_i
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wb_we_i
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 24.520 547.300 25.120 ;
    END
  END x[0]
  PIN x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 486.920 547.300 487.520 ;
    END
  END x[10]
  PIN x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 533.160 547.300 533.760 ;
    END
  END x[11]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 70.760 547.300 71.360 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 117.000 547.300 117.600 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 163.240 547.300 163.840 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 209.480 547.300 210.080 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 255.720 547.300 256.320 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 301.960 547.300 302.560 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 348.200 547.300 348.800 ;
    END
  END x[7]
  PIN x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 394.440 547.300 395.040 ;
    END
  END x[8]
  PIN x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 543.300 440.680 547.300 441.280 ;
    END
  END x[9]
  PIN y[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 554.020 64.310 558.020 ;
    END
  END y[0]
  PIN y[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 554.020 482.910 558.020 ;
    END
  END y[10]
  PIN y[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 554.020 524.770 558.020 ;
    END
  END y[11]
  PIN y[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 554.020 106.170 558.020 ;
    END
  END y[1]
  PIN y[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 554.020 148.030 558.020 ;
    END
  END y[2]
  PIN y[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 554.020 189.890 558.020 ;
    END
  END y[3]
  PIN y[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 554.020 231.750 558.020 ;
    END
  END y[4]
  PIN y[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 554.020 273.610 558.020 ;
    END
  END y[5]
  PIN y[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 554.020 315.470 558.020 ;
    END
  END y[6]
  PIN y[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 554.020 357.330 558.020 ;
    END
  END y[7]
  PIN y[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 554.020 399.190 558.020 ;
    END
  END y[8]
  PIN y[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 554.020 441.050 558.020 ;
    END
  END y[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 541.420 546.805 ;
      LAYER met1 ;
        RECT 1.450 2.760 541.420 549.400 ;
      LAYER met2 ;
        RECT 1.470 553.740 21.890 556.765 ;
        RECT 22.730 553.740 63.750 556.765 ;
        RECT 64.590 553.740 105.610 556.765 ;
        RECT 106.450 553.740 147.470 556.765 ;
        RECT 148.310 553.740 189.330 556.765 ;
        RECT 190.170 553.740 231.190 556.765 ;
        RECT 232.030 553.740 273.050 556.765 ;
        RECT 273.890 553.740 314.910 556.765 ;
        RECT 315.750 553.740 356.770 556.765 ;
        RECT 357.610 553.740 398.630 556.765 ;
        RECT 399.470 553.740 440.490 556.765 ;
        RECT 441.330 553.740 482.350 556.765 ;
        RECT 483.190 553.740 524.210 556.765 ;
        RECT 525.050 553.740 540.410 556.765 ;
        RECT 1.470 4.280 540.410 553.740 ;
        RECT 1.470 2.730 14.990 4.280 ;
        RECT 15.830 2.730 20.050 4.280 ;
        RECT 20.890 2.730 25.110 4.280 ;
        RECT 25.950 2.730 30.170 4.280 ;
        RECT 31.010 2.730 35.230 4.280 ;
        RECT 36.070 2.730 40.290 4.280 ;
        RECT 41.130 2.730 45.350 4.280 ;
        RECT 46.190 2.730 50.410 4.280 ;
        RECT 51.250 2.730 55.470 4.280 ;
        RECT 56.310 2.730 60.530 4.280 ;
        RECT 61.370 2.730 65.590 4.280 ;
        RECT 66.430 2.730 70.650 4.280 ;
        RECT 71.490 2.730 75.710 4.280 ;
        RECT 76.550 2.730 80.770 4.280 ;
        RECT 81.610 2.730 85.830 4.280 ;
        RECT 86.670 2.730 90.890 4.280 ;
        RECT 91.730 2.730 95.950 4.280 ;
        RECT 96.790 2.730 101.010 4.280 ;
        RECT 101.850 2.730 106.070 4.280 ;
        RECT 106.910 2.730 111.130 4.280 ;
        RECT 111.970 2.730 116.190 4.280 ;
        RECT 117.030 2.730 121.250 4.280 ;
        RECT 122.090 2.730 126.310 4.280 ;
        RECT 127.150 2.730 131.370 4.280 ;
        RECT 132.210 2.730 136.430 4.280 ;
        RECT 137.270 2.730 141.490 4.280 ;
        RECT 142.330 2.730 146.550 4.280 ;
        RECT 147.390 2.730 151.610 4.280 ;
        RECT 152.450 2.730 156.670 4.280 ;
        RECT 157.510 2.730 161.730 4.280 ;
        RECT 162.570 2.730 166.790 4.280 ;
        RECT 167.630 2.730 171.850 4.280 ;
        RECT 172.690 2.730 176.910 4.280 ;
        RECT 177.750 2.730 181.970 4.280 ;
        RECT 182.810 2.730 187.030 4.280 ;
        RECT 187.870 2.730 192.090 4.280 ;
        RECT 192.930 2.730 197.150 4.280 ;
        RECT 197.990 2.730 202.210 4.280 ;
        RECT 203.050 2.730 207.270 4.280 ;
        RECT 208.110 2.730 212.330 4.280 ;
        RECT 213.170 2.730 217.390 4.280 ;
        RECT 218.230 2.730 222.450 4.280 ;
        RECT 223.290 2.730 227.510 4.280 ;
        RECT 228.350 2.730 232.570 4.280 ;
        RECT 233.410 2.730 237.630 4.280 ;
        RECT 238.470 2.730 242.690 4.280 ;
        RECT 243.530 2.730 247.750 4.280 ;
        RECT 248.590 2.730 252.810 4.280 ;
        RECT 253.650 2.730 257.870 4.280 ;
        RECT 258.710 2.730 262.930 4.280 ;
        RECT 263.770 2.730 267.990 4.280 ;
        RECT 268.830 2.730 273.050 4.280 ;
        RECT 273.890 2.730 278.110 4.280 ;
        RECT 278.950 2.730 283.170 4.280 ;
        RECT 284.010 2.730 288.230 4.280 ;
        RECT 289.070 2.730 293.290 4.280 ;
        RECT 294.130 2.730 298.350 4.280 ;
        RECT 299.190 2.730 303.410 4.280 ;
        RECT 304.250 2.730 308.470 4.280 ;
        RECT 309.310 2.730 313.530 4.280 ;
        RECT 314.370 2.730 318.590 4.280 ;
        RECT 319.430 2.730 323.650 4.280 ;
        RECT 324.490 2.730 328.710 4.280 ;
        RECT 329.550 2.730 333.770 4.280 ;
        RECT 334.610 2.730 338.830 4.280 ;
        RECT 339.670 2.730 343.890 4.280 ;
        RECT 344.730 2.730 348.950 4.280 ;
        RECT 349.790 2.730 354.010 4.280 ;
        RECT 354.850 2.730 359.070 4.280 ;
        RECT 359.910 2.730 364.130 4.280 ;
        RECT 364.970 2.730 369.190 4.280 ;
        RECT 370.030 2.730 374.250 4.280 ;
        RECT 375.090 2.730 379.310 4.280 ;
        RECT 380.150 2.730 384.370 4.280 ;
        RECT 385.210 2.730 389.430 4.280 ;
        RECT 390.270 2.730 394.490 4.280 ;
        RECT 395.330 2.730 399.550 4.280 ;
        RECT 400.390 2.730 404.610 4.280 ;
        RECT 405.450 2.730 409.670 4.280 ;
        RECT 410.510 2.730 414.730 4.280 ;
        RECT 415.570 2.730 419.790 4.280 ;
        RECT 420.630 2.730 424.850 4.280 ;
        RECT 425.690 2.730 429.910 4.280 ;
        RECT 430.750 2.730 434.970 4.280 ;
        RECT 435.810 2.730 440.030 4.280 ;
        RECT 440.870 2.730 445.090 4.280 ;
        RECT 445.930 2.730 450.150 4.280 ;
        RECT 450.990 2.730 455.210 4.280 ;
        RECT 456.050 2.730 460.270 4.280 ;
        RECT 461.110 2.730 465.330 4.280 ;
        RECT 466.170 2.730 470.390 4.280 ;
        RECT 471.230 2.730 475.450 4.280 ;
        RECT 476.290 2.730 480.510 4.280 ;
        RECT 481.350 2.730 485.570 4.280 ;
        RECT 486.410 2.730 490.630 4.280 ;
        RECT 491.470 2.730 495.690 4.280 ;
        RECT 496.530 2.730 500.750 4.280 ;
        RECT 501.590 2.730 505.810 4.280 ;
        RECT 506.650 2.730 510.870 4.280 ;
        RECT 511.710 2.730 515.930 4.280 ;
        RECT 516.770 2.730 520.990 4.280 ;
        RECT 521.830 2.730 526.050 4.280 ;
        RECT 526.890 2.730 531.110 4.280 ;
        RECT 531.950 2.730 540.410 4.280 ;
      LAYER met3 ;
        RECT 1.445 534.160 543.300 556.745 ;
        RECT 1.445 532.760 542.900 534.160 ;
        RECT 1.445 487.920 543.300 532.760 ;
        RECT 1.445 486.520 542.900 487.920 ;
        RECT 1.445 441.680 543.300 486.520 ;
        RECT 1.445 440.280 542.900 441.680 ;
        RECT 1.445 395.440 543.300 440.280 ;
        RECT 1.445 394.040 542.900 395.440 ;
        RECT 1.445 349.200 543.300 394.040 ;
        RECT 1.445 347.800 542.900 349.200 ;
        RECT 1.445 302.960 543.300 347.800 ;
        RECT 1.445 301.560 542.900 302.960 ;
        RECT 1.445 256.720 543.300 301.560 ;
        RECT 1.445 255.320 542.900 256.720 ;
        RECT 1.445 210.480 543.300 255.320 ;
        RECT 1.445 209.080 542.900 210.480 ;
        RECT 1.445 164.240 543.300 209.080 ;
        RECT 1.445 162.840 542.900 164.240 ;
        RECT 1.445 118.000 543.300 162.840 ;
        RECT 1.445 116.600 542.900 118.000 ;
        RECT 1.445 71.760 543.300 116.600 ;
        RECT 1.445 70.360 542.900 71.760 ;
        RECT 1.445 25.520 543.300 70.360 ;
        RECT 1.445 24.120 542.900 25.520 ;
        RECT 1.445 4.935 543.300 24.120 ;
      LAYER met4 ;
        RECT 2.135 547.360 532.385 556.745 ;
        RECT 2.135 10.240 20.640 547.360 ;
        RECT 23.040 10.240 97.440 547.360 ;
        RECT 99.840 10.240 174.240 547.360 ;
        RECT 176.640 10.240 251.040 547.360 ;
        RECT 253.440 10.240 327.840 547.360 ;
        RECT 330.240 10.240 404.640 547.360 ;
        RECT 407.040 10.240 481.440 547.360 ;
        RECT 483.840 10.240 532.385 547.360 ;
        RECT 2.135 5.615 532.385 10.240 ;
  END
END bqmain
END LIBRARY

